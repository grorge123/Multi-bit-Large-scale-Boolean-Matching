//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 , n513 , n514 , n515 , n516 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 , n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 , n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n299 , n300 , n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 , n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 , n332 , n333 , n334 , n335 , n336 , n337 , n338 , n339 , n340 , n341 , n342 , n343 , n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 , n354 , n355 , n356 , n357 , n358 , n359 , n360 , n361 , n362 , n363 , n364 , n365 , n366 , n367 , n368 , n369 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n377 , n378 , n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n388 , n389 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 , n398 , n399 , n400 , n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 , n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 , n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 , n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 , n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 , n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 ;
output n512 , n513 , n514 , n515 , n516 ;

wire n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 ,
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 ,
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 ,
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 ,
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 ,
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 ,
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 ,
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 ,
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 ,
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 ,
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 ,
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 ,
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 ,
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 ,
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 ,
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 ,
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 ,
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 ,
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 ,
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 ,
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 ,
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 ,
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 ,
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 ,
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 ,
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 ,
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 ,
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 ,
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 ,
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 ,
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 ,
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 ,
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 ,
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 ,
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 ,
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 ,
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 ,
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 ,
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 ,
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 ,
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 ,
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 ,
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 ,
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 ,
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 ,
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 ,
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 ,
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 ,
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 ,
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 ,
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 ,
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 ,
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 ,
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 ,
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 ,
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 ,
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 ,
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 ,
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 ,
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 ,
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 ,
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 ,
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 ,
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 ,
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 ,
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 ,
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 ,
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 ,
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 ,
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 ,
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 ,
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 ,
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 ,
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 ,
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 ,
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 ,
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 ,
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 ,
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 ,
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 ,
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 ,
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 ,
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 ,
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 ,
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 ,
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 ,
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 ,
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 ,
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 ,
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 ,
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 ,
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 ,
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 ,
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 ,
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 ,
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 ,
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 ,
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 ,
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 ,
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 ,
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 ,
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 ,
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 ,
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 ,
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 ,
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 ,
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 ,
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 ,
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 ,
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 ,
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 ,
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 ,
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 ,
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 ,
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 ,
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 ,
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 ,
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 ,
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 ,
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 ,
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 ,
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 ,
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 ,
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 ,
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 ,
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 ,
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 ,
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 ,
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 ,
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 ,
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 ,
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 ,
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 ,
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 ,
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 ,
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 ,
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 ,
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 ,
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 ,
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 ,
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 ,
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 ,
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 ,
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 ,
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 ,
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 ,
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 ,
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 ,
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 ,
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 ,
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 ,
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 ,
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 ,
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 ,
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 ,
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 ,
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 ,
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 ,
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 ,
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 ,
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 ,
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 ,
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 ,
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 ,
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 ,
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 ,
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 ,
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 ,
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 ,
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 ,
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 ,
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 ,
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 ,
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 ,
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 ,
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 ,
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 ,
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 ,
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 ,
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 ,
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 ,
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 ,
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 ,
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 ,
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 ,
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 ,
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 ,
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 ,
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 ,
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 ,
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 ,
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 ,
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 ,
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 ,
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 ,
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 ,
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 ,
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 ,
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 ,
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 ,
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 ,
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 ,
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 ,
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 ,
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 ,
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 ,
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 ;
buf ( n512 , n2322 );
buf ( n516 , n3095 );
buf ( n513 , n3097 );
buf ( n515 , n3098 );
buf ( n514 , n3099 );
buf ( n1036 , n49 );
buf ( n1037 , n369 );
buf ( n1038 , n424 );
buf ( n1039 , n418 );
buf ( n1040 , n110 );
buf ( n1041 , n35 );
buf ( n1042 , n340 );
buf ( n1043 , n23 );
buf ( n1044 , n203 );
buf ( n1045 , n335 );
buf ( n1046 , n252 );
buf ( n1047 , n127 );
buf ( n1048 , n124 );
buf ( n1049 , n435 );
buf ( n1050 , n158 );
buf ( n1051 , n276 );
buf ( n1052 , n156 );
buf ( n1053 , n474 );
buf ( n1054 , n388 );
buf ( n1055 , n257 );
buf ( n1056 , n209 );
buf ( n1057 , n204 );
buf ( n1058 , n217 );
buf ( n1059 , n25 );
buf ( n1060 , n337 );
buf ( n1061 , n3 );
buf ( n1062 , n432 );
buf ( n1063 , n415 );
buf ( n1064 , n459 );
buf ( n1065 , n228 );
buf ( n1066 , n472 );
buf ( n1067 , n147 );
buf ( n1068 , n342 );
buf ( n1069 , n333 );
buf ( n1070 , n270 );
buf ( n1071 , n201 );
buf ( n1072 , n28 );
buf ( n1073 , n155 );
buf ( n1074 , n114 );
buf ( n1075 , n401 );
buf ( n1076 , n338 );
buf ( n1077 , n419 );
buf ( n1078 , n251 );
buf ( n1079 , n458 );
buf ( n1080 , n414 );
buf ( n1081 , n133 );
buf ( n1082 , n407 );
buf ( n1083 , n215 );
buf ( n1084 , n399 );
buf ( n1085 , n40 );
buf ( n1086 , n403 );
buf ( n1087 , n265 );
buf ( n1088 , n76 );
buf ( n1089 , n96 );
buf ( n1090 , n165 );
buf ( n1091 , n151 );
buf ( n1092 , n320 );
buf ( n1093 , n150 );
buf ( n1094 , n42 );
buf ( n1095 , n447 );
buf ( n1096 , n352 );
buf ( n1097 , n17 );
buf ( n1098 , n461 );
buf ( n1099 , n81 );
buf ( n1100 , n346 );
buf ( n1101 , n285 );
buf ( n1102 , n341 );
buf ( n1103 , n487 );
buf ( n1104 , n308 );
buf ( n1105 , n16 );
buf ( n1106 , n121 );
buf ( n1107 , n375 );
buf ( n1108 , n400 );
buf ( n1109 , n446 );
buf ( n1110 , n50 );
buf ( n1111 , n59 );
buf ( n1112 , n98 );
buf ( n1113 , n421 );
buf ( n1114 , n505 );
buf ( n1115 , n488 );
buf ( n1116 , n454 );
buf ( n1117 , n259 );
buf ( n1118 , n148 );
buf ( n1119 , n166 );
buf ( n1120 , n370 );
buf ( n1121 , n326 );
buf ( n1122 , n317 );
buf ( n1123 , n425 );
buf ( n1124 , n188 );
buf ( n1125 , n267 );
buf ( n1126 , n85 );
buf ( n1127 , n227 );
buf ( n1128 , n360 );
buf ( n1129 , n385 );
buf ( n1130 , n218 );
buf ( n1131 , n345 );
buf ( n1132 , n119 );
buf ( n1133 , n327 );
buf ( n1134 , n36 );
buf ( n1135 , n138 );
buf ( n1136 , n371 );
buf ( n1137 , n210 );
buf ( n1138 , n469 );
buf ( n1139 , n193 );
buf ( n1140 , n64 );
buf ( n1141 , n316 );
buf ( n1142 , n103 );
buf ( n1143 , n154 );
buf ( n1144 , n495 );
buf ( n1145 , n355 );
buf ( n1146 , n236 );
buf ( n1147 , n69 );
buf ( n1148 , n329 );
buf ( n1149 , n384 );
buf ( n1150 , n245 );
buf ( n1151 , n483 );
buf ( n1152 , n373 );
buf ( n1153 , n467 );
buf ( n1154 , n485 );
buf ( n1155 , n168 );
buf ( n1156 , n428 );
buf ( n1157 , n288 );
buf ( n1158 , n475 );
buf ( n1159 , n184 );
buf ( n1160 , n164 );
buf ( n1161 , n309 );
buf ( n1162 , n240 );
buf ( n1163 , n264 );
buf ( n1164 , n0 );
buf ( n1165 , n490 );
buf ( n1166 , n13 );
buf ( n1167 , n125 );
buf ( n1168 , n420 );
buf ( n1169 , n139 );
buf ( n1170 , n113 );
buf ( n1171 , n160 );
buf ( n1172 , n492 );
buf ( n1173 , n176 );
buf ( n1174 , n398 );
buf ( n1175 , n496 );
buf ( n1176 , n79 );
buf ( n1177 , n61 );
buf ( n1178 , n412 );
buf ( n1179 , n444 );
buf ( n1180 , n476 );
buf ( n1181 , n43 );
buf ( n1182 , n304 );
buf ( n1183 , n12 );
buf ( n1184 , n299 );
buf ( n1185 , n260 );
buf ( n1186 , n357 );
buf ( n1187 , n292 );
buf ( n1188 , n54 );
buf ( n1189 , n429 );
buf ( n1190 , n301 );
buf ( n1191 , n136 );
buf ( n1192 , n282 );
buf ( n1193 , n510 );
buf ( n1194 , n508 );
buf ( n1195 , n438 );
buf ( n1196 , n501 );
buf ( n1197 , n499 );
buf ( n1198 , n293 );
buf ( n1199 , n281 );
buf ( n1200 , n239 );
buf ( n1201 , n468 );
buf ( n1202 , n170 );
buf ( n1203 , n55 );
buf ( n1204 , n464 );
buf ( n1205 , n318 );
buf ( n1206 , n153 );
buf ( n1207 , n161 );
buf ( n1208 , n343 );
buf ( n1209 , n45 );
buf ( n1210 , n427 );
buf ( n1211 , n186 );
buf ( n1212 , n75 );
buf ( n1213 , n394 );
buf ( n1214 , n319 );
buf ( n1215 , n365 );
buf ( n1216 , n406 );
buf ( n1217 , n417 );
buf ( n1218 , n135 );
buf ( n1219 , n46 );
buf ( n1220 , n323 );
buf ( n1221 , n33 );
buf ( n1222 , n26 );
buf ( n1223 , n256 );
buf ( n1224 , n248 );
buf ( n1225 , n500 );
buf ( n1226 , n185 );
buf ( n1227 , n233 );
buf ( n1228 , n137 );
buf ( n1229 , n387 );
buf ( n1230 , n72 );
buf ( n1231 , n167 );
buf ( n1232 , n269 );
buf ( n1233 , n405 );
buf ( n1234 , n354 );
buf ( n1235 , n90 );
buf ( n1236 , n111 );
buf ( n1237 , n295 );
buf ( n1238 , n53 );
buf ( n1239 , n241 );
buf ( n1240 , n141 );
buf ( n1241 , n32 );
buf ( n1242 , n440 );
buf ( n1243 , n63 );
buf ( n1244 , n325 );
buf ( n1245 , n68 );
buf ( n1246 , n367 );
buf ( n1247 , n220 );
buf ( n1248 , n208 );
buf ( n1249 , n258 );
buf ( n1250 , n284 );
buf ( n1251 , n213 );
buf ( n1252 , n416 );
buf ( n1253 , n163 );
buf ( n1254 , n348 );
buf ( n1255 , n30 );
buf ( n1256 , n381 );
buf ( n1257 , n249 );
buf ( n1258 , n142 );
buf ( n1259 , n9 );
buf ( n1260 , n242 );
buf ( n1261 , n392 );
buf ( n1262 , n408 );
buf ( n1263 , n272 );
buf ( n1264 , n38 );
buf ( n1265 , n312 );
buf ( n1266 , n92 );
buf ( n1267 , n489 );
buf ( n1268 , n196 );
buf ( n1269 , n253 );
buf ( n1270 , n291 );
buf ( n1271 , n306 );
buf ( n1272 , n455 );
buf ( n1273 , n149 );
buf ( n1274 , n361 );
buf ( n1275 , n83 );
buf ( n1276 , n102 );
buf ( n1277 , n441 );
buf ( n1278 , n497 );
buf ( n1279 , n99 );
buf ( n1280 , n192 );
buf ( n1281 , n443 );
buf ( n1282 , n177 );
buf ( n1283 , n122 );
buf ( n1284 , n378 );
buf ( n1285 , n509 );
buf ( n1286 , n145 );
buf ( n1287 , n511 );
buf ( n1288 , n277 );
buf ( n1289 , n198 );
buf ( n1290 , n87 );
buf ( n1291 , n101 );
buf ( n1292 , n332 );
buf ( n1293 , n238 );
buf ( n1294 , n307 );
buf ( n1295 , n391 );
buf ( n1296 , n351 );
buf ( n1297 , n200 );
buf ( n1298 , n462 );
buf ( n1299 , n181 );
buf ( n1300 , n411 );
buf ( n1301 , n10 );
buf ( n1302 , n20 );
buf ( n1303 , n237 );
buf ( n1304 , n216 );
buf ( n1305 , n132 );
buf ( n1306 , n465 );
buf ( n1307 , n104 );
buf ( n1308 , n449 );
buf ( n1309 , n274 );
buf ( n1310 , n356 );
buf ( n1311 , n73 );
buf ( n1312 , n115 );
buf ( n1313 , n169 );
buf ( n1314 , n51 );
buf ( n1315 , n305 );
buf ( n1316 , n100 );
buf ( n1317 , n479 );
buf ( n1318 , n377 );
buf ( n1319 , n456 );
buf ( n1320 , n437 );
buf ( n1321 , n224 );
buf ( n1322 , n182 );
buf ( n1323 , n362 );
buf ( n1324 , n179 );
buf ( n1325 , n66 );
buf ( n1326 , n254 );
buf ( n1327 , n117 );
buf ( n1328 , n347 );
buf ( n1329 , n222 );
buf ( n1330 , n266 );
buf ( n1331 , n157 );
buf ( n1332 , n290 );
buf ( n1333 , n402 );
buf ( n1334 , n359 );
buf ( n1335 , n24 );
buf ( n1336 , n19 );
buf ( n1337 , n262 );
buf ( n1338 , n97 );
buf ( n1339 , n108 );
buf ( n1340 , n48 );
buf ( n1341 , n350 );
buf ( n1342 , n162 );
buf ( n1343 , n128 );
buf ( n1344 , n436 );
buf ( n1345 , n60 );
buf ( n1346 , n175 );
buf ( n1347 , n382 );
buf ( n1348 , n34 );
buf ( n1349 , n413 );
buf ( n1350 , n470 );
buf ( n1351 , n390 );
buf ( n1352 , n8 );
buf ( n1353 , n383 );
buf ( n1354 , n280 );
buf ( n1355 , n1 );
buf ( n1356 , n334 );
buf ( n1357 , n255 );
buf ( n1358 , n67 );
buf ( n1359 , n4 );
buf ( n1360 , n273 );
buf ( n1361 , n278 );
buf ( n1362 , n322 );
buf ( n1363 , n70 );
buf ( n1364 , n453 );
buf ( n1365 , n297 );
buf ( n1366 , n279 );
buf ( n1367 , n144 );
buf ( n1368 , n225 );
buf ( n1369 , n21 );
buf ( n1370 , n29 );
buf ( n1371 , n105 );
buf ( n1372 , n263 );
buf ( n1373 , n380 );
buf ( n1374 , n302 );
buf ( n1375 , n477 );
buf ( n1376 , n74 );
buf ( n1377 , n18 );
buf ( n1378 , n2 );
buf ( n1379 , n116 );
buf ( n1380 , n106 );
buf ( n1381 , n211 );
buf ( n1382 , n31 );
buf ( n1383 , n130 );
buf ( n1384 , n275 );
buf ( n1385 , n120 );
buf ( n1386 , n199 );
buf ( n1387 , n466 );
buf ( n1388 , n503 );
buf ( n1389 , n143 );
buf ( n1390 , n212 );
buf ( n1391 , n298 );
buf ( n1392 , n460 );
buf ( n1393 , n77 );
buf ( n1394 , n506 );
buf ( n1395 , n39 );
buf ( n1396 , n58 );
buf ( n1397 , n174 );
buf ( n1398 , n129 );
buf ( n1399 , n314 );
buf ( n1400 , n71 );
buf ( n1401 , n109 );
buf ( n1402 , n404 );
buf ( n1403 , n47 );
buf ( n1404 , n422 );
buf ( n1405 , n313 );
buf ( n1406 , n431 );
buf ( n1407 , n324 );
buf ( n1408 , n80 );
buf ( n1409 , n7 );
buf ( n1410 , n95 );
buf ( n1411 , n271 );
buf ( n1412 , n250 );
buf ( n1413 , n336 );
buf ( n1414 , n56 );
buf ( n1415 , n190 );
buf ( n1416 , n439 );
buf ( n1417 , n393 );
buf ( n1418 , n423 );
buf ( n1419 , n300 );
buf ( n1420 , n146 );
buf ( n1421 , n374 );
buf ( n1422 , n52 );
buf ( n1423 , n134 );
buf ( n1424 , n183 );
buf ( n1425 , n172 );
buf ( n1426 , n206 );
buf ( n1427 , n498 );
buf ( n1428 , n448 );
buf ( n1429 , n395 );
buf ( n1430 , n397 );
buf ( n1431 , n389 );
buf ( n1432 , n246 );
buf ( n1433 , n235 );
buf ( n1434 , n219 );
buf ( n1435 , n223 );
buf ( n1436 , n303 );
buf ( n1437 , n434 );
buf ( n1438 , n502 );
buf ( n1439 , n6 );
buf ( n1440 , n315 );
buf ( n1441 , n283 );
buf ( n1442 , n62 );
buf ( n1443 , n386 );
buf ( n1444 , n214 );
buf ( n1445 , n178 );
buf ( n1446 , n15 );
buf ( n1447 , n328 );
buf ( n1448 , n287 );
buf ( n1449 , n234 );
buf ( n1450 , n473 );
buf ( n1451 , n88 );
buf ( n1452 , n491 );
buf ( n1453 , n202 );
buf ( n1454 , n159 );
buf ( n1455 , n91 );
buf ( n1456 , n207 );
buf ( n1457 , n409 );
buf ( n1458 , n37 );
buf ( n1459 , n118 );
buf ( n1460 , n478 );
buf ( n1461 , n152 );
buf ( n1462 , n442 );
buf ( n1463 , n171 );
buf ( n1464 , n244 );
buf ( n1465 , n11 );
buf ( n1466 , n221 );
buf ( n1467 , n430 );
buf ( n1468 , n331 );
buf ( n1469 , n123 );
buf ( n1470 , n344 );
buf ( n1471 , n426 );
buf ( n1472 , n376 );
buf ( n1473 , n195 );
buf ( n1474 , n450 );
buf ( n1475 , n187 );
buf ( n1476 , n286 );
buf ( n1477 , n57 );
buf ( n1478 , n232 );
buf ( n1479 , n247 );
buf ( n1480 , n268 );
buf ( n1481 , n364 );
buf ( n1482 , n231 );
buf ( n1483 , n44 );
buf ( n1484 , n349 );
buf ( n1485 , n5 );
buf ( n1486 , n494 );
buf ( n1487 , n82 );
buf ( n1488 , n504 );
buf ( n1489 , n433 );
buf ( n1490 , n493 );
buf ( n1491 , n14 );
buf ( n1492 , n229 );
buf ( n1493 , n65 );
buf ( n1494 , n296 );
buf ( n1495 , n358 );
buf ( n1496 , n451 );
buf ( n1497 , n481 );
buf ( n1498 , n372 );
buf ( n1499 , n482 );
buf ( n1500 , n140 );
buf ( n1501 , n294 );
buf ( n1502 , n112 );
buf ( n1503 , n366 );
buf ( n1504 , n84 );
buf ( n1505 , n310 );
buf ( n1506 , n94 );
buf ( n1507 , n197 );
buf ( n1508 , n189 );
buf ( n1509 , n27 );
buf ( n1510 , n339 );
buf ( n1511 , n330 );
buf ( n1512 , n107 );
buf ( n1513 , n410 );
buf ( n1514 , n22 );
buf ( n1515 , n230 );
buf ( n1516 , n93 );
buf ( n1517 , n86 );
buf ( n1518 , n480 );
buf ( n1519 , n368 );
buf ( n1520 , n486 );
buf ( n1521 , n457 );
buf ( n1522 , n379 );
buf ( n1523 , n311 );
buf ( n1524 , n463 );
buf ( n1525 , n89 );
buf ( n1526 , n205 );
buf ( n1527 , n191 );
buf ( n1528 , n321 );
buf ( n1529 , n452 );
buf ( n1530 , n396 );
buf ( n1531 , n180 );
buf ( n1532 , n41 );
buf ( n1533 , n126 );
buf ( n1534 , n194 );
buf ( n1535 , n471 );
buf ( n1536 , n363 );
buf ( n1537 , n289 );
buf ( n1538 , n131 );
buf ( n1539 , n484 );
buf ( n1540 , n353 );
buf ( n1541 , n507 );
buf ( n1542 , n78 );
buf ( n1543 , n445 );
buf ( n1544 , n243 );
buf ( n1545 , n173 );
buf ( n1546 , n261 );
buf ( n1547 , n226 );
xor ( n1548 , n1036 , n1164 );
buf ( n1549 , n1548 );
xor ( n1550 , n1292 , n1420 );
buf ( n1551 , n1550 );
xor ( n1552 , n1549 , n1551 );
xor ( n1553 , n1037 , n1165 );
buf ( n1554 , n1553 );
xor ( n1555 , n1293 , n1421 );
buf ( n1556 , n1555 );
xor ( n1557 , n1554 , n1556 );
or ( n1558 , n1552 , n1557 );
xor ( n1559 , n1038 , n1166 );
buf ( n1560 , n1559 );
xor ( n1561 , n1294 , n1422 );
buf ( n1562 , n1561 );
xor ( n1563 , n1560 , n1562 );
or ( n1564 , n1558 , n1563 );
xor ( n1565 , n1039 , n1167 );
buf ( n1566 , n1565 );
xor ( n1567 , n1295 , n1423 );
buf ( n1568 , n1567 );
xor ( n1569 , n1566 , n1568 );
or ( n1570 , n1564 , n1569 );
xor ( n1571 , n1040 , n1168 );
buf ( n1572 , n1571 );
xor ( n1573 , n1296 , n1424 );
buf ( n1574 , n1573 );
xor ( n1575 , n1572 , n1574 );
or ( n1576 , n1570 , n1575 );
xor ( n1577 , n1041 , n1169 );
buf ( n1578 , n1577 );
xor ( n1579 , n1297 , n1425 );
buf ( n1580 , n1579 );
xor ( n1581 , n1578 , n1580 );
or ( n1582 , n1576 , n1581 );
xor ( n1583 , n1042 , n1170 );
buf ( n1584 , n1583 );
xor ( n1585 , n1298 , n1426 );
buf ( n1586 , n1585 );
xor ( n1587 , n1584 , n1586 );
or ( n1588 , n1582 , n1587 );
xor ( n1589 , n1043 , n1171 );
buf ( n1590 , n1589 );
xor ( n1591 , n1299 , n1427 );
buf ( n1592 , n1591 );
xor ( n1593 , n1590 , n1592 );
or ( n1594 , n1588 , n1593 );
xor ( n1595 , n1044 , n1172 );
buf ( n1596 , n1595 );
xor ( n1597 , n1300 , n1428 );
buf ( n1598 , n1597 );
xor ( n1599 , n1596 , n1598 );
or ( n1600 , n1594 , n1599 );
xor ( n1601 , n1045 , n1173 );
buf ( n1602 , n1601 );
xor ( n1603 , n1301 , n1429 );
buf ( n1604 , n1603 );
xor ( n1605 , n1602 , n1604 );
or ( n1606 , n1600 , n1605 );
xor ( n1607 , n1046 , n1174 );
buf ( n1608 , n1607 );
xor ( n1609 , n1302 , n1430 );
buf ( n1610 , n1609 );
xor ( n1611 , n1608 , n1610 );
or ( n1612 , n1606 , n1611 );
xor ( n1613 , n1047 , n1175 );
buf ( n1614 , n1613 );
xor ( n1615 , n1303 , n1431 );
buf ( n1616 , n1615 );
xor ( n1617 , n1614 , n1616 );
or ( n1618 , n1612 , n1617 );
xor ( n1619 , n1048 , n1176 );
buf ( n1620 , n1619 );
xor ( n1621 , n1304 , n1432 );
buf ( n1622 , n1621 );
xor ( n1623 , n1620 , n1622 );
or ( n1624 , n1618 , n1623 );
xor ( n1625 , n1049 , n1177 );
buf ( n1626 , n1625 );
xor ( n1627 , n1305 , n1433 );
buf ( n1628 , n1627 );
xor ( n1629 , n1626 , n1628 );
or ( n1630 , n1624 , n1629 );
xor ( n1631 , n1050 , n1178 );
buf ( n1632 , n1631 );
xor ( n1633 , n1306 , n1434 );
buf ( n1634 , n1633 );
xor ( n1635 , n1632 , n1634 );
or ( n1636 , n1630 , n1635 );
xor ( n1637 , n1051 , n1179 );
buf ( n1638 , n1637 );
xor ( n1639 , n1307 , n1435 );
buf ( n1640 , n1639 );
xor ( n1641 , n1638 , n1640 );
or ( n1642 , n1636 , n1641 );
xor ( n1643 , n1052 , n1180 );
buf ( n1644 , n1643 );
xor ( n1645 , n1308 , n1436 );
buf ( n1646 , n1645 );
xor ( n1647 , n1644 , n1646 );
or ( n1648 , n1642 , n1647 );
xor ( n1649 , n1053 , n1181 );
buf ( n1650 , n1649 );
xor ( n1651 , n1309 , n1437 );
buf ( n1652 , n1651 );
xor ( n1653 , n1650 , n1652 );
or ( n1654 , n1648 , n1653 );
xor ( n1655 , n1054 , n1182 );
buf ( n1656 , n1655 );
xor ( n1657 , n1310 , n1438 );
buf ( n1658 , n1657 );
xor ( n1659 , n1656 , n1658 );
or ( n1660 , n1654 , n1659 );
xor ( n1661 , n1055 , n1183 );
buf ( n1662 , n1661 );
xor ( n1663 , n1311 , n1439 );
buf ( n1664 , n1663 );
xor ( n1665 , n1662 , n1664 );
or ( n1666 , n1660 , n1665 );
xor ( n1667 , n1056 , n1184 );
buf ( n1668 , n1667 );
xor ( n1669 , n1312 , n1440 );
buf ( n1670 , n1669 );
xor ( n1671 , n1668 , n1670 );
or ( n1672 , n1666 , n1671 );
xor ( n1673 , n1057 , n1185 );
buf ( n1674 , n1673 );
xor ( n1675 , n1313 , n1441 );
buf ( n1676 , n1675 );
xor ( n1677 , n1674 , n1676 );
or ( n1678 , n1672 , n1677 );
xor ( n1679 , n1058 , n1186 );
buf ( n1680 , n1679 );
xor ( n1681 , n1314 , n1442 );
buf ( n1682 , n1681 );
xor ( n1683 , n1680 , n1682 );
or ( n1684 , n1678 , n1683 );
xor ( n1685 , n1059 , n1187 );
buf ( n1686 , n1685 );
xor ( n1687 , n1315 , n1443 );
buf ( n1688 , n1687 );
xor ( n1689 , n1686 , n1688 );
or ( n1690 , n1684 , n1689 );
xor ( n1691 , n1060 , n1188 );
buf ( n1692 , n1691 );
xor ( n1693 , n1316 , n1444 );
buf ( n1694 , n1693 );
xor ( n1695 , n1692 , n1694 );
or ( n1696 , n1690 , n1695 );
xor ( n1697 , n1061 , n1189 );
buf ( n1698 , n1697 );
xor ( n1699 , n1317 , n1445 );
buf ( n1700 , n1699 );
xor ( n1701 , n1698 , n1700 );
or ( n1702 , n1696 , n1701 );
xor ( n1703 , n1062 , n1190 );
buf ( n1704 , n1703 );
xor ( n1705 , n1318 , n1446 );
buf ( n1706 , n1705 );
xor ( n1707 , n1704 , n1706 );
or ( n1708 , n1702 , n1707 );
xor ( n1709 , n1063 , n1191 );
buf ( n1710 , n1709 );
xor ( n1711 , n1319 , n1447 );
buf ( n1712 , n1711 );
xor ( n1713 , n1710 , n1712 );
or ( n1714 , n1708 , n1713 );
xor ( n1715 , n1064 , n1192 );
buf ( n1716 , n1715 );
xor ( n1717 , n1320 , n1448 );
buf ( n1718 , n1717 );
xor ( n1719 , n1716 , n1718 );
or ( n1720 , n1714 , n1719 );
xor ( n1721 , n1065 , n1193 );
buf ( n1722 , n1721 );
xor ( n1723 , n1321 , n1449 );
buf ( n1724 , n1723 );
xor ( n1725 , n1722 , n1724 );
or ( n1726 , n1720 , n1725 );
xor ( n1727 , n1066 , n1194 );
buf ( n1728 , n1727 );
xor ( n1729 , n1322 , n1450 );
buf ( n1730 , n1729 );
xor ( n1731 , n1728 , n1730 );
or ( n1732 , n1726 , n1731 );
xor ( n1733 , n1067 , n1195 );
buf ( n1734 , n1733 );
xor ( n1735 , n1323 , n1451 );
buf ( n1736 , n1735 );
xor ( n1737 , n1734 , n1736 );
or ( n1738 , n1732 , n1737 );
xor ( n1739 , n1068 , n1196 );
buf ( n1740 , n1739 );
xor ( n1741 , n1324 , n1452 );
buf ( n1742 , n1741 );
xor ( n1743 , n1740 , n1742 );
or ( n1744 , n1738 , n1743 );
xor ( n1745 , n1069 , n1197 );
buf ( n1746 , n1745 );
xor ( n1747 , n1325 , n1453 );
buf ( n1748 , n1747 );
xor ( n1749 , n1746 , n1748 );
or ( n1750 , n1744 , n1749 );
xor ( n1751 , n1070 , n1198 );
buf ( n1752 , n1751 );
xor ( n1753 , n1326 , n1454 );
buf ( n1754 , n1753 );
xor ( n1755 , n1752 , n1754 );
or ( n1756 , n1750 , n1755 );
xor ( n1757 , n1071 , n1199 );
buf ( n1758 , n1757 );
xor ( n1759 , n1327 , n1455 );
buf ( n1760 , n1759 );
xor ( n1761 , n1758 , n1760 );
or ( n1762 , n1756 , n1761 );
xor ( n1763 , n1072 , n1200 );
buf ( n1764 , n1763 );
xor ( n1765 , n1328 , n1456 );
buf ( n1766 , n1765 );
xor ( n1767 , n1764 , n1766 );
or ( n1768 , n1762 , n1767 );
xor ( n1769 , n1073 , n1201 );
buf ( n1770 , n1769 );
xor ( n1771 , n1329 , n1457 );
buf ( n1772 , n1771 );
xor ( n1773 , n1770 , n1772 );
or ( n1774 , n1768 , n1773 );
xor ( n1775 , n1074 , n1202 );
buf ( n1776 , n1775 );
xor ( n1777 , n1330 , n1458 );
buf ( n1778 , n1777 );
xor ( n1779 , n1776 , n1778 );
or ( n1780 , n1774 , n1779 );
xor ( n1781 , n1075 , n1203 );
buf ( n1782 , n1781 );
xor ( n1783 , n1331 , n1459 );
buf ( n1784 , n1783 );
xor ( n1785 , n1782 , n1784 );
or ( n1786 , n1780 , n1785 );
xor ( n1787 , n1076 , n1204 );
buf ( n1788 , n1787 );
xor ( n1789 , n1332 , n1460 );
buf ( n1790 , n1789 );
xor ( n1791 , n1788 , n1790 );
or ( n1792 , n1786 , n1791 );
xor ( n1793 , n1077 , n1205 );
buf ( n1794 , n1793 );
xor ( n1795 , n1333 , n1461 );
buf ( n1796 , n1795 );
xor ( n1797 , n1794 , n1796 );
or ( n1798 , n1792 , n1797 );
xor ( n1799 , n1078 , n1206 );
buf ( n1800 , n1799 );
xor ( n1801 , n1334 , n1462 );
buf ( n1802 , n1801 );
xor ( n1803 , n1800 , n1802 );
or ( n1804 , n1798 , n1803 );
xor ( n1805 , n1079 , n1207 );
buf ( n1806 , n1805 );
xor ( n1807 , n1335 , n1463 );
buf ( n1808 , n1807 );
xor ( n1809 , n1806 , n1808 );
or ( n1810 , n1804 , n1809 );
xor ( n1811 , n1080 , n1208 );
buf ( n1812 , n1811 );
xor ( n1813 , n1336 , n1464 );
buf ( n1814 , n1813 );
xor ( n1815 , n1812 , n1814 );
or ( n1816 , n1810 , n1815 );
xor ( n1817 , n1081 , n1209 );
buf ( n1818 , n1817 );
xor ( n1819 , n1337 , n1465 );
buf ( n1820 , n1819 );
xor ( n1821 , n1818 , n1820 );
or ( n1822 , n1816 , n1821 );
xor ( n1823 , n1082 , n1210 );
buf ( n1824 , n1823 );
xor ( n1825 , n1338 , n1466 );
buf ( n1826 , n1825 );
xor ( n1827 , n1824 , n1826 );
or ( n1828 , n1822 , n1827 );
xor ( n1829 , n1083 , n1211 );
buf ( n1830 , n1829 );
xor ( n1831 , n1339 , n1467 );
buf ( n1832 , n1831 );
xor ( n1833 , n1830 , n1832 );
or ( n1834 , n1828 , n1833 );
xor ( n1835 , n1084 , n1212 );
buf ( n1836 , n1835 );
xor ( n1837 , n1340 , n1468 );
buf ( n1838 , n1837 );
xor ( n1839 , n1836 , n1838 );
or ( n1840 , n1834 , n1839 );
xor ( n1841 , n1085 , n1213 );
buf ( n1842 , n1841 );
xor ( n1843 , n1341 , n1469 );
buf ( n1844 , n1843 );
xor ( n1845 , n1842 , n1844 );
or ( n1846 , n1840 , n1845 );
xor ( n1847 , n1086 , n1214 );
buf ( n1848 , n1847 );
xor ( n1849 , n1342 , n1470 );
buf ( n1850 , n1849 );
xor ( n1851 , n1848 , n1850 );
or ( n1852 , n1846 , n1851 );
xor ( n1853 , n1087 , n1215 );
buf ( n1854 , n1853 );
xor ( n1855 , n1343 , n1471 );
buf ( n1856 , n1855 );
xor ( n1857 , n1854 , n1856 );
or ( n1858 , n1852 , n1857 );
xor ( n1859 , n1088 , n1216 );
buf ( n1860 , n1859 );
xor ( n1861 , n1344 , n1472 );
buf ( n1862 , n1861 );
xor ( n1863 , n1860 , n1862 );
or ( n1864 , n1858 , n1863 );
xor ( n1865 , n1089 , n1217 );
buf ( n1866 , n1865 );
xor ( n1867 , n1345 , n1473 );
buf ( n1868 , n1867 );
xor ( n1869 , n1866 , n1868 );
or ( n1870 , n1864 , n1869 );
xor ( n1871 , n1090 , n1218 );
buf ( n1872 , n1871 );
xor ( n1873 , n1346 , n1474 );
buf ( n1874 , n1873 );
xor ( n1875 , n1872 , n1874 );
or ( n1876 , n1870 , n1875 );
xor ( n1877 , n1091 , n1219 );
buf ( n1878 , n1877 );
xor ( n1879 , n1347 , n1475 );
buf ( n1880 , n1879 );
xor ( n1881 , n1878 , n1880 );
or ( n1882 , n1876 , n1881 );
xor ( n1883 , n1092 , n1220 );
buf ( n1884 , n1883 );
xor ( n1885 , n1348 , n1476 );
buf ( n1886 , n1885 );
xor ( n1887 , n1884 , n1886 );
or ( n1888 , n1882 , n1887 );
xor ( n1889 , n1093 , n1221 );
buf ( n1890 , n1889 );
xor ( n1891 , n1349 , n1477 );
buf ( n1892 , n1891 );
xor ( n1893 , n1890 , n1892 );
or ( n1894 , n1888 , n1893 );
xor ( n1895 , n1094 , n1222 );
buf ( n1896 , n1895 );
xor ( n1897 , n1350 , n1478 );
buf ( n1898 , n1897 );
xor ( n1899 , n1896 , n1898 );
or ( n1900 , n1894 , n1899 );
xor ( n1901 , n1095 , n1223 );
buf ( n1902 , n1901 );
xor ( n1903 , n1351 , n1479 );
buf ( n1904 , n1903 );
xor ( n1905 , n1902 , n1904 );
or ( n1906 , n1900 , n1905 );
xor ( n1907 , n1096 , n1224 );
buf ( n1908 , n1907 );
xor ( n1909 , n1352 , n1480 );
buf ( n1910 , n1909 );
xor ( n1911 , n1908 , n1910 );
or ( n1912 , n1906 , n1911 );
xor ( n1913 , n1097 , n1225 );
buf ( n1914 , n1913 );
xor ( n1915 , n1353 , n1481 );
buf ( n1916 , n1915 );
xor ( n1917 , n1914 , n1916 );
or ( n1918 , n1912 , n1917 );
xor ( n1919 , n1098 , n1226 );
buf ( n1920 , n1919 );
xor ( n1921 , n1354 , n1482 );
buf ( n1922 , n1921 );
xor ( n1923 , n1920 , n1922 );
or ( n1924 , n1918 , n1923 );
xor ( n1925 , n1099 , n1227 );
buf ( n1926 , n1925 );
xor ( n1927 , n1355 , n1483 );
buf ( n1928 , n1927 );
xor ( n1929 , n1926 , n1928 );
or ( n1930 , n1924 , n1929 );
xor ( n1931 , n1100 , n1228 );
buf ( n1932 , n1931 );
xor ( n1933 , n1356 , n1484 );
buf ( n1934 , n1933 );
xor ( n1935 , n1932 , n1934 );
or ( n1936 , n1930 , n1935 );
xor ( n1937 , n1101 , n1229 );
buf ( n1938 , n1937 );
xor ( n1939 , n1357 , n1485 );
buf ( n1940 , n1939 );
xor ( n1941 , n1938 , n1940 );
or ( n1942 , n1936 , n1941 );
xor ( n1943 , n1102 , n1230 );
buf ( n1944 , n1943 );
xor ( n1945 , n1358 , n1486 );
buf ( n1946 , n1945 );
xor ( n1947 , n1944 , n1946 );
or ( n1948 , n1942 , n1947 );
xor ( n1949 , n1103 , n1231 );
buf ( n1950 , n1949 );
xor ( n1951 , n1359 , n1487 );
buf ( n1952 , n1951 );
xor ( n1953 , n1950 , n1952 );
or ( n1954 , n1948 , n1953 );
xor ( n1955 , n1104 , n1232 );
buf ( n1956 , n1955 );
xor ( n1957 , n1360 , n1488 );
buf ( n1958 , n1957 );
xor ( n1959 , n1956 , n1958 );
or ( n1960 , n1954 , n1959 );
xor ( n1961 , n1105 , n1233 );
buf ( n1962 , n1961 );
xor ( n1963 , n1361 , n1489 );
buf ( n1964 , n1963 );
xor ( n1965 , n1962 , n1964 );
or ( n1966 , n1960 , n1965 );
xor ( n1967 , n1106 , n1234 );
buf ( n1968 , n1967 );
xor ( n1969 , n1362 , n1490 );
buf ( n1970 , n1969 );
xor ( n1971 , n1968 , n1970 );
or ( n1972 , n1966 , n1971 );
xor ( n1973 , n1107 , n1235 );
buf ( n1974 , n1973 );
xor ( n1975 , n1363 , n1491 );
buf ( n1976 , n1975 );
xor ( n1977 , n1974 , n1976 );
or ( n1978 , n1972 , n1977 );
xor ( n1979 , n1108 , n1236 );
buf ( n1980 , n1979 );
xor ( n1981 , n1364 , n1492 );
buf ( n1982 , n1981 );
xor ( n1983 , n1980 , n1982 );
or ( n1984 , n1978 , n1983 );
xor ( n1985 , n1109 , n1237 );
buf ( n1986 , n1985 );
xor ( n1987 , n1365 , n1493 );
buf ( n1988 , n1987 );
xor ( n1989 , n1986 , n1988 );
or ( n1990 , n1984 , n1989 );
xor ( n1991 , n1110 , n1238 );
buf ( n1992 , n1991 );
xor ( n1993 , n1366 , n1494 );
buf ( n1994 , n1993 );
xor ( n1995 , n1992 , n1994 );
or ( n1996 , n1990 , n1995 );
xor ( n1997 , n1111 , n1239 );
buf ( n1998 , n1997 );
xor ( n1999 , n1367 , n1495 );
buf ( n2000 , n1999 );
xor ( n2001 , n1998 , n2000 );
or ( n2002 , n1996 , n2001 );
xor ( n2003 , n1112 , n1240 );
buf ( n2004 , n2003 );
xor ( n2005 , n1368 , n1496 );
buf ( n2006 , n2005 );
xor ( n2007 , n2004 , n2006 );
or ( n2008 , n2002 , n2007 );
xor ( n2009 , n1113 , n1241 );
buf ( n2010 , n2009 );
xor ( n2011 , n1369 , n1497 );
buf ( n2012 , n2011 );
xor ( n2013 , n2010 , n2012 );
or ( n2014 , n2008 , n2013 );
xor ( n2015 , n1114 , n1242 );
buf ( n2016 , n2015 );
xor ( n2017 , n1370 , n1498 );
buf ( n2018 , n2017 );
xor ( n2019 , n2016 , n2018 );
or ( n2020 , n2014 , n2019 );
xor ( n2021 , n1115 , n1243 );
buf ( n2022 , n2021 );
xor ( n2023 , n1371 , n1499 );
buf ( n2024 , n2023 );
xor ( n2025 , n2022 , n2024 );
or ( n2026 , n2020 , n2025 );
xor ( n2027 , n1116 , n1244 );
buf ( n2028 , n2027 );
xor ( n2029 , n1372 , n1500 );
buf ( n2030 , n2029 );
xor ( n2031 , n2028 , n2030 );
or ( n2032 , n2026 , n2031 );
xor ( n2033 , n1117 , n1245 );
buf ( n2034 , n2033 );
xor ( n2035 , n1373 , n1501 );
buf ( n2036 , n2035 );
xor ( n2037 , n2034 , n2036 );
or ( n2038 , n2032 , n2037 );
xor ( n2039 , n1118 , n1246 );
buf ( n2040 , n2039 );
xor ( n2041 , n1374 , n1502 );
buf ( n2042 , n2041 );
xor ( n2043 , n2040 , n2042 );
or ( n2044 , n2038 , n2043 );
xor ( n2045 , n1119 , n1247 );
buf ( n2046 , n2045 );
xor ( n2047 , n1375 , n1503 );
buf ( n2048 , n2047 );
xor ( n2049 , n2046 , n2048 );
or ( n2050 , n2044 , n2049 );
xor ( n2051 , n1120 , n1248 );
buf ( n2052 , n2051 );
xor ( n2053 , n1376 , n1504 );
buf ( n2054 , n2053 );
xor ( n2055 , n2052 , n2054 );
or ( n2056 , n2050 , n2055 );
xor ( n2057 , n1121 , n1249 );
buf ( n2058 , n2057 );
xor ( n2059 , n1377 , n1505 );
buf ( n2060 , n2059 );
xor ( n2061 , n2058 , n2060 );
or ( n2062 , n2056 , n2061 );
xor ( n2063 , n1122 , n1250 );
buf ( n2064 , n2063 );
xor ( n2065 , n1378 , n1506 );
buf ( n2066 , n2065 );
xor ( n2067 , n2064 , n2066 );
or ( n2068 , n2062 , n2067 );
xor ( n2069 , n1123 , n1251 );
buf ( n2070 , n2069 );
xor ( n2071 , n1379 , n1507 );
buf ( n2072 , n2071 );
xor ( n2073 , n2070 , n2072 );
or ( n2074 , n2068 , n2073 );
xor ( n2075 , n1124 , n1252 );
buf ( n2076 , n2075 );
xor ( n2077 , n1380 , n1508 );
buf ( n2078 , n2077 );
xor ( n2079 , n2076 , n2078 );
or ( n2080 , n2074 , n2079 );
xor ( n2081 , n1125 , n1253 );
buf ( n2082 , n2081 );
xor ( n2083 , n1381 , n1509 );
buf ( n2084 , n2083 );
xor ( n2085 , n2082 , n2084 );
or ( n2086 , n2080 , n2085 );
xor ( n2087 , n1126 , n1254 );
buf ( n2088 , n2087 );
xor ( n2089 , n1382 , n1510 );
buf ( n2090 , n2089 );
xor ( n2091 , n2088 , n2090 );
or ( n2092 , n2086 , n2091 );
xor ( n2093 , n1127 , n1255 );
buf ( n2094 , n2093 );
xor ( n2095 , n1383 , n1511 );
buf ( n2096 , n2095 );
xor ( n2097 , n2094 , n2096 );
or ( n2098 , n2092 , n2097 );
xor ( n2099 , n1128 , n1256 );
buf ( n2100 , n2099 );
xor ( n2101 , n1384 , n1512 );
buf ( n2102 , n2101 );
xor ( n2103 , n2100 , n2102 );
or ( n2104 , n2098 , n2103 );
xor ( n2105 , n1129 , n1257 );
buf ( n2106 , n2105 );
xor ( n2107 , n1385 , n1513 );
buf ( n2108 , n2107 );
xor ( n2109 , n2106 , n2108 );
or ( n2110 , n2104 , n2109 );
xor ( n2111 , n1130 , n1258 );
buf ( n2112 , n2111 );
xor ( n2113 , n1386 , n1514 );
buf ( n2114 , n2113 );
xor ( n2115 , n2112 , n2114 );
or ( n2116 , n2110 , n2115 );
xor ( n2117 , n1131 , n1259 );
buf ( n2118 , n2117 );
xor ( n2119 , n1387 , n1515 );
buf ( n2120 , n2119 );
xor ( n2121 , n2118 , n2120 );
or ( n2122 , n2116 , n2121 );
xor ( n2123 , n1132 , n1260 );
buf ( n2124 , n2123 );
xor ( n2125 , n1388 , n1516 );
buf ( n2126 , n2125 );
xor ( n2127 , n2124 , n2126 );
or ( n2128 , n2122 , n2127 );
xor ( n2129 , n1133 , n1261 );
buf ( n2130 , n2129 );
xor ( n2131 , n1389 , n1517 );
buf ( n2132 , n2131 );
xor ( n2133 , n2130 , n2132 );
or ( n2134 , n2128 , n2133 );
xor ( n2135 , n1134 , n1262 );
buf ( n2136 , n2135 );
xor ( n2137 , n1390 , n1518 );
buf ( n2138 , n2137 );
xor ( n2139 , n2136 , n2138 );
or ( n2140 , n2134 , n2139 );
xor ( n2141 , n1135 , n1263 );
buf ( n2142 , n2141 );
xor ( n2143 , n1391 , n1519 );
buf ( n2144 , n2143 );
xor ( n2145 , n2142 , n2144 );
or ( n2146 , n2140 , n2145 );
xor ( n2147 , n1136 , n1264 );
buf ( n2148 , n2147 );
xor ( n2149 , n1392 , n1520 );
buf ( n2150 , n2149 );
xor ( n2151 , n2148 , n2150 );
or ( n2152 , n2146 , n2151 );
xor ( n2153 , n1137 , n1265 );
buf ( n2154 , n2153 );
xor ( n2155 , n1393 , n1521 );
buf ( n2156 , n2155 );
xor ( n2157 , n2154 , n2156 );
or ( n2158 , n2152 , n2157 );
xor ( n2159 , n1138 , n1266 );
buf ( n2160 , n2159 );
xor ( n2161 , n1394 , n1522 );
buf ( n2162 , n2161 );
xor ( n2163 , n2160 , n2162 );
or ( n2164 , n2158 , n2163 );
xor ( n2165 , n1139 , n1267 );
buf ( n2166 , n2165 );
xor ( n2167 , n1395 , n1523 );
buf ( n2168 , n2167 );
xor ( n2169 , n2166 , n2168 );
or ( n2170 , n2164 , n2169 );
xor ( n2171 , n1140 , n1268 );
buf ( n2172 , n2171 );
xor ( n2173 , n1396 , n1524 );
buf ( n2174 , n2173 );
xor ( n2175 , n2172 , n2174 );
or ( n2176 , n2170 , n2175 );
xor ( n2177 , n1141 , n1269 );
buf ( n2178 , n2177 );
xor ( n2179 , n1397 , n1525 );
buf ( n2180 , n2179 );
xor ( n2181 , n2178 , n2180 );
or ( n2182 , n2176 , n2181 );
xor ( n2183 , n1142 , n1270 );
buf ( n2184 , n2183 );
xor ( n2185 , n1398 , n1526 );
buf ( n2186 , n2185 );
xor ( n2187 , n2184 , n2186 );
or ( n2188 , n2182 , n2187 );
xor ( n2189 , n1143 , n1271 );
buf ( n2190 , n2189 );
xor ( n2191 , n1399 , n1527 );
buf ( n2192 , n2191 );
xor ( n2193 , n2190 , n2192 );
or ( n2194 , n2188 , n2193 );
xor ( n2195 , n1144 , n1272 );
buf ( n2196 , n2195 );
xor ( n2197 , n1400 , n1528 );
buf ( n2198 , n2197 );
xor ( n2199 , n2196 , n2198 );
or ( n2200 , n2194 , n2199 );
xor ( n2201 , n1145 , n1273 );
buf ( n2202 , n2201 );
xor ( n2203 , n1401 , n1529 );
buf ( n2204 , n2203 );
xor ( n2205 , n2202 , n2204 );
or ( n2206 , n2200 , n2205 );
xor ( n2207 , n1146 , n1274 );
buf ( n2208 , n2207 );
xor ( n2209 , n1402 , n1530 );
buf ( n2210 , n2209 );
xor ( n2211 , n2208 , n2210 );
or ( n2212 , n2206 , n2211 );
xor ( n2213 , n1147 , n1275 );
buf ( n2214 , n2213 );
xor ( n2215 , n1403 , n1531 );
buf ( n2216 , n2215 );
xor ( n2217 , n2214 , n2216 );
or ( n2218 , n2212 , n2217 );
xor ( n2219 , n1148 , n1276 );
buf ( n2220 , n2219 );
xor ( n2221 , n1404 , n1532 );
buf ( n2222 , n2221 );
xor ( n2223 , n2220 , n2222 );
or ( n2224 , n2218 , n2223 );
xor ( n2225 , n1149 , n1277 );
buf ( n2226 , n2225 );
xor ( n2227 , n1405 , n1533 );
buf ( n2228 , n2227 );
xor ( n2229 , n2226 , n2228 );
or ( n2230 , n2224 , n2229 );
xor ( n2231 , n1150 , n1278 );
buf ( n2232 , n2231 );
xor ( n2233 , n1406 , n1534 );
buf ( n2234 , n2233 );
xor ( n2235 , n2232 , n2234 );
or ( n2236 , n2230 , n2235 );
xor ( n2237 , n1151 , n1279 );
buf ( n2238 , n2237 );
xor ( n2239 , n1407 , n1535 );
buf ( n2240 , n2239 );
xor ( n2241 , n2238 , n2240 );
or ( n2242 , n2236 , n2241 );
xor ( n2243 , n1152 , n1280 );
buf ( n2244 , n2243 );
xor ( n2245 , n1408 , n1536 );
buf ( n2246 , n2245 );
xor ( n2247 , n2244 , n2246 );
or ( n2248 , n2242 , n2247 );
xor ( n2249 , n1153 , n1281 );
buf ( n2250 , n2249 );
xor ( n2251 , n1409 , n1537 );
buf ( n2252 , n2251 );
xor ( n2253 , n2250 , n2252 );
or ( n2254 , n2248 , n2253 );
xor ( n2255 , n1154 , n1282 );
buf ( n2256 , n2255 );
xor ( n2257 , n1410 , n1538 );
buf ( n2258 , n2257 );
xor ( n2259 , n2256 , n2258 );
or ( n2260 , n2254 , n2259 );
xor ( n2261 , n1155 , n1283 );
buf ( n2262 , n2261 );
xor ( n2263 , n1411 , n1539 );
buf ( n2264 , n2263 );
xor ( n2265 , n2262 , n2264 );
or ( n2266 , n2260 , n2265 );
xor ( n2267 , n1156 , n1284 );
buf ( n2268 , n2267 );
xor ( n2269 , n1412 , n1540 );
buf ( n2270 , n2269 );
xor ( n2271 , n2268 , n2270 );
or ( n2272 , n2266 , n2271 );
xor ( n2273 , n1157 , n1285 );
buf ( n2274 , n2273 );
xor ( n2275 , n1413 , n1541 );
buf ( n2276 , n2275 );
xor ( n2277 , n2274 , n2276 );
or ( n2278 , n2272 , n2277 );
xor ( n2279 , n1158 , n1286 );
buf ( n2280 , n2279 );
xor ( n2281 , n1414 , n1542 );
buf ( n2282 , n2281 );
xor ( n2283 , n2280 , n2282 );
or ( n2284 , n2278 , n2283 );
xor ( n2285 , n1159 , n1287 );
buf ( n2286 , n2285 );
xor ( n2287 , n1415 , n1543 );
buf ( n2288 , n2287 );
xor ( n2289 , n2286 , n2288 );
or ( n2290 , n2284 , n2289 );
xor ( n2291 , n1160 , n1288 );
buf ( n2292 , n2291 );
xor ( n2293 , n1416 , n1544 );
buf ( n2294 , n2293 );
xor ( n2295 , n2292 , n2294 );
or ( n2296 , n2290 , n2295 );
xor ( n2297 , n1161 , n1289 );
buf ( n2298 , n2297 );
xor ( n2299 , n1417 , n1545 );
buf ( n2300 , n2299 );
xor ( n2301 , n2298 , n2300 );
or ( n2302 , n2296 , n2301 );
xor ( n2303 , n1162 , n1290 );
buf ( n2304 , n2303 );
xor ( n2305 , n1418 , n1546 );
buf ( n2306 , n2305 );
xor ( n2307 , n2304 , n2306 );
or ( n2308 , n2302 , n2307 );
xor ( n2309 , n1163 , n1291 );
buf ( n2310 , n2309 );
xor ( n2311 , n1419 , n1547 );
buf ( n2312 , n2311 );
xor ( n2313 , n2310 , n2312 );
or ( n2314 , n2308 , n2313 );
not ( n2315 , n2314 );
buf ( n2316 , n2315 );
not ( n2317 , n2316 );
and ( n2318 , n2317 , n1269 );
not ( n2319 , n1406 );
and ( n2320 , n2318 , n2319 );
buf ( n2321 , n2320 );
buf ( n2322 , n2321 );
xor ( n2323 , n1036 , n1420 );
buf ( n2324 , n2323 );
xor ( n2325 , n1164 , n1292 );
buf ( n2326 , n2325 );
xor ( n2327 , n2324 , n2326 );
xor ( n2328 , n1037 , n1421 );
buf ( n2329 , n2328 );
xor ( n2330 , n1165 , n1293 );
buf ( n2331 , n2330 );
xor ( n2332 , n2329 , n2331 );
or ( n2333 , n2327 , n2332 );
xor ( n2334 , n1038 , n1422 );
buf ( n2335 , n2334 );
xor ( n2336 , n1166 , n1294 );
buf ( n2337 , n2336 );
xor ( n2338 , n2335 , n2337 );
or ( n2339 , n2333 , n2338 );
xor ( n2340 , n1039 , n1423 );
buf ( n2341 , n2340 );
xor ( n2342 , n1167 , n1295 );
buf ( n2343 , n2342 );
xor ( n2344 , n2341 , n2343 );
or ( n2345 , n2339 , n2344 );
xor ( n2346 , n1040 , n1424 );
buf ( n2347 , n2346 );
xor ( n2348 , n1168 , n1296 );
buf ( n2349 , n2348 );
xor ( n2350 , n2347 , n2349 );
or ( n2351 , n2345 , n2350 );
xor ( n2352 , n1041 , n1425 );
buf ( n2353 , n2352 );
xor ( n2354 , n1169 , n1297 );
buf ( n2355 , n2354 );
xor ( n2356 , n2353 , n2355 );
or ( n2357 , n2351 , n2356 );
xor ( n2358 , n1042 , n1426 );
buf ( n2359 , n2358 );
xor ( n2360 , n1170 , n1298 );
buf ( n2361 , n2360 );
xor ( n2362 , n2359 , n2361 );
or ( n2363 , n2357 , n2362 );
xor ( n2364 , n1043 , n1427 );
buf ( n2365 , n2364 );
xor ( n2366 , n1171 , n1299 );
buf ( n2367 , n2366 );
xor ( n2368 , n2365 , n2367 );
or ( n2369 , n2363 , n2368 );
xor ( n2370 , n1044 , n1428 );
buf ( n2371 , n2370 );
xor ( n2372 , n1172 , n1300 );
buf ( n2373 , n2372 );
xor ( n2374 , n2371 , n2373 );
or ( n2375 , n2369 , n2374 );
xor ( n2376 , n1045 , n1429 );
buf ( n2377 , n2376 );
xor ( n2378 , n1173 , n1301 );
buf ( n2379 , n2378 );
xor ( n2380 , n2377 , n2379 );
or ( n2381 , n2375 , n2380 );
xor ( n2382 , n1046 , n1430 );
buf ( n2383 , n2382 );
xor ( n2384 , n1174 , n1302 );
buf ( n2385 , n2384 );
xor ( n2386 , n2383 , n2385 );
or ( n2387 , n2381 , n2386 );
xor ( n2388 , n1047 , n1431 );
buf ( n2389 , n2388 );
xor ( n2390 , n1175 , n1303 );
buf ( n2391 , n2390 );
xor ( n2392 , n2389 , n2391 );
or ( n2393 , n2387 , n2392 );
xor ( n2394 , n1048 , n1432 );
buf ( n2395 , n2394 );
xor ( n2396 , n1176 , n1304 );
buf ( n2397 , n2396 );
xor ( n2398 , n2395 , n2397 );
or ( n2399 , n2393 , n2398 );
xor ( n2400 , n1049 , n1433 );
buf ( n2401 , n2400 );
xor ( n2402 , n1177 , n1305 );
buf ( n2403 , n2402 );
xor ( n2404 , n2401 , n2403 );
or ( n2405 , n2399 , n2404 );
xor ( n2406 , n1050 , n1434 );
buf ( n2407 , n2406 );
xor ( n2408 , n1178 , n1306 );
buf ( n2409 , n2408 );
xor ( n2410 , n2407 , n2409 );
or ( n2411 , n2405 , n2410 );
xor ( n2412 , n1051 , n1435 );
buf ( n2413 , n2412 );
xor ( n2414 , n1179 , n1307 );
buf ( n2415 , n2414 );
xor ( n2416 , n2413 , n2415 );
or ( n2417 , n2411 , n2416 );
xor ( n2418 , n1052 , n1436 );
buf ( n2419 , n2418 );
xor ( n2420 , n1180 , n1308 );
buf ( n2421 , n2420 );
xor ( n2422 , n2419 , n2421 );
or ( n2423 , n2417 , n2422 );
xor ( n2424 , n1053 , n1437 );
buf ( n2425 , n2424 );
xor ( n2426 , n1181 , n1309 );
buf ( n2427 , n2426 );
xor ( n2428 , n2425 , n2427 );
or ( n2429 , n2423 , n2428 );
xor ( n2430 , n1054 , n1438 );
buf ( n2431 , n2430 );
xor ( n2432 , n1182 , n1310 );
buf ( n2433 , n2432 );
xor ( n2434 , n2431 , n2433 );
or ( n2435 , n2429 , n2434 );
xor ( n2436 , n1055 , n1439 );
buf ( n2437 , n2436 );
xor ( n2438 , n1183 , n1311 );
buf ( n2439 , n2438 );
xor ( n2440 , n2437 , n2439 );
or ( n2441 , n2435 , n2440 );
xor ( n2442 , n1056 , n1440 );
buf ( n2443 , n2442 );
xor ( n2444 , n1184 , n1312 );
buf ( n2445 , n2444 );
xor ( n2446 , n2443 , n2445 );
or ( n2447 , n2441 , n2446 );
xor ( n2448 , n1057 , n1441 );
buf ( n2449 , n2448 );
xor ( n2450 , n1185 , n1313 );
buf ( n2451 , n2450 );
xor ( n2452 , n2449 , n2451 );
or ( n2453 , n2447 , n2452 );
xor ( n2454 , n1058 , n1442 );
buf ( n2455 , n2454 );
xor ( n2456 , n1186 , n1314 );
buf ( n2457 , n2456 );
xor ( n2458 , n2455 , n2457 );
or ( n2459 , n2453 , n2458 );
xor ( n2460 , n1059 , n1443 );
buf ( n2461 , n2460 );
xor ( n2462 , n1187 , n1315 );
buf ( n2463 , n2462 );
xor ( n2464 , n2461 , n2463 );
or ( n2465 , n2459 , n2464 );
xor ( n2466 , n1060 , n1444 );
buf ( n2467 , n2466 );
xor ( n2468 , n1188 , n1316 );
buf ( n2469 , n2468 );
xor ( n2470 , n2467 , n2469 );
or ( n2471 , n2465 , n2470 );
xor ( n2472 , n1061 , n1445 );
buf ( n2473 , n2472 );
xor ( n2474 , n1189 , n1317 );
buf ( n2475 , n2474 );
xor ( n2476 , n2473 , n2475 );
or ( n2477 , n2471 , n2476 );
xor ( n2478 , n1062 , n1446 );
buf ( n2479 , n2478 );
xor ( n2480 , n1190 , n1318 );
buf ( n2481 , n2480 );
xor ( n2482 , n2479 , n2481 );
or ( n2483 , n2477 , n2482 );
xor ( n2484 , n1063 , n1447 );
buf ( n2485 , n2484 );
xor ( n2486 , n1191 , n1319 );
buf ( n2487 , n2486 );
xor ( n2488 , n2485 , n2487 );
or ( n2489 , n2483 , n2488 );
xor ( n2490 , n1064 , n1448 );
buf ( n2491 , n2490 );
xor ( n2492 , n1192 , n1320 );
buf ( n2493 , n2492 );
xor ( n2494 , n2491 , n2493 );
or ( n2495 , n2489 , n2494 );
xor ( n2496 , n1065 , n1449 );
buf ( n2497 , n2496 );
xor ( n2498 , n1193 , n1321 );
buf ( n2499 , n2498 );
xor ( n2500 , n2497 , n2499 );
or ( n2501 , n2495 , n2500 );
xor ( n2502 , n1066 , n1450 );
buf ( n2503 , n2502 );
xor ( n2504 , n1194 , n1322 );
buf ( n2505 , n2504 );
xor ( n2506 , n2503 , n2505 );
or ( n2507 , n2501 , n2506 );
xor ( n2508 , n1067 , n1451 );
buf ( n2509 , n2508 );
xor ( n2510 , n1195 , n1323 );
buf ( n2511 , n2510 );
xor ( n2512 , n2509 , n2511 );
or ( n2513 , n2507 , n2512 );
xor ( n2514 , n1068 , n1452 );
buf ( n2515 , n2514 );
xor ( n2516 , n1196 , n1324 );
buf ( n2517 , n2516 );
xor ( n2518 , n2515 , n2517 );
or ( n2519 , n2513 , n2518 );
xor ( n2520 , n1069 , n1453 );
buf ( n2521 , n2520 );
xor ( n2522 , n1197 , n1325 );
buf ( n2523 , n2522 );
xor ( n2524 , n2521 , n2523 );
or ( n2525 , n2519 , n2524 );
xor ( n2526 , n1070 , n1454 );
buf ( n2527 , n2526 );
xor ( n2528 , n1198 , n1326 );
buf ( n2529 , n2528 );
xor ( n2530 , n2527 , n2529 );
or ( n2531 , n2525 , n2530 );
xor ( n2532 , n1071 , n1455 );
buf ( n2533 , n2532 );
xor ( n2534 , n1199 , n1327 );
buf ( n2535 , n2534 );
xor ( n2536 , n2533 , n2535 );
or ( n2537 , n2531 , n2536 );
xor ( n2538 , n1072 , n1456 );
buf ( n2539 , n2538 );
xor ( n2540 , n1200 , n1328 );
buf ( n2541 , n2540 );
xor ( n2542 , n2539 , n2541 );
or ( n2543 , n2537 , n2542 );
xor ( n2544 , n1073 , n1457 );
buf ( n2545 , n2544 );
xor ( n2546 , n1201 , n1329 );
buf ( n2547 , n2546 );
xor ( n2548 , n2545 , n2547 );
or ( n2549 , n2543 , n2548 );
xor ( n2550 , n1074 , n1458 );
buf ( n2551 , n2550 );
xor ( n2552 , n1202 , n1330 );
buf ( n2553 , n2552 );
xor ( n2554 , n2551 , n2553 );
or ( n2555 , n2549 , n2554 );
xor ( n2556 , n1075 , n1459 );
buf ( n2557 , n2556 );
xor ( n2558 , n1203 , n1331 );
buf ( n2559 , n2558 );
xor ( n2560 , n2557 , n2559 );
or ( n2561 , n2555 , n2560 );
xor ( n2562 , n1076 , n1460 );
buf ( n2563 , n2562 );
xor ( n2564 , n1204 , n1332 );
buf ( n2565 , n2564 );
xor ( n2566 , n2563 , n2565 );
or ( n2567 , n2561 , n2566 );
xor ( n2568 , n1077 , n1461 );
buf ( n2569 , n2568 );
xor ( n2570 , n1205 , n1333 );
buf ( n2571 , n2570 );
xor ( n2572 , n2569 , n2571 );
or ( n2573 , n2567 , n2572 );
xor ( n2574 , n1078 , n1462 );
buf ( n2575 , n2574 );
xor ( n2576 , n1206 , n1334 );
buf ( n2577 , n2576 );
xor ( n2578 , n2575 , n2577 );
or ( n2579 , n2573 , n2578 );
xor ( n2580 , n1079 , n1463 );
buf ( n2581 , n2580 );
xor ( n2582 , n1207 , n1335 );
buf ( n2583 , n2582 );
xor ( n2584 , n2581 , n2583 );
or ( n2585 , n2579 , n2584 );
xor ( n2586 , n1080 , n1464 );
buf ( n2587 , n2586 );
xor ( n2588 , n1208 , n1336 );
buf ( n2589 , n2588 );
xor ( n2590 , n2587 , n2589 );
or ( n2591 , n2585 , n2590 );
xor ( n2592 , n1081 , n1465 );
buf ( n2593 , n2592 );
xor ( n2594 , n1209 , n1337 );
buf ( n2595 , n2594 );
xor ( n2596 , n2593 , n2595 );
or ( n2597 , n2591 , n2596 );
xor ( n2598 , n1082 , n1466 );
buf ( n2599 , n2598 );
xor ( n2600 , n1210 , n1338 );
buf ( n2601 , n2600 );
xor ( n2602 , n2599 , n2601 );
or ( n2603 , n2597 , n2602 );
xor ( n2604 , n1083 , n1467 );
buf ( n2605 , n2604 );
xor ( n2606 , n1211 , n1339 );
buf ( n2607 , n2606 );
xor ( n2608 , n2605 , n2607 );
or ( n2609 , n2603 , n2608 );
xor ( n2610 , n1084 , n1468 );
buf ( n2611 , n2610 );
xor ( n2612 , n1212 , n1340 );
buf ( n2613 , n2612 );
xor ( n2614 , n2611 , n2613 );
or ( n2615 , n2609 , n2614 );
xor ( n2616 , n1085 , n1469 );
buf ( n2617 , n2616 );
xor ( n2618 , n1213 , n1341 );
buf ( n2619 , n2618 );
xor ( n2620 , n2617 , n2619 );
or ( n2621 , n2615 , n2620 );
xor ( n2622 , n1086 , n1470 );
buf ( n2623 , n2622 );
xor ( n2624 , n1214 , n1342 );
buf ( n2625 , n2624 );
xor ( n2626 , n2623 , n2625 );
or ( n2627 , n2621 , n2626 );
xor ( n2628 , n1087 , n1471 );
buf ( n2629 , n2628 );
xor ( n2630 , n1215 , n1343 );
buf ( n2631 , n2630 );
xor ( n2632 , n2629 , n2631 );
or ( n2633 , n2627 , n2632 );
xor ( n2634 , n1088 , n1472 );
buf ( n2635 , n2634 );
xor ( n2636 , n1216 , n1344 );
buf ( n2637 , n2636 );
xor ( n2638 , n2635 , n2637 );
or ( n2639 , n2633 , n2638 );
xor ( n2640 , n1089 , n1473 );
buf ( n2641 , n2640 );
xor ( n2642 , n1217 , n1345 );
buf ( n2643 , n2642 );
xor ( n2644 , n2641 , n2643 );
or ( n2645 , n2639 , n2644 );
xor ( n2646 , n1090 , n1474 );
buf ( n2647 , n2646 );
xor ( n2648 , n1218 , n1346 );
buf ( n2649 , n2648 );
xor ( n2650 , n2647 , n2649 );
or ( n2651 , n2645 , n2650 );
xor ( n2652 , n1091 , n1475 );
buf ( n2653 , n2652 );
xor ( n2654 , n1219 , n1347 );
buf ( n2655 , n2654 );
xor ( n2656 , n2653 , n2655 );
or ( n2657 , n2651 , n2656 );
xor ( n2658 , n1092 , n1476 );
buf ( n2659 , n2658 );
xor ( n2660 , n1220 , n1348 );
buf ( n2661 , n2660 );
xor ( n2662 , n2659 , n2661 );
or ( n2663 , n2657 , n2662 );
xor ( n2664 , n1093 , n1477 );
buf ( n2665 , n2664 );
xor ( n2666 , n1221 , n1349 );
buf ( n2667 , n2666 );
xor ( n2668 , n2665 , n2667 );
or ( n2669 , n2663 , n2668 );
xor ( n2670 , n1094 , n1478 );
buf ( n2671 , n2670 );
xor ( n2672 , n1222 , n1350 );
buf ( n2673 , n2672 );
xor ( n2674 , n2671 , n2673 );
or ( n2675 , n2669 , n2674 );
xor ( n2676 , n1095 , n1479 );
buf ( n2677 , n2676 );
xor ( n2678 , n1223 , n1351 );
buf ( n2679 , n2678 );
xor ( n2680 , n2677 , n2679 );
or ( n2681 , n2675 , n2680 );
xor ( n2682 , n1096 , n1480 );
buf ( n2683 , n2682 );
xor ( n2684 , n1224 , n1352 );
buf ( n2685 , n2684 );
xor ( n2686 , n2683 , n2685 );
or ( n2687 , n2681 , n2686 );
xor ( n2688 , n1097 , n1481 );
buf ( n2689 , n2688 );
xor ( n2690 , n1225 , n1353 );
buf ( n2691 , n2690 );
xor ( n2692 , n2689 , n2691 );
or ( n2693 , n2687 , n2692 );
xor ( n2694 , n1098 , n1482 );
buf ( n2695 , n2694 );
xor ( n2696 , n1226 , n1354 );
buf ( n2697 , n2696 );
xor ( n2698 , n2695 , n2697 );
or ( n2699 , n2693 , n2698 );
xor ( n2700 , n1099 , n1483 );
buf ( n2701 , n2700 );
xor ( n2702 , n1227 , n1355 );
buf ( n2703 , n2702 );
xor ( n2704 , n2701 , n2703 );
or ( n2705 , n2699 , n2704 );
xor ( n2706 , n1100 , n1484 );
buf ( n2707 , n2706 );
xor ( n2708 , n1228 , n1356 );
buf ( n2709 , n2708 );
xor ( n2710 , n2707 , n2709 );
or ( n2711 , n2705 , n2710 );
xor ( n2712 , n1101 , n1485 );
buf ( n2713 , n2712 );
xor ( n2714 , n1229 , n1357 );
buf ( n2715 , n2714 );
xor ( n2716 , n2713 , n2715 );
or ( n2717 , n2711 , n2716 );
xor ( n2718 , n1102 , n1486 );
buf ( n2719 , n2718 );
xor ( n2720 , n1230 , n1358 );
buf ( n2721 , n2720 );
xor ( n2722 , n2719 , n2721 );
or ( n2723 , n2717 , n2722 );
xor ( n2724 , n1103 , n1487 );
buf ( n2725 , n2724 );
xor ( n2726 , n1231 , n1359 );
buf ( n2727 , n2726 );
xor ( n2728 , n2725 , n2727 );
or ( n2729 , n2723 , n2728 );
xor ( n2730 , n1104 , n1488 );
buf ( n2731 , n2730 );
xor ( n2732 , n1232 , n1360 );
buf ( n2733 , n2732 );
xor ( n2734 , n2731 , n2733 );
or ( n2735 , n2729 , n2734 );
xor ( n2736 , n1105 , n1489 );
buf ( n2737 , n2736 );
xor ( n2738 , n1233 , n1361 );
buf ( n2739 , n2738 );
xor ( n2740 , n2737 , n2739 );
or ( n2741 , n2735 , n2740 );
xor ( n2742 , n1106 , n1490 );
buf ( n2743 , n2742 );
xor ( n2744 , n1234 , n1362 );
buf ( n2745 , n2744 );
xor ( n2746 , n2743 , n2745 );
or ( n2747 , n2741 , n2746 );
xor ( n2748 , n1107 , n1491 );
buf ( n2749 , n2748 );
xor ( n2750 , n1235 , n1363 );
buf ( n2751 , n2750 );
xor ( n2752 , n2749 , n2751 );
or ( n2753 , n2747 , n2752 );
xor ( n2754 , n1108 , n1492 );
buf ( n2755 , n2754 );
xor ( n2756 , n1236 , n1364 );
buf ( n2757 , n2756 );
xor ( n2758 , n2755 , n2757 );
or ( n2759 , n2753 , n2758 );
xor ( n2760 , n1109 , n1493 );
buf ( n2761 , n2760 );
xor ( n2762 , n1237 , n1365 );
buf ( n2763 , n2762 );
xor ( n2764 , n2761 , n2763 );
or ( n2765 , n2759 , n2764 );
xor ( n2766 , n1110 , n1494 );
buf ( n2767 , n2766 );
xor ( n2768 , n1238 , n1366 );
buf ( n2769 , n2768 );
xor ( n2770 , n2767 , n2769 );
or ( n2771 , n2765 , n2770 );
xor ( n2772 , n1111 , n1495 );
buf ( n2773 , n2772 );
xor ( n2774 , n1239 , n1367 );
buf ( n2775 , n2774 );
xor ( n2776 , n2773 , n2775 );
or ( n2777 , n2771 , n2776 );
xor ( n2778 , n1112 , n1496 );
buf ( n2779 , n2778 );
xor ( n2780 , n1240 , n1368 );
buf ( n2781 , n2780 );
xor ( n2782 , n2779 , n2781 );
or ( n2783 , n2777 , n2782 );
xor ( n2784 , n1113 , n1497 );
buf ( n2785 , n2784 );
xor ( n2786 , n1241 , n1369 );
buf ( n2787 , n2786 );
xor ( n2788 , n2785 , n2787 );
or ( n2789 , n2783 , n2788 );
xor ( n2790 , n1114 , n1498 );
buf ( n2791 , n2790 );
xor ( n2792 , n1242 , n1370 );
buf ( n2793 , n2792 );
xor ( n2794 , n2791 , n2793 );
or ( n2795 , n2789 , n2794 );
xor ( n2796 , n1115 , n1499 );
buf ( n2797 , n2796 );
xor ( n2798 , n1243 , n1371 );
buf ( n2799 , n2798 );
xor ( n2800 , n2797 , n2799 );
or ( n2801 , n2795 , n2800 );
xor ( n2802 , n1116 , n1500 );
buf ( n2803 , n2802 );
xor ( n2804 , n1244 , n1372 );
buf ( n2805 , n2804 );
xor ( n2806 , n2803 , n2805 );
or ( n2807 , n2801 , n2806 );
xor ( n2808 , n1117 , n1501 );
buf ( n2809 , n2808 );
xor ( n2810 , n1245 , n1373 );
buf ( n2811 , n2810 );
xor ( n2812 , n2809 , n2811 );
or ( n2813 , n2807 , n2812 );
xor ( n2814 , n1118 , n1502 );
buf ( n2815 , n2814 );
xor ( n2816 , n1246 , n1374 );
buf ( n2817 , n2816 );
xor ( n2818 , n2815 , n2817 );
or ( n2819 , n2813 , n2818 );
xor ( n2820 , n1119 , n1503 );
buf ( n2821 , n2820 );
xor ( n2822 , n1247 , n1375 );
buf ( n2823 , n2822 );
xor ( n2824 , n2821 , n2823 );
or ( n2825 , n2819 , n2824 );
xor ( n2826 , n1120 , n1504 );
buf ( n2827 , n2826 );
xor ( n2828 , n1248 , n1376 );
buf ( n2829 , n2828 );
xor ( n2830 , n2827 , n2829 );
or ( n2831 , n2825 , n2830 );
xor ( n2832 , n1121 , n1505 );
buf ( n2833 , n2832 );
xor ( n2834 , n1249 , n1377 );
buf ( n2835 , n2834 );
xor ( n2836 , n2833 , n2835 );
or ( n2837 , n2831 , n2836 );
xor ( n2838 , n1122 , n1506 );
buf ( n2839 , n2838 );
xor ( n2840 , n1250 , n1378 );
buf ( n2841 , n2840 );
xor ( n2842 , n2839 , n2841 );
or ( n2843 , n2837 , n2842 );
xor ( n2844 , n1123 , n1507 );
buf ( n2845 , n2844 );
xor ( n2846 , n1251 , n1379 );
buf ( n2847 , n2846 );
xor ( n2848 , n2845 , n2847 );
or ( n2849 , n2843 , n2848 );
xor ( n2850 , n1124 , n1508 );
buf ( n2851 , n2850 );
xor ( n2852 , n1252 , n1380 );
buf ( n2853 , n2852 );
xor ( n2854 , n2851 , n2853 );
or ( n2855 , n2849 , n2854 );
xor ( n2856 , n1125 , n1509 );
buf ( n2857 , n2856 );
xor ( n2858 , n1253 , n1381 );
buf ( n2859 , n2858 );
xor ( n2860 , n2857 , n2859 );
or ( n2861 , n2855 , n2860 );
xor ( n2862 , n1126 , n1510 );
buf ( n2863 , n2862 );
xor ( n2864 , n1254 , n1382 );
buf ( n2865 , n2864 );
xor ( n2866 , n2863 , n2865 );
or ( n2867 , n2861 , n2866 );
xor ( n2868 , n1127 , n1511 );
buf ( n2869 , n2868 );
xor ( n2870 , n1255 , n1383 );
buf ( n2871 , n2870 );
xor ( n2872 , n2869 , n2871 );
or ( n2873 , n2867 , n2872 );
xor ( n2874 , n1128 , n1512 );
buf ( n2875 , n2874 );
xor ( n2876 , n1256 , n1384 );
buf ( n2877 , n2876 );
xor ( n2878 , n2875 , n2877 );
or ( n2879 , n2873 , n2878 );
xor ( n2880 , n1129 , n1513 );
buf ( n2881 , n2880 );
xor ( n2882 , n1257 , n1385 );
buf ( n2883 , n2882 );
xor ( n2884 , n2881 , n2883 );
or ( n2885 , n2879 , n2884 );
xor ( n2886 , n1130 , n1514 );
buf ( n2887 , n2886 );
xor ( n2888 , n1258 , n1386 );
buf ( n2889 , n2888 );
xor ( n2890 , n2887 , n2889 );
or ( n2891 , n2885 , n2890 );
xor ( n2892 , n1131 , n1515 );
buf ( n2893 , n2892 );
xor ( n2894 , n1259 , n1387 );
buf ( n2895 , n2894 );
xor ( n2896 , n2893 , n2895 );
or ( n2897 , n2891 , n2896 );
xor ( n2898 , n1132 , n1516 );
buf ( n2899 , n2898 );
xor ( n2900 , n1260 , n1388 );
buf ( n2901 , n2900 );
xor ( n2902 , n2899 , n2901 );
or ( n2903 , n2897 , n2902 );
xor ( n2904 , n1133 , n1517 );
buf ( n2905 , n2904 );
xor ( n2906 , n1261 , n1389 );
buf ( n2907 , n2906 );
xor ( n2908 , n2905 , n2907 );
or ( n2909 , n2903 , n2908 );
xor ( n2910 , n1134 , n1518 );
buf ( n2911 , n2910 );
xor ( n2912 , n1262 , n1390 );
buf ( n2913 , n2912 );
xor ( n2914 , n2911 , n2913 );
or ( n2915 , n2909 , n2914 );
xor ( n2916 , n1135 , n1519 );
buf ( n2917 , n2916 );
xor ( n2918 , n1263 , n1391 );
buf ( n2919 , n2918 );
xor ( n2920 , n2917 , n2919 );
or ( n2921 , n2915 , n2920 );
xor ( n2922 , n1136 , n1520 );
buf ( n2923 , n2922 );
xor ( n2924 , n1264 , n1392 );
buf ( n2925 , n2924 );
xor ( n2926 , n2923 , n2925 );
or ( n2927 , n2921 , n2926 );
xor ( n2928 , n1137 , n1521 );
buf ( n2929 , n2928 );
xor ( n2930 , n1265 , n1393 );
buf ( n2931 , n2930 );
xor ( n2932 , n2929 , n2931 );
or ( n2933 , n2927 , n2932 );
xor ( n2934 , n1138 , n1522 );
buf ( n2935 , n2934 );
xor ( n2936 , n1266 , n1394 );
buf ( n2937 , n2936 );
xor ( n2938 , n2935 , n2937 );
or ( n2939 , n2933 , n2938 );
xor ( n2940 , n1139 , n1523 );
buf ( n2941 , n2940 );
xor ( n2942 , n1267 , n1395 );
buf ( n2943 , n2942 );
xor ( n2944 , n2941 , n2943 );
or ( n2945 , n2939 , n2944 );
xor ( n2946 , n1140 , n1524 );
buf ( n2947 , n2946 );
xor ( n2948 , n1268 , n1396 );
buf ( n2949 , n2948 );
xor ( n2950 , n2947 , n2949 );
or ( n2951 , n2945 , n2950 );
xor ( n2952 , n1141 , n1525 );
buf ( n2953 , n2952 );
xor ( n2954 , n1269 , n1397 );
buf ( n2955 , n2954 );
xor ( n2956 , n2953 , n2955 );
or ( n2957 , n2951 , n2956 );
xor ( n2958 , n1142 , n1526 );
buf ( n2959 , n2958 );
xor ( n2960 , n1270 , n1398 );
buf ( n2961 , n2960 );
xor ( n2962 , n2959 , n2961 );
or ( n2963 , n2957 , n2962 );
xor ( n2964 , n1143 , n1527 );
buf ( n2965 , n2964 );
xor ( n2966 , n1271 , n1399 );
buf ( n2967 , n2966 );
xor ( n2968 , n2965 , n2967 );
or ( n2969 , n2963 , n2968 );
xor ( n2970 , n1144 , n1528 );
buf ( n2971 , n2970 );
xor ( n2972 , n1272 , n1400 );
buf ( n2973 , n2972 );
xor ( n2974 , n2971 , n2973 );
or ( n2975 , n2969 , n2974 );
xor ( n2976 , n1145 , n1529 );
buf ( n2977 , n2976 );
xor ( n2978 , n1273 , n1401 );
buf ( n2979 , n2978 );
xor ( n2980 , n2977 , n2979 );
or ( n2981 , n2975 , n2980 );
xor ( n2982 , n1146 , n1530 );
buf ( n2983 , n2982 );
xor ( n2984 , n1274 , n1402 );
buf ( n2985 , n2984 );
xor ( n2986 , n2983 , n2985 );
or ( n2987 , n2981 , n2986 );
xor ( n2988 , n1147 , n1531 );
buf ( n2989 , n2988 );
xor ( n2990 , n1275 , n1403 );
buf ( n2991 , n2990 );
xor ( n2992 , n2989 , n2991 );
or ( n2993 , n2987 , n2992 );
xor ( n2994 , n1148 , n1532 );
buf ( n2995 , n2994 );
xor ( n2996 , n1276 , n1404 );
buf ( n2997 , n2996 );
xor ( n2998 , n2995 , n2997 );
or ( n2999 , n2993 , n2998 );
xor ( n3000 , n1149 , n1533 );
buf ( n3001 , n3000 );
xor ( n3002 , n1277 , n1405 );
buf ( n3003 , n3002 );
xor ( n3004 , n3001 , n3003 );
or ( n3005 , n2999 , n3004 );
xor ( n3006 , n1150 , n1534 );
buf ( n3007 , n3006 );
xor ( n3008 , n1278 , n1406 );
buf ( n3009 , n3008 );
xor ( n3010 , n3007 , n3009 );
or ( n3011 , n3005 , n3010 );
xor ( n3012 , n1151 , n1535 );
buf ( n3013 , n3012 );
xor ( n3014 , n1279 , n1407 );
buf ( n3015 , n3014 );
xor ( n3016 , n3013 , n3015 );
or ( n3017 , n3011 , n3016 );
xor ( n3018 , n1152 , n1536 );
buf ( n3019 , n3018 );
xor ( n3020 , n1280 , n1408 );
buf ( n3021 , n3020 );
xor ( n3022 , n3019 , n3021 );
or ( n3023 , n3017 , n3022 );
xor ( n3024 , n1153 , n1537 );
buf ( n3025 , n3024 );
xor ( n3026 , n1281 , n1409 );
buf ( n3027 , n3026 );
xor ( n3028 , n3025 , n3027 );
or ( n3029 , n3023 , n3028 );
xor ( n3030 , n1154 , n1538 );
buf ( n3031 , n3030 );
xor ( n3032 , n1282 , n1410 );
buf ( n3033 , n3032 );
xor ( n3034 , n3031 , n3033 );
or ( n3035 , n3029 , n3034 );
xor ( n3036 , n1155 , n1539 );
buf ( n3037 , n3036 );
xor ( n3038 , n1283 , n1411 );
buf ( n3039 , n3038 );
xor ( n3040 , n3037 , n3039 );
or ( n3041 , n3035 , n3040 );
xor ( n3042 , n1156 , n1540 );
buf ( n3043 , n3042 );
xor ( n3044 , n1284 , n1412 );
buf ( n3045 , n3044 );
xor ( n3046 , n3043 , n3045 );
or ( n3047 , n3041 , n3046 );
xor ( n3048 , n1157 , n1541 );
buf ( n3049 , n3048 );
xor ( n3050 , n1285 , n1413 );
buf ( n3051 , n3050 );
xor ( n3052 , n3049 , n3051 );
or ( n3053 , n3047 , n3052 );
xor ( n3054 , n1158 , n1542 );
buf ( n3055 , n3054 );
xor ( n3056 , n1286 , n1414 );
buf ( n3057 , n3056 );
xor ( n3058 , n3055 , n3057 );
or ( n3059 , n3053 , n3058 );
xor ( n3060 , n1159 , n1543 );
buf ( n3061 , n3060 );
xor ( n3062 , n1287 , n1415 );
buf ( n3063 , n3062 );
xor ( n3064 , n3061 , n3063 );
or ( n3065 , n3059 , n3064 );
xor ( n3066 , n1160 , n1544 );
buf ( n3067 , n3066 );
xor ( n3068 , n1288 , n1416 );
buf ( n3069 , n3068 );
xor ( n3070 , n3067 , n3069 );
or ( n3071 , n3065 , n3070 );
xor ( n3072 , n1161 , n1545 );
buf ( n3073 , n3072 );
xor ( n3074 , n1289 , n1417 );
buf ( n3075 , n3074 );
xor ( n3076 , n3073 , n3075 );
or ( n3077 , n3071 , n3076 );
xor ( n3078 , n1162 , n1546 );
buf ( n3079 , n3078 );
xor ( n3080 , n1290 , n1418 );
buf ( n3081 , n3080 );
xor ( n3082 , n3079 , n3081 );
or ( n3083 , n3077 , n3082 );
xor ( n3084 , n1163 , n1547 );
buf ( n3085 , n3084 );
xor ( n3086 , n1291 , n1419 );
buf ( n3087 , n3086 );
xor ( n3088 , n3085 , n3087 );
or ( n3089 , n3083 , n3088 );
not ( n3090 , n3089 );
buf ( n3091 , n3090 );
or ( n3092 , n1160 , n1546 );
and ( n3093 , n3091 , n3092 );
buf ( n3094 , n3093 );
buf ( n3095 , n3094 );
buf ( n3096 , n2317 );
buf ( n3097 , n3096 );
buf ( n3098 , n2316 );
buf ( n3099 , n3091 );
endmodule
