module top( n2 , n11 , n13 , n16 , n21 , n44 , n45 , n46 , n55 ,
n74 , n75 , n81 , n84 , n85 , n87 , n93 , n96 , n98 , n101 ,
n105 , n111 , n123 , n128 , n131 , n134 , n139 , n148 , n153 , n159 ,
n163 , n177 , n191 , n196 , n199 , n206 , n211 , n216 , n223 , n226 ,
n240 , n243 , n254 , n260 , n264 , n266 , n280 , n282 , n283 , n287 ,
n290 , n291 , n299 , n309 , n336 , n346 , n349 , n360 , n368 , n369 ,
n377 , n388 , n394 , n409 , n428 , n435 , n442 , n447 , n449 , n454 ,
n457 , n468 , n471 , n481 , n484 , n494 , n500 , n507 , n511 , n518 ,
n519 , n525 , n534 , n542 , n547 , n557 , n561 , n568 , n569 , n571 ,
n575 , n581 , n582 , n583 , n587 , n600 , n603 , n609 , n613 , n614 ,
n616 , n627 , n635 , n646 , n659 , n661 , n664 , n672 , n673 );
    input n2 , n11 , n13 , n16 , n21 , n45 , n46 , n55 , n74 ,
n75 , n81 , n84 , n85 , n93 , n96 , n98 , n101 , n111 , n128 ,
n131 , n134 , n139 , n153 , n159 , n177 , n199 , n206 , n211 , n216 ,
n223 , n243 , n264 , n266 , n280 , n282 , n287 , n290 , n309 , n336 ,
n346 , n349 , n360 , n368 , n369 , n377 , n388 , n394 , n409 , n428 ,
n435 , n447 , n454 , n457 , n468 , n471 , n481 , n494 , n500 , n507 ,
n511 , n519 , n525 , n557 , n561 , n569 , n571 , n575 , n581 , n582 ,
n583 , n587 , n600 , n603 , n609 , n613 , n614 , n616 , n646 , n659 ,
n661 , n664 , n673 ;
    output n44 , n87 , n105 , n123 , n148 , n163 , n191 , n196 , n226 ,
n240 , n254 , n260 , n283 , n291 , n299 , n442 , n449 , n484 , n518 ,
n534 , n542 , n547 , n568 , n627 , n635 , n672 ;
    wire n0 , n1 , n3 , n4 , n5 , n6 , n7 , n8 , n9 ,
n10 , n12 , n14 , n15 , n17 , n18 , n19 , n20 , n22 , n23 ,
n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 ,
n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ,
n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n56 , n57 ,
n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 ,
n68 , n69 , n70 , n71 , n72 , n73 , n76 , n77 , n78 , n79 ,
n80 , n82 , n83 , n86 , n88 , n89 , n90 , n91 , n92 , n94 ,
n95 , n97 , n99 , n100 , n102 , n103 , n104 , n106 , n107 , n108 ,
n109 , n110 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 ,
n120 , n121 , n122 , n124 , n125 , n126 , n127 , n129 , n130 , n132 ,
n133 , n135 , n136 , n137 , n138 , n140 , n141 , n142 , n143 , n144 ,
n145 , n146 , n147 , n149 , n150 , n151 , n152 , n154 , n155 , n156 ,
n157 , n158 , n160 , n161 , n162 , n164 , n165 , n166 , n167 , n168 ,
n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n178 , n179 ,
n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 ,
n190 , n192 , n193 , n194 , n195 , n197 , n198 , n200 , n201 , n202 ,
n203 , n204 , n205 , n207 , n208 , n209 , n210 , n212 , n213 , n214 ,
n215 , n217 , n218 , n219 , n220 , n221 , n222 , n224 , n225 , n227 ,
n228 , n229 , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 ,
n238 , n239 , n241 , n242 , n244 , n245 , n246 , n247 , n248 , n249 ,
n250 , n251 , n252 , n253 , n255 , n256 , n257 , n258 , n259 , n261 ,
n262 , n263 , n265 , n267 , n268 , n269 , n270 , n271 , n272 , n273 ,
n274 , n275 , n276 , n277 , n278 , n279 , n281 , n284 , n285 , n286 ,
n288 , n289 , n292 , n293 , n294 , n295 , n296 , n297 , n298 , n300 ,
n301 , n302 , n303 , n304 , n305 , n306 , n307 , n308 , n310 , n311 ,
n312 , n313 , n314 , n315 , n316 , n317 , n318 , n319 , n320 , n321 ,
n322 , n323 , n324 , n325 , n326 , n327 , n328 , n329 , n330 , n331 ,
n332 , n333 , n334 , n335 , n337 , n338 , n339 , n340 , n341 , n342 ,
n343 , n344 , n345 , n347 , n348 , n350 , n351 , n352 , n353 , n354 ,
n355 , n356 , n357 , n358 , n359 , n361 , n362 , n363 , n364 , n365 ,
n366 , n367 , n370 , n371 , n372 , n373 , n374 , n375 , n376 , n378 ,
n379 , n380 , n381 , n382 , n383 , n384 , n385 , n386 , n387 , n389 ,
n390 , n391 , n392 , n393 , n395 , n396 , n397 , n398 , n399 , n400 ,
n401 , n402 , n403 , n404 , n405 , n406 , n407 , n408 , n410 , n411 ,
n412 , n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 ,
n422 , n423 , n424 , n425 , n426 , n427 , n429 , n430 , n431 , n432 ,
n433 , n434 , n436 , n437 , n438 , n439 , n440 , n441 , n443 , n444 ,
n445 , n446 , n448 , n450 , n451 , n452 , n453 , n455 , n456 , n458 ,
n459 , n460 , n461 , n462 , n463 , n464 , n465 , n466 , n467 , n469 ,
n470 , n472 , n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 ,
n482 , n483 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 ,
n493 , n495 , n496 , n497 , n498 , n499 , n501 , n502 , n503 , n504 ,
n505 , n506 , n508 , n509 , n510 , n512 , n513 , n514 , n515 , n516 ,
n517 , n520 , n521 , n522 , n523 , n524 , n526 , n527 , n528 , n529 ,
n530 , n531 , n532 , n533 , n535 , n536 , n537 , n538 , n539 , n540 ,
n541 , n543 , n544 , n545 , n546 , n548 , n549 , n550 , n551 , n552 ,
n553 , n554 , n555 , n556 , n558 , n559 , n560 , n562 , n563 , n564 ,
n565 , n566 , n567 , n570 , n572 , n573 , n574 , n576 , n577 , n578 ,
n579 , n580 , n584 , n585 , n586 , n588 , n589 , n590 , n591 , n592 ,
n593 , n594 , n595 , n596 , n597 , n598 , n599 , n601 , n602 , n604 ,
n605 , n606 , n607 , n608 , n610 , n611 , n612 , n615 , n617 , n618 ,
n619 , n620 , n621 , n622 , n623 , n624 , n625 , n626 , n628 , n629 ,
n630 , n631 , n632 , n633 , n634 , n636 , n637 , n638 , n639 , n640 ,
n641 , n642 , n643 , n644 , n645 , n647 , n648 , n649 , n650 , n651 ,
n652 , n653 , n654 , n655 , n656 , n657 , n658 , n660 , n662 , n663 ,
n665 , n666 , n667 , n668 , n669 , n670 , n671 ;
    and g0 ( n657 , n356 , n451 );
    and g1 ( n203 , n224 , n349 );
    and g2 ( n660 , n340 , n25 );
    nor g3 ( n347 , n468 , n417 );
    not g4 ( n253 , n54 );
    or g5 ( n6 , n48 , n383 );
    xnor g6 ( n291 , n339 , n668 );
    and g7 ( n308 , n515 , n168 );
    or g8 ( n629 , n253 , n652 );
    nor g9 ( n187 , n2 , n159 );
    not g10 ( n585 , n434 );
    buf g11 ( n570 , n389 );
    nor g12 ( n47 , n414 , n467 );
    xnor g13 ( n393 , n444 , n216 );
    not g14 ( n391 , n531 );
    not g15 ( n443 , n176 );
    xnor g16 ( n76 , n556 , n16 );
    xnor g17 ( n390 , n598 , n290 );
    not g18 ( n38 , n499 );
    or g19 ( n426 , n524 , n62 );
    nor g20 ( n117 , n93 , n396 );
    and g21 ( n89 , n9 , n72 );
    xnor g22 ( n628 , n107 , n531 );
    not g23 ( n550 , n159 );
    and g24 ( n365 , n321 , n253 );
    xnor g25 ( n163 , n0 , n479 );
    xnor g26 ( n61 , n7 , n613 );
    and g27 ( n648 , n127 , n125 );
    xnor g28 ( n283 , n31 , n648 );
    not g29 ( n608 , n31 );
    and g30 ( n327 , n638 , n367 );
    or g31 ( n444 , n285 , n412 );
    not g32 ( n373 , n639 );
    and g33 ( n602 , n570 , n101 );
    not g34 ( n251 , n75 );
    not g35 ( n107 , n520 );
    or g36 ( n427 , n608 , n125 );
    nor g37 ( n480 , n349 , n322 );
    and g38 ( n359 , n137 , n604 );
    nor g39 ( n95 , n13 , n2 );
    nor g40 ( n118 , n623 , n540 );
    not g41 ( n474 , n613 );
    nor g42 ( n115 , n93 , n37 );
    not g43 ( n398 , n0 );
    xnor g44 ( n289 , n280 , n287 );
    and g45 ( n543 , n390 , n266 );
    xnor g46 ( n60 , n624 , n464 );
    or g47 ( n141 , n538 , n452 );
    not g48 ( n572 , n466 );
    or g49 ( n339 , n5 , n492 );
    or g50 ( n31 , n559 , n424 );
    not g51 ( n514 , n206 );
    and g52 ( n234 , n198 , n326 );
    and g53 ( n258 , n19 , n266 );
    not g54 ( n300 , n428 );
    and g55 ( n651 , n526 , n570 );
    not g56 ( n197 , n138 );
    not g57 ( n351 , n508 );
    not g58 ( n649 , n225 );
    or g59 ( n100 , n413 , n179 );
    nor g60 ( n670 , n203 , n611 );
    or g61 ( n30 , n318 , n342 );
    or g62 ( n144 , n385 , n445 );
    or g63 ( n453 , n539 , n344 );
    not g64 ( n78 , n365 );
    and g65 ( n496 , n233 , n93 );
    nor g66 ( n179 , n570 , n330 );
    nor g67 ( n39 , n490 , n480 );
    not g68 ( n149 , n144 );
    nor g69 ( n182 , n183 , n370 );
    and g70 ( n9 , n513 , n551 );
    xnor g71 ( n152 , n356 , n616 );
    not g72 ( n576 , n100 );
    and g73 ( n662 , n580 , n264 );
    xnor g74 ( n123 , n182 , n463 );
    or g75 ( n65 , n201 , n439 );
    or g76 ( n259 , n58 , n1 );
    nor g77 ( n591 , n590 , n275 );
    and g78 ( n200 , n136 , n266 );
    not g79 ( n399 , n573 );
    or g80 ( n558 , n64 , n453 );
    or g81 ( n434 , n450 , n86 );
    or g82 ( n618 , n537 , n18 );
    and g83 ( n140 , n333 , n654 );
    xnor g84 ( n553 , n6 , n432 );
    or g85 ( n34 , n375 , n116 );
    and g86 ( n5 , n570 , n500 );
    nor g87 ( n530 , n472 , n327 );
    or g88 ( n626 , n384 , n642 );
    xnor g89 ( n401 , n582 , n2 );
    or g90 ( n450 , n190 , n307 );
    and g91 ( n106 , n465 , n608 );
    and g92 ( n40 , n421 , n93 );
    not g93 ( n520 , n248 );
    xnor g94 ( n299 , n395 , n175 );
    not g95 ( n501 , n171 );
    not g96 ( n420 , n45 );
    or g97 ( n169 , n319 , n629 );
    and g98 ( n637 , n124 , n335 );
    not g99 ( n621 , n380 );
    nor g100 ( n267 , n570 , n140 );
    xnor g101 ( n105 , n54 , n615 );
    or g102 ( n533 , n331 , n52 );
    or g103 ( n355 , n71 , n591 );
    xnor g104 ( n260 , n508 , n669 );
    or g105 ( n594 , n514 , n516 );
    nor g106 ( n395 , n431 , n663 );
    xnor g107 ( n302 , n453 , n336 );
    or g108 ( n363 , n526 , n239 );
    and g109 ( n238 , n42 , n93 );
    and g110 ( n424 , n61 , n266 );
    and g111 ( n567 , n77 , n569 );
    and g112 ( n79 , n29 , n266 );
    or g113 ( n598 , n298 , n460 );
    xnor g114 ( n620 , n632 , n392 );
    nor g115 ( n479 , n185 , n425 );
    not g116 ( n143 , n339 );
    buf g117 ( n77 , n389 );
    or g118 ( n624 , n285 , n305 );
    and g119 ( n218 , n249 , n266 );
    and g120 ( n3 , n147 , n266 );
    nor g121 ( n88 , n199 , n85 );
    xnor g122 ( n249 , n426 , n282 );
    or g123 ( n380 , n358 , n597 );
    or g124 ( n654 , n58 , n562 );
    or g125 ( n165 , n201 , n660 );
    nor g126 ( n212 , n75 , n131 );
    not g127 ( n623 , n577 );
    or g128 ( n7 , n636 , n477 );
    nor g129 ( n340 , n170 , n418 );
    or g130 ( n114 , n482 , n444 );
    not g131 ( n560 , n209 );
    and g132 ( n580 , n666 , n43 );
    and g133 ( n274 , n570 , n603 );
    not g134 ( n1 , n381 );
    xnor g135 ( n484 , n180 , n584 );
    or g136 ( n592 , n606 , n503 );
    and g137 ( n222 , n26 , n436 );
    or g138 ( n335 , n397 , n517 );
    not g139 ( n461 , n13 );
    nor g140 ( n650 , n665 , n15 );
    or g141 ( n552 , n220 , n461 );
    or g142 ( n475 , n227 , n637 );
    or g143 ( n386 , n231 , n323 );
    or g144 ( n130 , n440 , n548 );
    nor g145 ( n312 , n77 , n637 );
    or g146 ( n463 , n566 , n543 );
    or g147 ( n497 , n538 , n278 );
    or g148 ( n655 , n470 , n324 );
    or g149 ( n257 , n387 , n200 );
    and g150 ( n110 , n65 , n601 );
    and g151 ( n478 , n570 , n153 );
    or g152 ( n90 , n653 , n459 );
    and g153 ( n658 , n302 , n266 );
    xnor g154 ( n262 , n177 , n75 );
    not g155 ( n155 , n521 );
    not g156 ( n383 , n468 );
    or g157 ( n167 , n359 , n219 );
    not g158 ( n15 , n373 );
    or g159 ( n247 , n662 , n404 );
    and g160 ( n640 , n284 , n552 );
    not g161 ( n201 , n352 );
    nor g162 ( n415 , n194 , n133 );
    or g163 ( n367 , n625 , n209 );
    xnor g164 ( n635 , n12 , n4 );
    not g165 ( n207 , n641 );
    or g166 ( n344 , n429 , n353 );
    nor g167 ( n192 , n34 , n517 );
    and g168 ( n189 , n235 , n487 );
    or g169 ( n261 , n428 , n48 );
    not g170 ( n389 , n266 );
    xnor g171 ( n148 , n36 , n17 );
    and g172 ( n372 , n57 , n266 );
    or g173 ( n579 , n586 , n78 );
    and g174 ( n374 , n393 , n206 );
    or g175 ( n124 , n334 , n140 );
    not g176 ( n174 , n51 );
    and g177 ( n4 , n434 , n52 );
    not g178 ( n588 , n388 );
    and g179 ( n269 , n564 , n126 );
    or g180 ( n156 , n63 , n495 );
    and g181 ( n286 , n455 , n482 );
    nor g182 ( n161 , n657 , n438 );
    not g183 ( n483 , n6 );
    not g184 ( n509 , n368 );
    nor g185 ( n541 , n472 , n39 );
    not g186 ( n43 , n93 );
    not g187 ( n64 , n336 );
    or g188 ( n284 , n95 , n294 );
    not g189 ( n328 , n631 );
    xnor g190 ( n464 , n511 , n454 );
    and g191 ( n433 , n158 , n441 );
    not g192 ( n563 , n511 );
    and g193 ( n71 , n2 , n582 );
    and g194 ( n67 , n94 , n35 );
    or g195 ( n456 , n251 , n8 );
    nor g196 ( n217 , n135 , n419 );
    not g197 ( n448 , n595 );
    not g198 ( n310 , n533 );
    nor g199 ( n265 , n289 , n316 );
    or g200 ( n151 , n286 , n408 );
    or g201 ( n281 , n221 , n593 );
    xnor g202 ( n568 , n217 , n406 );
    and g203 ( n644 , n570 , n614 );
    not g204 ( n73 , n450 );
    xnor g205 ( n154 , n459 , n583 );
    and g206 ( n532 , n475 , n167 );
    xnor g207 ( n607 , n355 , n97 );
    and g208 ( n256 , n553 , n93 );
    and g209 ( n150 , n570 , n519 );
    nor g210 ( n304 , n107 , n219 );
    not g211 ( n80 , n352 );
    and g212 ( n667 , n639 , n174 );
    not g213 ( n248 , n359 );
    xnor g214 ( n87 , n156 , n49 );
    or g215 ( n168 , n359 , n271 );
    or g216 ( n403 , n451 , n295 );
    not g217 ( n324 , n560 );
    and g218 ( n593 , n546 , n527 );
    not g219 ( n215 , n235 );
    and g220 ( n32 , n659 , n93 );
    xnor g221 ( n458 , n294 , n112 );
    or g222 ( n513 , n187 , n632 );
    or g223 ( n467 , n206 , n509 );
    or g224 ( n385 , n237 , n129 );
    or g225 ( n72 , n251 , n121 );
    not g226 ( n517 , n197 );
    not g227 ( n8 , n177 );
    not g228 ( n482 , n216 );
    nor g229 ( n337 , n443 , n269 );
    or g230 ( n476 , n650 , n50 );
    nor g231 ( n638 , n229 , n265 );
    not g232 ( n319 , n586 );
    or g233 ( n157 , n212 , n89 );
    xnor g234 ( n240 , n341 , n402 );
    not g235 ( n24 , n491 );
    or g236 ( n295 , n493 , n114 );
    xnor g237 ( n627 , n130 , n366 );
    not g238 ( n625 , n664 );
    or g239 ( n178 , n616 , n66 );
    or g240 ( n642 , n505 , n90 );
    or g241 ( n311 , n228 , n363 );
    nor g242 ( n33 , n620 , n623 );
    nor g243 ( n18 , n77 , n60 );
    or g244 ( n171 , n351 , n169 );
    or g245 ( n341 , n343 , n345 );
    and g246 ( n68 , n570 , n581 );
    or g247 ( n556 , n102 , n329 );
    nor g248 ( n437 , n119 , n293 );
    not g249 ( n606 , n646 );
    not g250 ( n565 , n624 );
    not g251 ( n412 , n454 );
    not g252 ( n473 , n432 );
    not g253 ( n462 , n381 );
    or g254 ( n503 , n315 , n426 );
    not g255 ( n48 , n409 );
    not g256 ( n285 , n659 );
    nor g257 ( n27 , n119 , n356 );
    xnor g258 ( n263 , n626 , n388 );
    not g259 ( n430 , n579 );
    xnor g260 ( n112 , n13 , n2 );
    not g261 ( n536 , n561 );
    or g262 ( n527 , n478 , n574 );
    nor g263 ( n358 , n20 , n43 );
    or g264 ( n632 , n276 , n120 );
    not g265 ( n505 , n55 );
    and g266 ( n313 , n386 , n259 );
    or g267 ( n104 , n511 , n659 );
    nor g268 ( n296 , n435 , n75 );
    and g269 ( n146 , n454 , n511 );
    and g270 ( n307 , n272 , n266 );
    not g271 ( n321 , n656 );
    not g272 ( n554 , n555 );
    not g273 ( n276 , n287 );
    xnor g274 ( n442 , n172 , n382 );
    nor g275 ( n619 , n6 , n473 );
    and g276 ( n396 , n165 , n522 );
    and g277 ( n566 , n77 , n74 );
    not g278 ( n22 , n425 );
    not g279 ( n120 , n96 );
    nor g280 ( n323 , n306 , n562 );
    xor g281 ( n224 , n275 , n401 );
    not g282 ( n315 , n282 );
    and g283 ( n23 , n596 , n155 );
    or g284 ( n172 , n274 , n325 );
    not g285 ( n306 , n576 );
    or g286 ( n241 , n506 , n592 );
    or g287 ( n528 , n405 , n427 );
    and g288 ( n63 , n570 , n139 );
    and g289 ( n183 , n242 , n555 );
    nor g290 ( n378 , n292 , n193 );
    xnor g291 ( n20 , n428 , n454 );
    nor g292 ( n666 , n80 , n209 );
    and g293 ( n669 , n579 , n169 );
    or g294 ( n353 , n634 , n612 );
    not g295 ( n126 , n350 );
    and g296 ( n548 , n622 , n266 );
    xnor g297 ( n42 , n10 , n202 );
    or g298 ( n508 , n166 , n258 );
    and g299 ( n488 , n279 , n77 );
    xnor g300 ( n498 , n423 , n45 );
    nor g301 ( n116 , n77 , n76 );
    or g302 ( n489 , n437 , n10 );
    and g303 ( n37 , n273 , n594 );
    not g304 ( n510 , n211 );
    not g305 ( n278 , n38 );
    or g306 ( n460 , n230 , n558 );
    xnor g307 ( n226 , n213 , n245 );
    not g308 ( n397 , n448 );
    and g309 ( n559 , n77 , n609 );
    and g310 ( n371 , n77 , n11 );
    not g311 ( n405 , n172 );
    or g312 ( n555 , n486 , n647 );
    not g313 ( n268 , n629 );
    and g314 ( n589 , n106 , n405 );
    or g315 ( n205 , n422 , n241 );
    not g316 ( n665 , n51 );
    xnor g317 ( n421 , n455 , n103 );
    and g318 ( n186 , n580 , n21 );
    and g319 ( n417 , n409 , n428 );
    or g320 ( n209 , n85 , n349 );
    xnor g321 ( n293 , n261 , n468 );
    xnor g322 ( n516 , n214 , n114 );
    and g323 ( n135 , n231 , n77 );
    xnor g324 ( n518 , n555 , n195 );
    and g325 ( n633 , n624 , n104 );
    and g326 ( n438 , n489 , n178 );
    nor g327 ( n663 , n570 , n532 );
    or g328 ( n12 , n602 , n3 );
    nor g329 ( n82 , n160 , n312 );
    nor g330 ( n504 , n296 , n91 );
    nor g331 ( n250 , n177 , n75 );
    not g332 ( n384 , n128 );
    and g333 ( n142 , n236 , n497 );
    not g334 ( n599 , n216 );
    or g335 ( n645 , n59 , n228 );
    or g336 ( n436 , n485 , n23 );
    not g337 ( n564 , n132 );
    nor g338 ( n162 , n514 , n643 );
    and g339 ( n108 , n210 , n85 );
    and g340 ( n173 , n317 , n266 );
    or g341 ( n596 , n32 , n332 );
    nor g342 ( n50 , n667 , n532 );
    not g343 ( n230 , n494 );
    not g344 ( n305 , n511 );
    not g345 ( n298 , n223 );
    or g346 ( n350 , n68 , n529 );
    and g347 ( n160 , n67 , n77 );
    or g348 ( n326 , n599 , n305 );
    and g349 ( n366 , n144 , n184 );
    not g350 ( n485 , n618 );
    not g351 ( n577 , n467 );
    not g352 ( n109 , n527 );
    nor g353 ( n522 , n374 , n118 );
    and g354 ( n615 , n656 , n652 );
    and g355 ( n537 , n77 , n46 );
    and g356 ( n431 , n308 , n570 );
    or g357 ( n254 , n411 , n281 );
    nor g358 ( n597 , n93 , n110 );
    xnor g359 ( n147 , n344 , n369 );
    or g360 ( n499 , n40 , n117 );
    not g361 ( n121 , n131 );
    nor g362 ( n601 , n33 , n162 );
    not g363 ( n127 , n465 );
    or g364 ( n26 , n380 , n354 );
    xnor g365 ( n17 , n448 , n138 );
    and g366 ( n231 , n181 , n141 );
    not g367 ( n198 , n288 );
    and g368 ( n387 , n570 , n457 );
    not g369 ( n653 , n583 );
    nor g370 ( n590 , n582 , n2 );
    and g371 ( n361 , n28 , n53 );
    xnor g372 ( n136 , n288 , n113 );
    or g373 ( n652 , n266 , n415 );
    or g374 ( n531 , n186 , n256 );
    and g375 ( n166 , n570 , n571 );
    not g376 ( n610 , n138 );
    and g377 ( n297 , n498 , n266 );
    or g378 ( n94 , n192 , n313 );
    not g379 ( n145 , n130 );
    or g380 ( n193 , n47 , n530 );
    not g381 ( n232 , n377 );
    or g382 ( n342 , n145 , n184 );
    or g383 ( n138 , n247 , n496 );
    not g384 ( n470 , n525 );
    nor g385 ( n213 , n488 , n362 );
    and g386 ( n325 , n154 , n266 );
    and g387 ( n382 , n446 , n427 );
    not g388 ( n429 , n575 );
    not g389 ( n538 , n207 );
    xnor g390 ( n449 , n155 , n596 );
    and g391 ( n418 , n607 , n349 );
    or g392 ( n176 , n126 , n30 );
    and g393 ( n605 , n570 , n84 );
    or g394 ( n70 , n143 , n171 );
    and g395 ( n370 , n411 , n554 );
    not g396 ( n86 , n269 );
    not g397 ( n119 , n616 );
    nor g398 ( n273 , n502 , n541 );
    not g399 ( n441 , n239 );
    or g400 ( n316 , n349 , n92 );
    and g401 ( n630 , n149 , n145 );
    or g402 ( n294 , n276 , n545 );
    not g403 ( n318 , n341 );
    not g404 ( n219 , n391 );
    or g405 ( n604 , n266 , n232 );
    nor g406 ( n402 , n416 , n630 );
    xnor g407 ( n672 , n385 , n400 );
    not g408 ( n208 , n528 );
    xnor g409 ( n272 , n353 , n575 );
    not g410 ( n320 , n600 );
    xnor g411 ( n376 , n511 , n616 );
    or g412 ( n52 , n73 , n176 );
    not g413 ( n314 , n109 );
    not g414 ( n92 , n85 );
    nor g415 ( n611 , n458 , n316 );
    or g416 ( n181 , n122 , n279 );
    not g417 ( n53 , n180 );
    and g418 ( n338 , n75 , n435 );
    xnor g419 ( n245 , n207 , n499 );
    xnor g420 ( n244 , n558 , n494 );
    not g421 ( n521 , n526 );
    not g422 ( n14 , n23 );
    xnor g423 ( n540 , n9 , n164 );
    and g424 ( n574 , n244 , n266 );
    and g425 ( n303 , n77 , n346 );
    or g426 ( n132 , n341 , n56 );
    not g427 ( n422 , n557 );
    and g428 ( n529 , n469 , n266 );
    and g429 ( n671 , n313 , n77 );
    nor g430 ( n419 , n77 , n142 );
    nor g431 ( n354 , n618 , n14 );
    or g432 ( n255 , n563 , n348 );
    nor g433 ( n221 , n527 , n225 );
    or g434 ( n54 , n605 , n79 );
    nor g435 ( n102 , n563 , n214 );
    or g436 ( n25 , n510 , n324 );
    nor g437 ( n204 , n257 , n452 );
    nor g438 ( n362 , n570 , n222 );
    not g439 ( n636 , n471 );
    or g440 ( n252 , n599 , n455 );
    or g441 ( n356 , n483 , n347 );
    not g442 ( n524 , n111 );
    and g443 ( n413 , n77 , n507 );
    nor g444 ( n292 , n659 , n493 );
    xnor g445 ( n357 , n241 , n557 );
    nor g446 ( n133 , n99 , n308 );
    and g447 ( n647 , n410 , n266 );
    or g448 ( n639 , n277 , n549 );
    and g449 ( n495 , n357 , n266 );
    nor g450 ( n36 , n671 , n267 );
    not g451 ( n329 , n234 );
    or g452 ( n35 , n397 , n610 );
    and g453 ( n526 , n24 , n270 );
    or g454 ( n0 , n303 , n173 );
    not g455 ( n379 , n156 );
    or g456 ( n586 , n371 , n218 );
    and g457 ( n28 , n585 , n331 );
    xnor g458 ( n57 , n477 , n471 );
    or g459 ( n472 , n368 , n206 );
    or g460 ( n180 , n567 , n658 );
    xnor g461 ( n535 , n90 , n55 );
    or g462 ( n656 , n77 , n476 );
    nor g463 ( n91 , n338 , n355 );
    xnor g464 ( n44 , n466 , n189 );
    not g465 ( n41 , n16 );
    or g466 ( n381 , n238 , n115 );
    not g467 ( n56 , n630 );
    not g468 ( n451 , n616 );
    and g469 ( n99 , n373 , n174 );
    not g470 ( n348 , n423 );
    or g471 ( n322 , n88 , n108 );
    xnor g472 ( n233 , n438 , n152 );
    not g473 ( n220 , n2 );
    not g474 ( n506 , n243 );
    or g475 ( n235 , n0 , n22 );
    or g476 ( n184 , n69 , n528 );
    not g477 ( n539 , n369 );
    or g478 ( n270 , n266 , n83 );
    or g479 ( n551 , n220 , n550 );
    nor g480 ( n188 , n268 , n365 );
    and g481 ( n465 , n215 , n572 );
    xnor g482 ( n410 , n460 , n223 );
    nor g483 ( n195 , n242 , n411 );
    nor g484 ( n122 , n257 , n278 );
    or g485 ( n288 , n146 , n565 );
    xnor g486 ( n408 , n428 , n409 );
    and g487 ( n49 , n573 , n70 );
    and g488 ( n578 , n640 , n456 );
    xnor g489 ( n547 , n82 , n628 );
    not g490 ( n493 , n206 );
    not g491 ( n331 , n12 );
    nor g492 ( n400 , n208 , n589 );
    not g493 ( n66 , n293 );
    or g494 ( n51 , n150 , n297 );
    and g495 ( n631 , n430 , n351 );
    not g496 ( n214 , n616 );
    or g497 ( n236 , n204 , n222 );
    and g498 ( n343 , n77 , n360 );
    nor g499 ( n668 , n501 , n631 );
    or g500 ( n137 , n77 , n255 );
    xnor g501 ( n406 , n306 , n381 );
    not g502 ( n185 , n544 );
    not g503 ( n641 , n257 );
    or g504 ( n62 , n420 , n423 );
    xnor g505 ( n246 , n640 , n262 );
    and g506 ( n229 , n364 , n349 );
    or g507 ( n59 , n491 , n651 );
    not g508 ( n271 , n531 );
    nor g509 ( n227 , n248 , n271 );
    or g510 ( n158 , n407 , n621 );
    and g511 ( n242 , n649 , n314 );
    and g512 ( n277 , n580 , n98 );
    xnor g513 ( n29 , n62 , n111 );
    and g514 ( n190 , n570 , n134 );
    and g515 ( n491 , n633 , n266 );
    and g516 ( n549 , n619 , n93 );
    not g517 ( n634 , n661 );
    or g518 ( n333 , n617 , n142 );
    xnor g519 ( n202 , n293 , n616 );
    xnor g520 ( n196 , n645 , n433 );
    not g521 ( n58 , n100 );
    or g522 ( n459 , n474 , n7 );
    xor g523 ( n364 , n600 , n287 );
    xnor g524 ( n622 , n642 , n128 );
    xnor g525 ( n643 , n659 , n454 );
    and g526 ( n486 , n77 , n309 );
    or g527 ( n515 , n304 , n67 );
    xnor g528 ( n414 , n287 , n96 );
    and g529 ( n194 , n15 , n51 );
    and g530 ( n490 , n504 , n349 );
    nor g531 ( n584 , n310 , n28 );
    not g532 ( n446 , n106 );
    xnor g533 ( n191 , n350 , n523 );
    or g534 ( n125 , n572 , n487 );
    xnor g535 ( n103 , n408 , n216 );
    xnor g536 ( n469 , n612 , n661 );
    not g537 ( n228 , n596 );
    nor g538 ( n332 , n93 , n378 );
    nor g539 ( n502 , n467 , n157 );
    and g540 ( n10 , n151 , n252 );
    not g541 ( n512 , n556 );
    and g542 ( n237 , n570 , n447 );
    or g543 ( n573 , n339 , n328 );
    xnor g544 ( n164 , n75 , n131 );
    not g545 ( n69 , n385 );
    or g546 ( n225 , n53 , n533 );
    and g547 ( n239 , n621 , n407 );
    or g548 ( n466 , n644 , n372 );
    not g549 ( n407 , n618 );
    and g550 ( n523 , n132 , n30 );
    or g551 ( n175 , n99 , n194 );
    and g552 ( n440 , n570 , n394 );
    or g553 ( n544 , n379 , n70 );
    or g554 ( n487 , n398 , n544 );
    not g555 ( n545 , n280 );
    xnor g556 ( n534 , n586 , n188 );
    or g557 ( n210 , n250 , n578 );
    xnor g558 ( n542 , n450 , n337 );
    and g559 ( n279 , n311 , n158 );
    or g560 ( n275 , n276 , n320 );
    xnor g561 ( n330 , n234 , n376 );
    not g562 ( n416 , n342 );
    nor g563 ( n546 , n649 , n361 );
    or g564 ( n477 , n536 , n205 );
    and g565 ( n411 , n361 , n109 );
    not g566 ( n352 , n472 );
    or g567 ( n612 , n588 , n626 );
    not g568 ( n452 , n499 );
    or g569 ( n423 , n41 , n512 );
    and g570 ( n375 , n77 , n81 );
    and g571 ( n492 , n301 , n266 );
    xnor g572 ( n392 , n2 , n159 );
    and g573 ( n129 , n535 , n266 );
    not g574 ( n562 , n462 );
    nor g575 ( n334 , n34 , n610 );
    xnor g576 ( n113 , n511 , n216 );
    and g577 ( n439 , n670 , n655 );
    or g578 ( n455 , n300 , n412 );
    and g579 ( n345 , n263 , n266 );
    nor g580 ( n617 , n100 , n1 );
    xnor g581 ( n97 , n435 , n75 );
    and g582 ( n425 , n399 , n379 );
    or g583 ( n432 , n27 , n161 );
    xnor g584 ( n301 , n592 , n243 );
    not g585 ( n445 , n589 );
    xnor g586 ( n317 , n205 , n561 );
    xnor g587 ( n19 , n503 , n646 );
    not g588 ( n595 , n34 );
    nor g589 ( n404 , n93 , n403 );
    nor g590 ( n170 , n316 , n246 );
    not g591 ( n83 , n673 );
endmodule