//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 ;
output n36 , n37 , n38 , n39 , n40 , n41 , n42 ;

wire n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 ,
     n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 ,
     n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ,
     n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 ,
     n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 ,
     n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 ,
     n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 ,
     n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 ,
     n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 ,
     n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 ,
     n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 ,
     n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 ,
     n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 ,
     n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 ,
     n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , n234 ,
     n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 ,
     n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 ,
     n255 , n256 , n257 , n258 , n259 , n260 , n261 , n262 , n263 , n264 ,
     n265 , n266 , n267 , n268 , n269 , n270 , n271 , n272 , n273 , n274 ,
     n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 , n283 , n284 ,
     n285 , n286 , n287 , n288 , n289 , n290 , n291 , n292 , n293 , n294 ,
     n295 , n296 , n297 ;
buf ( n36 , n145 );
buf ( n41 , n186 );
buf ( n39 , n236 );
buf ( n42 , n280 );
buf ( n37 , n285 );
buf ( n38 , n292 );
buf ( n40 , n297 );
buf ( n88 , n35 );
buf ( n89 , n3 );
buf ( n90 , n13 );
buf ( n91 , n25 );
buf ( n92 , n21 );
buf ( n93 , n4 );
buf ( n94 , n33 );
buf ( n95 , n6 );
buf ( n96 , n11 );
buf ( n97 , n15 );
buf ( n98 , n24 );
buf ( n99 , n29 );
buf ( n100 , n19 );
buf ( n101 , n18 );
buf ( n102 , n10 );
buf ( n103 , n0 );
buf ( n104 , n9 );
buf ( n105 , n31 );
buf ( n106 , n5 );
buf ( n107 , n14 );
buf ( n108 , n16 );
buf ( n109 , n12 );
buf ( n110 , n23 );
buf ( n111 , n34 );
buf ( n112 , n28 );
buf ( n113 , n1 );
buf ( n114 , n22 );
buf ( n115 , n8 );
buf ( n116 , n7 );
buf ( n117 , n30 );
buf ( n118 , n27 );
buf ( n119 , n26 );
buf ( n120 , n20 );
buf ( n121 , n17 );
buf ( n122 , n32 );
buf ( n123 , n2 );
not ( n124 , n88 );
nand ( n125 , n124 , n89 );
not ( n126 , n91 );
nand ( n127 , n126 , n93 );
not ( n128 , n95 );
nand ( n129 , n128 , n97 );
not ( n130 , n99 );
nand ( n131 , n130 , n101 );
not ( n132 , n103 );
nand ( n133 , n132 , n105 );
not ( n134 , n107 );
nand ( n135 , n134 , n109 );
not ( n136 , n111 );
nand ( n137 , n136 , n113 );
not ( n138 , n115 );
nand ( n139 , n138 , n117 );
not ( n140 , n119 );
nand ( n141 , n140 , n121 );
and ( n142 , n125 , n127 , n129 , n131 , n133 , n135 , n137 , n139 , n141 );
not ( n143 , n142 );
buf ( n144 , n143 );
buf ( n145 , n144 );
not ( n146 , n142 );
xor ( n147 , n146 , n125 );
not ( n148 , n89 );
nor ( n149 , n90 , n148 );
nand ( n150 , n147 , n149 );
xor ( n151 , n146 , n127 );
not ( n152 , n93 );
nor ( n153 , n94 , n152 );
nand ( n154 , n151 , n153 );
xor ( n155 , n146 , n129 );
not ( n156 , n97 );
nor ( n157 , n98 , n156 );
nand ( n158 , n155 , n157 );
xor ( n159 , n146 , n131 );
not ( n160 , n101 );
nor ( n161 , n102 , n160 );
nand ( n162 , n159 , n161 );
xor ( n163 , n146 , n133 );
not ( n164 , n105 );
nor ( n165 , n106 , n164 );
nand ( n166 , n163 , n165 );
xor ( n167 , n146 , n135 );
not ( n168 , n109 );
nor ( n169 , n110 , n168 );
nand ( n170 , n167 , n169 );
xor ( n171 , n146 , n137 );
not ( n172 , n113 );
nor ( n173 , n114 , n172 );
nand ( n174 , n171 , n173 );
xor ( n175 , n146 , n139 );
not ( n176 , n117 );
nor ( n177 , n118 , n176 );
nand ( n178 , n175 , n177 );
xor ( n179 , n146 , n141 );
not ( n180 , n121 );
nor ( n181 , n122 , n180 );
nand ( n182 , n179 , n181 );
and ( n183 , n150 , n154 , n158 , n162 , n166 , n170 , n174 , n178 , n182 );
not ( n184 , n183 );
buf ( n185 , n184 );
buf ( n186 , n185 );
not ( n187 , n183 );
xor ( n188 , n187 , n150 );
nor ( n189 , n92 , n148 );
nand ( n190 , n147 , n189 );
not ( n191 , n190 );
nand ( n192 , n188 , n191 );
xor ( n193 , n187 , n154 );
nor ( n194 , n96 , n152 );
nand ( n195 , n151 , n194 );
not ( n196 , n195 );
nand ( n197 , n193 , n196 );
xor ( n198 , n187 , n158 );
nor ( n199 , n100 , n156 );
nand ( n200 , n155 , n199 );
not ( n201 , n200 );
nand ( n202 , n198 , n201 );
xor ( n203 , n187 , n162 );
nor ( n204 , n104 , n160 );
nand ( n205 , n159 , n204 );
not ( n206 , n205 );
nand ( n207 , n203 , n206 );
xor ( n208 , n187 , n166 );
nor ( n209 , n108 , n164 );
nand ( n210 , n163 , n209 );
not ( n211 , n210 );
nand ( n212 , n208 , n211 );
xor ( n213 , n187 , n170 );
nor ( n214 , n112 , n168 );
nand ( n215 , n167 , n214 );
not ( n216 , n215 );
nand ( n217 , n213 , n216 );
xor ( n218 , n187 , n174 );
nor ( n219 , n116 , n172 );
nand ( n220 , n171 , n219 );
not ( n221 , n220 );
nand ( n222 , n218 , n221 );
xor ( n223 , n187 , n178 );
nor ( n224 , n120 , n176 );
nand ( n225 , n175 , n224 );
not ( n226 , n225 );
nand ( n227 , n223 , n226 );
xor ( n228 , n187 , n182 );
nor ( n229 , n123 , n180 );
nand ( n230 , n179 , n229 );
not ( n231 , n230 );
nand ( n232 , n228 , n231 );
and ( n233 , n192 , n197 , n202 , n207 , n212 , n217 , n222 , n227 , n232 );
not ( n234 , n233 );
buf ( n235 , n234 );
buf ( n236 , n235 );
not ( n237 , n142 );
nand ( n238 , n88 , n237 );
not ( n239 , n183 );
nand ( n240 , n90 , n239 );
not ( n241 , n233 );
nand ( n242 , n92 , n241 );
nand ( n243 , n89 , n238 , n240 , n242 );
not ( n244 , n243 );
nand ( n245 , n237 , n91 );
nand ( n246 , n239 , n94 );
nand ( n247 , n241 , n96 );
nand ( n248 , n245 , n246 , n247 , n93 );
nand ( n249 , n237 , n95 );
nand ( n250 , n239 , n98 );
nand ( n251 , n241 , n100 );
nand ( n252 , n249 , n250 , n251 , n97 );
nand ( n253 , n237 , n99 );
nand ( n254 , n239 , n102 );
nand ( n255 , n241 , n104 );
nand ( n256 , n253 , n254 , n255 , n101 );
nand ( n257 , n237 , n103 );
nand ( n258 , n239 , n106 );
nand ( n259 , n241 , n108 );
nand ( n260 , n257 , n258 , n259 , n105 );
nand ( n261 , n237 , n107 );
nand ( n262 , n239 , n110 );
nand ( n263 , n241 , n112 );
nand ( n264 , n261 , n262 , n263 , n109 );
nand ( n265 , n237 , n111 );
nand ( n266 , n239 , n114 );
nand ( n267 , n241 , n116 );
nand ( n268 , n265 , n266 , n267 , n113 );
nand ( n269 , n237 , n115 );
nand ( n270 , n239 , n118 );
nand ( n271 , n241 , n120 );
nand ( n272 , n269 , n270 , n271 , n117 );
nand ( n273 , n237 , n119 );
nand ( n274 , n239 , n122 );
nand ( n275 , n241 , n123 );
nand ( n276 , n273 , n274 , n275 , n121 );
and ( n277 , n248 , n252 , n256 , n260 , n264 , n268 , n272 , n276 );
nor ( n278 , n244 , n277 );
buf ( n279 , n278 );
buf ( n280 , n279 );
not ( n281 , n256 );
nand ( n282 , n252 , n281 );
nand ( n283 , n248 , n252 , n282 , n260 );
buf ( n284 , n283 );
buf ( n285 , n284 );
not ( n286 , n264 );
nand ( n287 , n252 , n256 , n286 , n260 );
not ( n288 , n268 );
nand ( n289 , n260 , n256 , n288 );
nand ( n290 , n248 , n252 , n287 , n289 );
buf ( n291 , n290 );
buf ( n292 , n291 );
not ( n293 , n272 );
nand ( n294 , n252 , n256 , n268 , n293 );
nand ( n295 , n248 , n282 , n287 , n294 );
buf ( n296 , n295 );
buf ( n297 , n296 );
endmodule
