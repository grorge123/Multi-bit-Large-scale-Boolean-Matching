//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n9999, n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , PI_PI_clock , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , PI_DFF_state_reg_Q , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , PI_PI_reset , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , PI_DFF_B_reg_Q , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , PI_DFF_rd_reg_Q , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , PI_DFF_wr_reg_Q , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 );
input n9999, n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , PI_PI_clock , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , PI_DFF_state_reg_Q , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , PI_PI_reset , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , PI_DFF_B_reg_Q , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , PI_DFF_rd_reg_Q , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , PI_DFF_wr_reg_Q , n230 , n231 , n232 , n233 , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 ;
output n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 ;

wire n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 ,
     n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 ,
     n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 ,
     n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 ,
     n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 ,
     n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 ,
     n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 ,
     n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 ,
     n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 ,
     n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 ,
     n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 ,
     n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 ,
     n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 ,
     n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 ,
     n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 ,
     n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 ,
     n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 ,
     n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 ,
     n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 ,
     n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 ,
     n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 ,
     n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 ,
     n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 ,
     n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 ,
     n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 ,
     n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 ,
     n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 ,
     n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 ,
     n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 ,
     n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 ,
     n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 ,
     n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 ,
     n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 ,
     n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 ,
     n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 ,
     n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 ,
     n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 ,
     n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 ,
     n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 ,
     n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 ,
     n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 ,
     n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 ,
     n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 ,
     n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 ,
     n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 ,
     n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 ,
     n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 ,
     n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 ,
     n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 ,
     n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 ,
     n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 ,
     n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 ,
     n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 ,
     n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 ,
     n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 ,
     n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 ,
     n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 ,
     n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 ,
     n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 ,
     n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 ,
     n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 ,
     n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 ,
     n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 ,
     n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 ,
     n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 ,
     n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 ,
     n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 ,
     n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 ,
     n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 ,
     n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 ,
     n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 ,
     n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 ,
     n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 ,
     n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 ,
     n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 ,
     n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 ,
     n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 ,
     n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 ,
     n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 ,
     n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 ,
     n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 ,
     n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 ,
     n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 ,
     n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 ,
     n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 ,
     n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 ,
     n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 ,
     n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 ,
     n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 ,
     n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 ,
     n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 ,
     n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 ,
     n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 ,
     n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 ,
     n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 ,
     n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 ,
     n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 ,
     n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 ,
     n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 ,
     n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 ,
     n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 ,
     n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 ,
     n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 ,
     n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 ,
     n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 ,
     n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 ,
     n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 ,
     n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 ,
     n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 ,
     n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 ,
     n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 ,
     n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 ,
     n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 ,
     n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 ,
     n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 ,
     n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 ,
     n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 ,
     n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 ,
     n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 ,
     n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 ,
     n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 ,
     n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 ,
     n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 ,
     n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 ,
     n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 ,
     n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 ,
     n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 ,
     n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 ,
     n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 ,
     n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 ,
     n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 ,
     n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 ,
     n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 ,
     n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 ,
     n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 ,
     n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 ,
     n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 ,
     n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 ,
     n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 ,
     n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 ,
     n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 ,
     n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 ,
     n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 ,
     n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 ,
     n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 ,
     n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 ,
     n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 ,
     n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 ,
     n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 ,
     n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 ,
     n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 ,
     n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 ,
     n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 ,
     n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 ,
     n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 ,
     n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 ,
     n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 ,
     n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 ,
     n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 ,
     n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 ,
     n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 ,
     n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 ,
     n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 ,
     n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 ,
     n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 ,
     n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 ,
     n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 ,
     n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 ,
     n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 ,
     n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 ,
     n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 ,
     n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 ,
     n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 ,
     n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 ,
     n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 ,
     n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 ,
     n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 ,
     n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 ,
     n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 ,
     n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 ,
     n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 ,
     n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 ,
     n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 ,
     n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 ,
     n2355 , n2356 , n2357 , n2358 , n2359 , n2360 ;
buf ( n246 , n699 );
buf ( n249 , n2058 );
buf ( n251 , n9999 );
buf ( n247 , n2063 );
buf ( n243 , n2064 );
buf ( n244 , n2150 );
buf ( n245 , n9999 );
buf ( n250 , n2153 );
buf ( n256 , n2154 );
buf ( n255 , n2242 );
buf ( n252 , n9999 );
buf ( n253 , n2245 );
buf ( n257 , n2246 );
buf ( n254 , n2360 );
buf ( n248 , n9999 );
buf ( n530 , PI_PI_clock);
buf ( n531 , PI_PI_reset);
buf ( n532 , n6 );
buf ( n533 , n168 );
buf ( n534 , n233 );
buf ( n535 , n223 );
buf ( n536 , n85 );
buf ( n537 , PI_DFF_state_reg_Q);
buf ( n538 , n169 );
buf ( n539 , n95 );
buf ( n540 , n73 );
buf ( n541 , n93 );
buf ( n542 , n239 );
buf ( n543 , n99 );
buf ( n544 , n88 );
buf ( n545 , n174 );
buf ( n546 , n234 );
buf ( n547 , n2 );
buf ( n548 , n49 );
buf ( n549 , n108 );
buf ( n550 , n109 );
buf ( n551 , n61 );
buf ( n552 , n1 );
buf ( n553 , n198 );
buf ( n554 , n229 );
buf ( n555 , n113 );
buf ( n556 , n29 );
buf ( n557 , n143 );
buf ( n558 , n154 );
buf ( n559 , n151 );
buf ( n560 , n240 );
buf ( n561 , n64 );
buf ( n562 , n130 );
buf ( n563 , n48 );
buf ( n564 , n27 );
buf ( n565 , n30 );
buf ( n566 , n204 );
buf ( n567 , n19 );
buf ( n568 , n12 );
buf ( n569 , n105 );
buf ( n570 , n191 );
buf ( n571 , n206 );
buf ( n572 , n153 );
buf ( n573 , n179 );
buf ( n574 , n242 );
buf ( n575 , n180 );
buf ( n576 , n117 );
buf ( n577 , n101 );
buf ( n578 , n44 );
buf ( n579 , n33 );
buf ( n580 , n43 );
buf ( n581 , n173 );
buf ( n582 , n147 );
buf ( n583 , n120 );
buf ( n584 , n7 );
buf ( n585 , n196 );
buf ( n586 , n31 );
buf ( n587 , n82 );
buf ( n588 , n138 );
buf ( n589 , n25 );
buf ( n590 , n32 );
buf ( n591 , n228 );
buf ( n592 , n241 );
buf ( n593 , n189 );
buf ( n594 , n167 );
buf ( n595 , n76 );
buf ( n596 , n87 );
buf ( n597 , n127 );
buf ( n598 , n103 );
buf ( n599 , n152 );
buf ( n600 , n186 );
buf ( n601 , n129 );
buf ( n602 , n209 );
buf ( n603 , n146 );
buf ( n604 , n10 );
buf ( n605 , n83 );
buf ( n606 , n45 );
buf ( n607 , n157 );
buf ( n608 , n67 );
buf ( n609 , n115 );
buf ( n610 , n238 );
buf ( n611 , n94 );
buf ( n612 , n70 );
buf ( n613 , n3 );
buf ( n614 , n222 );
buf ( n615 , n11 );
buf ( n616 , n140 );
buf ( n617 , n177 );
buf ( n618 , n142 );
buf ( n619 , n216 );
buf ( n620 , n71 );
buf ( n621 , n116 );
buf ( n622 , n16 );
buf ( n623 , n205 );
buf ( n624 , n14 );
buf ( n625 , n53 );
buf ( n626 , n56 );
buf ( n627 , n195 );
buf ( n628 , n51 );
buf ( n629 , n21 );
buf ( n630 , n28 );
buf ( n631 , n207 );
buf ( n632 , n100 );
buf ( n633 , n59 );
buf ( n634 , n125 );
buf ( n635 , n96 );
buf ( n636 , n97 );
buf ( n637 , n200 );
buf ( n638 , n75 );
buf ( n639 , n26 );
buf ( n640 , n42 );
buf ( n641 , n72 );
buf ( n642 , n24 );
buf ( n643 , n54 );
buf ( n644 , n217 );
buf ( n645 , n5 );
buf ( n646 , n193 );
buf ( n647 , n35 );
buf ( n648 , n163 );
buf ( n649 , n60 );
buf ( n650 , n77 );
buf ( n651 , n92 );
buf ( n652 , n91 );
buf ( n653 , n185 );
buf ( n654 , n215 );
buf ( n655 , n156 );
buf ( n656 , n74 );
buf ( n657 , n212 );
buf ( n658 , n231 );
buf ( n659 , n34 );
buf ( n660 , n62 );
buf ( n661 , n237 );
buf ( n662 , n126 );
buf ( n663 , n172 );
buf ( n664 , n55 );
buf ( n665 , PI_DFF_B_reg_Q);
buf ( n666 , n122 );
buf ( n667 , n175 );
buf ( n668 , n178 );
buf ( n669 , n123 );
buf ( n670 , n37 );
buf ( n671 , n134 );
buf ( n672 , n194 );
buf ( n673 , n176 );
buf ( n674 , n213 );
buf ( n675 , n57 );
buf ( n676 , n81 );
buf ( n677 , n136 );
buf ( n678 , n40 );
buf ( n679 , n104 );
buf ( n680 , n135 );
buf ( n681 , n47 );
buf ( n682 , n39 );
buf ( n683 , n166 );
buf ( n684 , n79 );
buf ( n685 , n144 );
buf ( n686 , n208 );
buf ( n687 , n121 );
buf ( n688 , n23 );
buf ( n689 , n203 );
buf ( n690 , n235 );
buf ( n691 , n86 );
buf ( n692 , n9 );
buf ( n693 , n236 );
buf ( n694 , n8 );
buf ( n695 , n149 );
buf ( n696 , n165 );
buf ( n697 , n20 );
buf ( n698 , n530 );
buf ( n699 , n698 );
buf ( n700 , n569 );
not ( n701 , n700 );
not ( n702 , n701 );
not ( n703 , n702 );
buf ( n704 , n542 );
not ( n705 , n704 );
not ( n706 , n705 );
buf ( n707 , n543 );
not ( n708 , n707 );
not ( n709 , n708 );
not ( n710 , n709 );
not ( n711 , n710 );
nor ( n712 , n706 , n711 );
buf ( n713 , n545 );
not ( n714 , n713 );
not ( n715 , n714 );
not ( n716 , n715 );
not ( n717 , n716 );
buf ( n718 , n544 );
not ( n719 , n718 );
not ( n720 , n719 );
not ( n721 , n720 );
not ( n722 , n721 );
nor ( n723 , n717 , n722 );
nand ( n724 , n712 , n723 );
buf ( n725 , n538 );
not ( n726 , n725 );
buf ( n727 , n539 );
not ( n728 , n727 );
nand ( n729 , n726 , n728 );
not ( n730 , n729 );
buf ( n731 , n540 );
not ( n732 , n731 );
not ( n733 , n732 );
buf ( n734 , n541 );
not ( n735 , n734 );
not ( n736 , n735 );
nor ( n737 , n733 , n736 );
nand ( n738 , n730 , n737 );
or ( n739 , n724 , n738 );
not ( n740 , n739 );
buf ( n741 , n547 );
not ( n742 , n741 );
buf ( n743 , n546 );
not ( n744 , n743 );
not ( n745 , n744 );
not ( n746 , n745 );
nand ( n747 , n742 , n746 );
buf ( n748 , n549 );
not ( n749 , n748 );
buf ( n750 , n548 );
not ( n751 , n750 );
nand ( n752 , n749 , n751 );
nor ( n753 , n747 , n752 );
nand ( n754 , n740 , n753 );
buf ( n755 , n550 );
and ( n756 , n754 , n755 );
not ( n757 , n754 );
not ( n758 , n755 );
and ( n759 , n757 , n758 );
nor ( n760 , n756 , n759 );
not ( n761 , n760 );
not ( n762 , n761 );
not ( n763 , n762 );
or ( n764 , n703 , n763 );
nand ( n765 , n701 , n755 );
nand ( n766 , n764 , n765 );
not ( n767 , n766 );
not ( n768 , n767 );
not ( n769 , n701 );
not ( n770 , n769 );
buf ( n771 , n553 );
not ( n772 , n771 );
not ( n773 , n772 );
not ( n774 , n738 );
not ( n775 , n724 );
nand ( n776 , n774 , n775 );
not ( n777 , n776 );
buf ( n778 , n551 );
not ( n779 , n778 );
nand ( n780 , n779 , n758 );
buf ( n781 , n552 );
nor ( n782 , n780 , n781 );
and ( n783 , n753 , n782 );
nand ( n784 , n777 , n783 );
not ( n785 , n784 );
or ( n786 , n773 , n785 );
or ( n787 , n784 , n772 );
nand ( n788 , n786 , n787 );
not ( n789 , n788 );
or ( n790 , n770 , n789 );
nand ( n791 , n701 , n771 );
nand ( n792 , n790 , n791 );
nor ( n793 , n768 , n792 );
not ( n794 , n702 );
not ( n795 , n753 );
nor ( n796 , n795 , n755 );
nand ( n797 , n777 , n796 );
and ( n798 , n797 , n778 );
not ( n799 , n797 );
and ( n800 , n799 , n779 );
nor ( n801 , n798 , n800 );
not ( n802 , n801 );
or ( n803 , n794 , n802 );
nand ( n804 , n701 , n778 );
nand ( n805 , n803 , n804 );
not ( n806 , n805 );
not ( n807 , n806 );
not ( n808 , n702 );
nor ( n809 , n795 , n780 );
nand ( n810 , n777 , n809 );
and ( n811 , n810 , n781 );
not ( n812 , n810 );
not ( n813 , n781 );
and ( n814 , n812 , n813 );
nor ( n815 , n811 , n814 );
not ( n816 , n815 );
or ( n817 , n808 , n816 );
nand ( n818 , n701 , n781 );
nand ( n819 , n817 , n818 );
nor ( n820 , n807 , n819 );
not ( n821 , n702 );
not ( n822 , n751 );
nor ( n823 , n822 , n747 );
nand ( n824 , n740 , n823 );
not ( n825 , n749 );
and ( n826 , n824 , n825 );
not ( n827 , n824 );
and ( n828 , n827 , n749 );
nor ( n829 , n826 , n828 );
not ( n830 , n829 );
not ( n831 , n830 );
not ( n832 , n831 );
or ( n833 , n821 , n832 );
nand ( n834 , n701 , n748 );
nand ( n835 , n833 , n834 );
not ( n836 , n835 );
not ( n837 , n745 );
not ( n838 , n701 );
or ( n839 , n837 , n838 );
not ( n840 , n745 );
not ( n841 , n740 );
or ( n842 , n840 , n841 );
or ( n843 , n777 , n745 );
nand ( n844 , n842 , n843 );
nand ( n845 , n844 , n700 );
nand ( n846 , n839 , n845 );
and ( n847 , n701 , n715 );
not ( n848 , n701 );
not ( n849 , n717 );
not ( n850 , n849 );
not ( n851 , n710 );
nor ( n852 , n851 , n706 );
not ( n853 , n852 );
nor ( n854 , n853 , n722 );
not ( n855 , n736 );
not ( n856 , n727 );
not ( n857 , n725 );
not ( n858 , n733 );
and ( n859 , n855 , n856 , n857 , n858 );
nand ( n860 , n854 , n859 );
not ( n861 , n860 );
or ( n862 , n850 , n861 );
nand ( n863 , n859 , n854 );
or ( n864 , n863 , n849 );
nand ( n865 , n862 , n864 );
and ( n866 , n848 , n865 );
nor ( n867 , n847 , n866 );
not ( n868 , n867 );
not ( n869 , n868 );
and ( n870 , n701 , n709 );
not ( n871 , n701 );
not ( n872 , n851 );
not ( n873 , n872 );
not ( n874 , n706 );
nand ( n875 , n859 , n874 );
not ( n876 , n875 );
or ( n877 , n873 , n876 );
nand ( n878 , n859 , n874 );
or ( n879 , n878 , n872 );
nand ( n880 , n877 , n879 );
and ( n881 , n871 , n880 );
nor ( n882 , n870 , n881 );
not ( n883 , n882 );
not ( n884 , n883 );
nand ( n885 , n869 , n884 );
nor ( n886 , n846 , n885 );
and ( n887 , n836 , n886 );
nand ( n888 , n793 , n820 , n887 );
not ( n889 , n888 );
not ( n890 , n702 );
not ( n891 , n751 );
not ( n892 , n747 );
nand ( n893 , n892 , n740 );
not ( n894 , n893 );
or ( n895 , n891 , n894 );
or ( n896 , n893 , n751 );
nand ( n897 , n895 , n896 );
not ( n898 , n897 );
not ( n899 , n898 );
not ( n900 , n899 );
or ( n901 , n890 , n900 );
nand ( n902 , n701 , n750 );
nand ( n903 , n901 , n902 );
not ( n904 , n903 );
and ( n905 , n701 , n720 );
not ( n906 , n701 );
not ( n907 , n722 );
not ( n908 , n907 );
nand ( n909 , n859 , n852 );
not ( n910 , n909 );
or ( n911 , n908 , n910 );
nand ( n912 , n859 , n852 );
or ( n913 , n912 , n907 );
nand ( n914 , n911 , n913 );
and ( n915 , n906 , n914 );
nor ( n916 , n905 , n915 );
not ( n917 , n916 );
not ( n918 , n700 );
and ( n919 , n918 , n736 );
not ( n920 , n918 );
not ( n921 , n858 );
nor ( n922 , n921 , n729 );
and ( n923 , n922 , n855 );
not ( n924 , n922 );
not ( n925 , n855 );
and ( n926 , n924 , n925 );
nor ( n927 , n923 , n926 );
and ( n928 , n920 , n927 );
nor ( n929 , n919 , n928 );
not ( n930 , n929 );
not ( n931 , n930 );
not ( n932 , n874 );
not ( n933 , n738 );
or ( n934 , n932 , n933 );
or ( n935 , n874 , n738 );
nand ( n936 , n934 , n935 );
and ( n937 , n700 , n936 );
not ( n938 , n700 );
and ( n939 , n938 , n706 );
nor ( n940 , n937 , n939 );
not ( n941 , n940 );
not ( n942 , n941 );
not ( n943 , n700 );
not ( n944 , n858 );
not ( n945 , n729 );
or ( n946 , n944 , n945 );
or ( n947 , n729 , n858 );
nand ( n948 , n946 , n947 );
not ( n949 , n948 );
or ( n950 , n943 , n949 );
not ( n951 , n700 );
nand ( n952 , n951 , n733 );
nand ( n953 , n950 , n952 );
not ( n954 , n700 );
not ( n955 , n856 );
not ( n956 , n955 );
not ( n957 , n857 );
or ( n958 , n956 , n957 );
or ( n959 , n955 , n857 );
nand ( n960 , n958 , n959 );
not ( n961 , n960 );
or ( n962 , n954 , n961 );
nand ( n963 , n951 , n727 );
nand ( n964 , n962 , n963 );
not ( n965 , n964 );
not ( n966 , n725 );
nand ( n967 , n965 , n966 );
nor ( n968 , n953 , n967 );
nand ( n969 , n931 , n942 , n968 );
nor ( n970 , n917 , n969 );
and ( n971 , n904 , n970 );
not ( n972 , n702 );
nand ( n973 , n777 , n746 );
and ( n974 , n973 , n741 );
not ( n975 , n973 );
and ( n976 , n975 , n742 );
nor ( n977 , n974 , n976 );
not ( n978 , n977 );
or ( n979 , n972 , n978 );
nand ( n980 , n701 , n741 );
nand ( n981 , n979 , n980 );
not ( n982 , n981 );
not ( n983 , n702 );
nand ( n984 , n751 , n721 );
nand ( n985 , n749 , n716 );
nor ( n986 , n984 , n985 );
not ( n987 , n729 );
nor ( n988 , n745 , n706 );
nand ( n989 , n986 , n987 , n988 );
nor ( n990 , n733 , n755 );
nor ( n991 , n778 , n736 );
nor ( n992 , n771 , n781 );
nor ( n993 , n741 , n709 );
nand ( n994 , n990 , n991 , n992 , n993 );
nor ( n995 , n989 , n994 );
buf ( n996 , n555 );
buf ( n997 , n554 );
not ( n998 , n997 );
not ( n999 , n998 );
nor ( n1000 , n996 , n999 );
not ( n1001 , n1000 );
not ( n1002 , n1001 );
nand ( n1003 , n995 , n1002 );
buf ( n1004 , n556 );
not ( n1005 , n1004 );
not ( n1006 , n1005 );
and ( n1007 , n1003 , n1006 );
not ( n1008 , n1003 );
not ( n1009 , n1006 );
and ( n1010 , n1008 , n1009 );
nor ( n1011 , n1007 , n1010 );
not ( n1012 , n1011 );
or ( n1013 , n983 , n1012 );
nand ( n1014 , n701 , n1006 );
nand ( n1015 , n1013 , n1014 );
not ( n1016 , n1015 );
and ( n1017 , n982 , n1016 );
not ( n1018 , n702 );
not ( n1019 , n995 );
nor ( n1020 , n1019 , n999 );
or ( n1021 , n1020 , n996 );
nand ( n1022 , n991 , n992 , n988 , n993 );
not ( n1023 , n1022 );
not ( n1024 , n986 );
not ( n1025 , n999 );
nand ( n1026 , n1025 , n857 , n856 , n996 );
not ( n1027 , n990 );
nor ( n1028 , n1024 , n1026 , n1027 );
nand ( n1029 , n1023 , n1028 );
nand ( n1030 , n1021 , n1029 );
not ( n1031 , n1030 );
or ( n1032 , n1018 , n1031 );
nand ( n1033 , n701 , n996 );
nand ( n1034 , n1032 , n1033 );
not ( n1035 , n1034 );
not ( n1036 , n999 );
not ( n1037 , n701 );
or ( n1038 , n1036 , n1037 );
not ( n1039 , n999 );
not ( n1040 , n995 );
or ( n1041 , n1039 , n1040 );
or ( n1042 , n995 , n999 );
nand ( n1043 , n1041 , n1042 );
nand ( n1044 , n1043 , n700 );
nand ( n1045 , n1038 , n1044 );
not ( n1046 , n1045 );
and ( n1047 , n1035 , n1046 );
nand ( n1048 , n971 , n1017 , n1047 );
not ( n1049 , n1048 );
and ( n1050 , n889 , n1049 );
not ( n1051 , n1019 );
buf ( n1052 , n563 );
buf ( n1053 , n562 );
nor ( n1054 , n1052 , n1053 );
buf ( n1055 , n564 );
buf ( n1056 , n565 );
nor ( n1057 , n1055 , n1056 );
nand ( n1058 , n1054 , n1057 );
not ( n1059 , n1058 );
buf ( n1060 , n567 );
buf ( n1061 , n566 );
or ( n1062 , n1060 , n1061 );
buf ( n1063 , n568 );
nor ( n1064 , n1062 , n1063 );
nand ( n1065 , n1059 , n1064 );
buf ( n1066 , n559 );
not ( n1067 , n1066 );
not ( n1068 , n1067 );
buf ( n1069 , n557 );
nor ( n1070 , n1068 , n1069 );
buf ( n1071 , n560 );
nor ( n1072 , n1071 , n999 );
buf ( n1073 , n561 );
nor ( n1074 , n1073 , n996 );
buf ( n1075 , n558 );
not ( n1076 , n1075 );
not ( n1077 , n1076 );
nor ( n1078 , n1077 , n1006 );
nand ( n1079 , n1070 , n1072 , n1074 , n1078 );
nor ( n1080 , n1065 , n1079 );
nand ( n1081 , n1051 , n1080 );
and ( n1082 , n1081 , n700 );
not ( n1083 , n1081 );
not ( n1084 , n700 );
and ( n1085 , n1083 , n1084 );
nor ( n1086 , n1082 , n1085 );
nand ( n1087 , n1086 , n702 );
not ( n1088 , n1087 );
not ( n1089 , n1088 );
nor ( n1090 , n1050 , n1089 );
not ( n1091 , n1069 );
not ( n1092 , n701 );
or ( n1093 , n1091 , n1092 );
nor ( n1094 , n1001 , n1006 );
nand ( n1095 , n995 , n1094 );
xor ( n1096 , n1095 , n1069 );
nand ( n1097 , n1096 , n702 );
nand ( n1098 , n1093 , n1097 );
not ( n1099 , n1098 );
not ( n1100 , n769 );
nor ( n1101 , n1006 , n1069 );
nand ( n1102 , n1000 , n1101 );
not ( n1103 , n1102 );
nand ( n1104 , n1103 , n995 );
and ( n1105 , n1104 , n1077 );
not ( n1106 , n1104 );
not ( n1107 , n1077 );
and ( n1108 , n1106 , n1107 );
nor ( n1109 , n1105 , n1108 );
not ( n1110 , n1109 );
or ( n1111 , n1100 , n1110 );
not ( n1112 , n702 );
nand ( n1113 , n1112 , n1077 );
nand ( n1114 , n1111 , n1113 );
not ( n1115 , n1114 );
not ( n1116 , n769 );
nor ( n1117 , n1102 , n1077 );
nand ( n1118 , n995 , n1117 );
xor ( n1119 , n1118 , n1068 );
not ( n1120 , n1119 );
or ( n1121 , n1116 , n1120 );
nand ( n1122 , n701 , n1068 );
nand ( n1123 , n1121 , n1122 );
not ( n1124 , n1123 );
not ( n1125 , n769 );
nor ( n1126 , n1068 , n1077 );
not ( n1127 , n1126 );
nor ( n1128 , n1127 , n1102 );
nand ( n1129 , n995 , n1128 );
not ( n1130 , n1071 );
xnor ( n1131 , n1129 , n1130 );
not ( n1132 , n1131 );
or ( n1133 , n1125 , n1132 );
nand ( n1134 , n701 , n1071 );
nand ( n1135 , n1133 , n1134 );
not ( n1136 , n1135 );
and ( n1137 , n1099 , n1115 , n1124 , n1136 );
not ( n1138 , n702 );
nand ( n1139 , n1126 , n1130 );
nor ( n1140 , n1102 , n1139 );
nand ( n1141 , n995 , n1140 );
not ( n1142 , n1073 );
xnor ( n1143 , n1141 , n1142 );
not ( n1144 , n1143 );
or ( n1145 , n1138 , n1144 );
nand ( n1146 , n1112 , n1073 );
nand ( n1147 , n1145 , n1146 );
not ( n1148 , n769 );
nor ( n1149 , n1079 , n1053 );
nand ( n1150 , n995 , n1149 );
not ( n1151 , n1052 );
xnor ( n1152 , n1150 , n1151 );
not ( n1153 , n1152 );
or ( n1154 , n1148 , n1153 );
nand ( n1155 , n701 , n1052 );
nand ( n1156 , n1154 , n1155 );
not ( n1157 , n769 );
not ( n1158 , n1053 );
not ( n1159 , n1158 );
not ( n1160 , n1079 );
nand ( n1161 , n1160 , n995 );
not ( n1162 , n1161 );
or ( n1163 , n1159 , n1162 );
or ( n1164 , n1161 , n1158 );
nand ( n1165 , n1163 , n1164 );
not ( n1166 , n1165 );
or ( n1167 , n1157 , n1166 );
nand ( n1168 , n701 , n1053 );
nand ( n1169 , n1167 , n1168 );
or ( n1170 , n1147 , n1156 , n1169 );
not ( n1171 , n702 );
not ( n1172 , n1054 );
nor ( n1173 , n1172 , n1079 );
nand ( n1174 , n995 , n1173 );
not ( n1175 , n1055 );
xnor ( n1176 , n1174 , n1175 );
not ( n1177 , n1176 );
not ( n1178 , n1177 );
not ( n1179 , n1178 );
or ( n1180 , n1171 , n1179 );
nand ( n1181 , n701 , n1055 );
nand ( n1182 , n1180 , n1181 );
nor ( n1183 , n1170 , n1182 );
and ( n1184 , n1137 , n1183 );
nor ( n1185 , n1184 , n1089 );
nor ( n1186 , n1090 , n1185 );
not ( n1187 , n1186 );
not ( n1188 , n1056 );
not ( n1189 , n1112 );
or ( n1190 , n1188 , n1189 );
nand ( n1191 , n1054 , n1175 );
nor ( n1192 , n1079 , n1191 );
nand ( n1193 , n995 , n1192 );
xor ( n1194 , n1193 , n1056 );
nand ( n1195 , n1194 , n702 );
nand ( n1196 , n1190 , n1195 );
nand ( n1197 , n1187 , n1196 );
and ( n1198 , n701 , n1061 );
not ( n1199 , n701 );
nor ( n1200 , n1079 , n1058 );
nand ( n1201 , n995 , n1200 );
not ( n1202 , n1061 );
not ( n1203 , n1202 );
and ( n1204 , n1201 , n1203 );
not ( n1205 , n1201 );
and ( n1206 , n1205 , n1202 );
nor ( n1207 , n1204 , n1206 );
and ( n1208 , n1199 , n1207 );
nor ( n1209 , n1198 , n1208 );
not ( n1210 , n1209 );
not ( n1211 , n1210 );
and ( n1212 , n1197 , n1211 );
not ( n1213 , n1197 );
and ( n1214 , n1213 , n1210 );
nor ( n1215 , n1212 , n1214 );
not ( n1216 , n1215 );
not ( n1217 , n1216 );
buf ( n1218 , n572 );
not ( n1219 , n1218 );
not ( n1220 , n1219 );
not ( n1221 , n1220 );
nand ( n1222 , n1044 , n867 );
not ( n1223 , n1222 );
not ( n1224 , n845 );
nand ( n1225 , n916 , n882 );
nor ( n1226 , n1224 , n1225 );
nor ( n1227 , n788 , n1152 );
nand ( n1228 , n1223 , n1226 , n1227 );
nor ( n1229 , n1143 , n725 );
nand ( n1230 , n1229 , n1177 , n898 , n761 );
nor ( n1231 , n1228 , n1230 );
nor ( n1232 , n1165 , n1119 );
nor ( n1233 , n1109 , n1011 );
nand ( n1234 , n1209 , n1195 , n1232 , n1233 );
not ( n1235 , n1234 );
not ( n1236 , n977 );
nor ( n1237 , n953 , n964 );
and ( n1238 , n940 , n929 , n1237 );
nand ( n1239 , n1097 , n1236 , n830 , n1238 );
nor ( n1240 , n801 , n815 );
nor ( n1241 , n1131 , n1030 );
nand ( n1242 , n1240 , n1241 );
nor ( n1243 , n1239 , n1242 );
nand ( n1244 , n1231 , n1235 , n1243 );
nand ( n1245 , n1244 , n1088 );
nand ( n1246 , n1059 , n1202 );
nor ( n1247 , n1246 , n1079 );
nand ( n1248 , n1051 , n1247 );
xor ( n1249 , n1248 , n1060 );
and ( n1250 , n1249 , n769 );
and ( n1251 , n701 , n1060 );
nor ( n1252 , n1250 , n1251 );
and ( n1253 , n1245 , n1252 );
not ( n1254 , n1245 );
not ( n1255 , n1252 );
and ( n1256 , n1254 , n1255 );
nor ( n1257 , n1253 , n1256 );
not ( n1258 , n1257 );
not ( n1259 , n1258 );
nor ( n1260 , n1252 , n1087 );
nand ( n1261 , n1244 , n1260 );
not ( n1262 , n1261 );
not ( n1263 , n1062 );
nand ( n1264 , n1263 , n1059 );
nor ( n1265 , n1264 , n1079 );
nand ( n1266 , n1051 , n1265 );
xor ( n1267 , n1266 , n1063 );
nand ( n1268 , n1267 , n769 );
nand ( n1269 , n701 , n1063 );
nand ( n1270 , n1268 , n1269 );
not ( n1271 , n1270 );
and ( n1272 , n1262 , n1271 );
and ( n1273 , n1261 , n1270 );
nor ( n1274 , n1272 , n1273 );
not ( n1275 , n1274 );
nand ( n1276 , n1259 , n1275 );
not ( n1277 , n1276 );
not ( n1278 , n1277 );
or ( n1279 , n1221 , n1278 );
not ( n1280 , n1274 );
nand ( n1281 , n1280 , n1258 );
not ( n1282 , n1281 );
buf ( n1283 , n666 );
nand ( n1284 , n1282 , n1283 );
nand ( n1285 , n1279 , n1284 );
buf ( n1286 , n601 );
not ( n1287 , n1286 );
not ( n1288 , n1257 );
nor ( n1289 , n1275 , n1288 );
not ( n1290 , n1289 );
not ( n1291 , n1290 );
not ( n1292 , n1291 );
or ( n1293 , n1287 , n1292 );
nand ( n1294 , n1274 , n1258 );
not ( n1295 , n1294 );
buf ( n1296 , n633 );
not ( n1297 , n1296 );
not ( n1298 , n1297 );
nand ( n1299 , n1295 , n1298 );
nand ( n1300 , n1293 , n1299 );
nor ( n1301 , n1285 , n1300 );
not ( n1302 , n1301 );
and ( n1303 , n1217 , n1302 );
not ( n1304 , n1217 );
buf ( n1305 , n574 );
not ( n1306 , n1305 );
not ( n1307 , n1277 );
or ( n1308 , n1306 , n1307 );
buf ( n1309 , n668 );
nand ( n1310 , n1282 , n1309 );
nand ( n1311 , n1308 , n1310 );
buf ( n1312 , n635 );
not ( n1313 , n1312 );
not ( n1314 , n1313 );
not ( n1315 , n1314 );
not ( n1316 , n1295 );
or ( n1317 , n1315 , n1316 );
buf ( n1318 , n603 );
not ( n1319 , n1318 );
not ( n1320 , n1319 );
nand ( n1321 , n1291 , n1320 );
nand ( n1322 , n1317 , n1321 );
nor ( n1323 , n1311 , n1322 );
not ( n1324 , n1323 );
not ( n1325 , n1324 );
not ( n1326 , n1274 );
nand ( n1327 , n1326 , n1288 );
not ( n1328 , n1327 );
buf ( n1329 , n671 );
nand ( n1330 , n1328 , n1329 );
nor ( n1331 , n1288 , n1280 );
not ( n1332 , n1331 );
not ( n1333 , n1332 );
buf ( n1334 , n606 );
nand ( n1335 , n1333 , n1334 );
nand ( n1336 , n1326 , n1259 );
not ( n1337 , n1336 );
buf ( n1338 , n577 );
nand ( n1339 , n1337 , n1338 );
nand ( n1340 , n1274 , n1288 );
not ( n1341 , n1340 );
buf ( n1342 , n638 );
not ( n1343 , n1342 );
not ( n1344 , n1343 );
nand ( n1345 , n1341 , n1344 );
nand ( n1346 , n1330 , n1335 , n1339 , n1345 );
not ( n1347 , n1281 );
buf ( n1348 , n674 );
nand ( n1349 , n1347 , n1348 );
buf ( n1350 , n609 );
nand ( n1351 , n1289 , n1350 );
not ( n1352 , n1276 );
buf ( n1353 , n580 );
nand ( n1354 , n1352 , n1353 );
buf ( n1355 , n641 );
nand ( n1356 , n1295 , n1355 );
nand ( n1357 , n1349 , n1351 , n1354 , n1356 );
not ( n1358 , n1340 );
buf ( n1359 , n637 );
not ( n1360 , n1359 );
not ( n1361 , n1360 );
nand ( n1362 , n1358 , n1361 );
not ( n1363 , n1332 );
buf ( n1364 , n605 );
nand ( n1365 , n1363 , n1364 );
not ( n1366 , n1336 );
buf ( n1367 , n576 );
nand ( n1368 , n1366 , n1367 );
not ( n1369 , n1327 );
buf ( n1370 , n670 );
nand ( n1371 , n1369 , n1370 );
nand ( n1372 , n1362 , n1365 , n1368 , n1371 );
buf ( n1373 , n675 );
nand ( n1374 , n1347 , n1373 );
buf ( n1375 , n610 );
nand ( n1376 , n1289 , n1375 );
not ( n1377 , n1276 );
buf ( n1378 , n581 );
nand ( n1379 , n1377 , n1378 );
buf ( n1380 , n642 );
not ( n1381 , n1380 );
not ( n1382 , n1381 );
nand ( n1383 , n1295 , n1382 );
nand ( n1384 , n1374 , n1376 , n1379 , n1383 );
nand ( n1385 , n1346 , n1357 , n1372 , n1384 );
not ( n1386 , n1281 );
not ( n1387 , n1386 );
buf ( n1388 , n679 );
not ( n1389 , n1388 );
nor ( n1390 , n1387 , n1389 );
not ( n1391 , n1289 );
buf ( n1392 , n614 );
not ( n1393 , n1392 );
nor ( n1394 , n1391 , n1393 );
nor ( n1395 , n1390 , n1394 );
not ( n1396 , n1276 );
buf ( n1397 , n585 );
and ( n1398 , n1396 , n1397 );
not ( n1399 , n1295 );
buf ( n1400 , n646 );
not ( n1401 , n1400 );
not ( n1402 , n1401 );
not ( n1403 , n1402 );
nor ( n1404 , n1399 , n1403 );
nor ( n1405 , n1398 , n1404 );
nand ( n1406 , n1395 , n1405 );
not ( n1407 , n1281 );
buf ( n1408 , n678 );
nand ( n1409 , n1407 , n1408 );
buf ( n1410 , n613 );
nand ( n1411 , n1289 , n1410 );
not ( n1412 , n1276 );
buf ( n1413 , n584 );
nand ( n1414 , n1412 , n1413 );
not ( n1415 , n1294 );
buf ( n1416 , n645 );
not ( n1417 , n1416 );
not ( n1418 , n1417 );
nand ( n1419 , n1415 , n1418 );
nand ( n1420 , n1409 , n1411 , n1414 , n1419 );
nand ( n1421 , n1406 , n1420 );
nor ( n1422 , n1385 , n1421 );
buf ( n1423 , n677 );
nand ( n1424 , n1407 , n1423 );
buf ( n1425 , n612 );
nand ( n1426 , n1289 , n1425 );
buf ( n1427 , n583 );
nand ( n1428 , n1412 , n1427 );
not ( n1429 , n1294 );
buf ( n1430 , n644 );
not ( n1431 , n1430 );
not ( n1432 , n1431 );
nand ( n1433 , n1429 , n1432 );
nand ( n1434 , n1424 , n1426 , n1428 , n1433 );
buf ( n1435 , n582 );
nand ( n1436 , n1412 , n1435 );
buf ( n1437 , n676 );
nand ( n1438 , n1407 , n1437 );
buf ( n1439 , n611 );
nand ( n1440 , n1289 , n1439 );
buf ( n1441 , n643 );
not ( n1442 , n1441 );
not ( n1443 , n1442 );
nand ( n1444 , n1415 , n1443 );
nand ( n1445 , n1436 , n1438 , n1440 , n1444 );
nand ( n1446 , n1434 , n1445 );
buf ( n1447 , n587 );
nand ( n1448 , n1277 , n1447 );
buf ( n1449 , n681 );
nand ( n1450 , n1369 , n1449 );
not ( n1451 , n1331 );
not ( n1452 , n1451 );
buf ( n1453 , n616 );
nand ( n1454 , n1452 , n1453 );
buf ( n1455 , n648 );
not ( n1456 , n1455 );
not ( n1457 , n1456 );
nand ( n1458 , n1358 , n1457 );
nand ( n1459 , n1448 , n1450 , n1454 , n1458 );
buf ( n1460 , n680 );
nand ( n1461 , n1386 , n1460 );
buf ( n1462 , n615 );
nand ( n1463 , n1289 , n1462 );
buf ( n1464 , n586 );
nand ( n1465 , n1366 , n1464 );
buf ( n1466 , n647 );
not ( n1467 , n1466 );
not ( n1468 , n1467 );
nand ( n1469 , n1358 , n1468 );
nand ( n1470 , n1461 , n1463 , n1465 , n1469 );
nand ( n1471 , n1459 , n1470 );
nor ( n1472 , n1446 , n1471 );
buf ( n1473 , n672 );
nand ( n1474 , n1369 , n1473 );
buf ( n1475 , n607 );
nand ( n1476 , n1452 , n1475 );
buf ( n1477 , n578 );
nand ( n1478 , n1366 , n1477 );
buf ( n1479 , n639 );
not ( n1480 , n1479 );
not ( n1481 , n1480 );
nand ( n1482 , n1295 , n1481 );
nand ( n1483 , n1474 , n1476 , n1478 , n1482 );
not ( n1484 , n1327 );
buf ( n1485 , n669 );
nand ( n1486 , n1484 , n1485 );
not ( n1487 , n1451 );
buf ( n1488 , n604 );
nand ( n1489 , n1487 , n1488 );
not ( n1490 , n1336 );
buf ( n1491 , n575 );
nand ( n1492 , n1490 , n1491 );
not ( n1493 , n1340 );
buf ( n1494 , n636 );
not ( n1495 , n1494 );
not ( n1496 , n1495 );
nand ( n1497 , n1493 , n1496 );
nand ( n1498 , n1486 , n1489 , n1492 , n1497 );
nand ( n1499 , n1483 , n1498 );
buf ( n1500 , n608 );
nand ( n1501 , n1289 , n1500 );
buf ( n1502 , n673 );
nand ( n1503 , n1347 , n1502 );
buf ( n1504 , n579 );
nand ( n1505 , n1377 , n1504 );
not ( n1506 , n1294 );
buf ( n1507 , n640 );
not ( n1508 , n1507 );
not ( n1509 , n1508 );
nand ( n1510 , n1506 , n1509 );
nand ( n1511 , n1501 , n1503 , n1505 , n1510 );
nand ( n1512 , n1511 , n1277 );
nor ( n1513 , n1499 , n1512 );
and ( n1514 , n1422 , n1472 , n1513 );
not ( n1515 , n1391 );
buf ( n1516 , n627 );
not ( n1517 , n1516 );
not ( n1518 , n1517 );
and ( n1519 , n1515 , n1518 );
not ( n1520 , n1407 );
buf ( n1521 , n692 );
not ( n1522 , n1521 );
not ( n1523 , n1522 );
not ( n1524 , n1523 );
nor ( n1525 , n1520 , n1524 );
nor ( n1526 , n1519 , n1525 );
buf ( n1527 , n598 );
not ( n1528 , n1527 );
not ( n1529 , n1528 );
and ( n1530 , n1396 , n1529 );
not ( n1531 , n1295 );
buf ( n1532 , n659 );
not ( n1533 , n1532 );
not ( n1534 , n1533 );
not ( n1535 , n1534 );
nor ( n1536 , n1531 , n1535 );
nor ( n1537 , n1530 , n1536 );
nand ( n1538 , n1526 , n1537 );
buf ( n1539 , n693 );
not ( n1540 , n1539 );
not ( n1541 , n1540 );
not ( n1542 , n1541 );
nor ( n1543 , n1281 , n1542 );
buf ( n1544 , n628 );
not ( n1545 , n1544 );
not ( n1546 , n1545 );
not ( n1547 , n1546 );
nor ( n1548 , n1391 , n1547 );
nor ( n1549 , n1543 , n1548 );
buf ( n1550 , n660 );
not ( n1551 , n1550 );
nor ( n1552 , n1399 , n1551 );
buf ( n1553 , n599 );
not ( n1554 , n1553 );
not ( n1555 , n1554 );
not ( n1556 , n1555 );
nor ( n1557 , n1276 , n1556 );
nor ( n1558 , n1552 , n1557 );
nand ( n1559 , n1549 , n1558 );
nand ( n1560 , n1538 , n1559 );
buf ( n1561 , n694 );
not ( n1562 , n1561 );
not ( n1563 , n1562 );
not ( n1564 , n1563 );
nor ( n1565 , n1281 , n1564 );
buf ( n1566 , n629 );
not ( n1567 , n1566 );
not ( n1568 , n1567 );
not ( n1569 , n1568 );
nor ( n1570 , n1391 , n1569 );
nor ( n1571 , n1565 , n1570 );
buf ( n1572 , n600 );
not ( n1573 , n1572 );
not ( n1574 , n1573 );
and ( n1575 , n1396 , n1574 );
buf ( n1576 , n661 );
not ( n1577 , n1576 );
not ( n1578 , n1577 );
not ( n1579 , n1578 );
nor ( n1580 , n1531 , n1579 );
nor ( n1581 , n1575 , n1580 );
nand ( n1582 , n1571 , n1581 );
buf ( n1583 , n662 );
not ( n1584 , n1583 );
not ( n1585 , n1584 );
nand ( n1586 , n1415 , n1585 );
not ( n1587 , n1391 );
buf ( n1588 , n630 );
not ( n1589 , n1588 );
not ( n1590 , n1589 );
nand ( n1591 , n1587 , n1590 );
buf ( n1592 , n695 );
not ( n1593 , n1592 );
not ( n1594 , n1593 );
nand ( n1595 , n1407 , n1594 );
nand ( n1596 , n1586 , n1591 , n1595 );
nand ( n1597 , n1582 , n1596 );
nor ( n1598 , n1560 , n1597 );
not ( n1599 , n1387 );
buf ( n1600 , n689 );
not ( n1601 , n1600 );
not ( n1602 , n1601 );
not ( n1603 , n1602 );
not ( n1604 , n1603 );
and ( n1605 , n1599 , n1604 );
buf ( n1606 , n624 );
not ( n1607 , n1606 );
not ( n1608 , n1607 );
and ( n1609 , n1291 , n1608 );
nor ( n1610 , n1605 , n1609 );
not ( n1611 , n1294 );
buf ( n1612 , n656 );
not ( n1613 , n1612 );
not ( n1614 , n1613 );
not ( n1615 , n1614 );
not ( n1616 , n1615 );
and ( n1617 , n1611 , n1616 );
not ( n1618 , n1276 );
buf ( n1619 , n595 );
and ( n1620 , n1618 , n1619 );
nor ( n1621 , n1617 , n1620 );
nand ( n1622 , n1610 , n1621 );
buf ( n1623 , n594 );
not ( n1624 , n1623 );
not ( n1625 , n1624 );
not ( n1626 , n1625 );
nor ( n1627 , n1276 , n1626 );
not ( n1628 , n1289 );
buf ( n1629 , n623 );
not ( n1630 , n1629 );
not ( n1631 , n1630 );
not ( n1632 , n1631 );
nor ( n1633 , n1628 , n1632 );
nor ( n1634 , n1627 , n1633 );
buf ( n1635 , n688 );
not ( n1636 , n1635 );
not ( n1637 , n1636 );
not ( n1638 , n1637 );
nor ( n1639 , n1281 , n1638 );
buf ( n1640 , n655 );
not ( n1641 , n1640 );
not ( n1642 , n1641 );
not ( n1643 , n1642 );
nor ( n1644 , n1294 , n1643 );
nor ( n1645 , n1639 , n1644 );
nand ( n1646 , n1634 , n1645 );
nand ( n1647 , n1622 , n1646 );
buf ( n1648 , n652 );
not ( n1649 , n1648 );
not ( n1650 , n1649 );
nand ( n1651 , n1295 , n1650 );
buf ( n1652 , n685 );
nand ( n1653 , n1386 , n1652 );
buf ( n1654 , n620 );
nand ( n1655 , n1291 , n1654 );
buf ( n1656 , n591 );
nand ( n1657 , n1396 , n1656 );
nand ( n1658 , n1651 , n1653 , n1655 , n1657 );
not ( n1659 , n1347 );
not ( n1660 , n1659 );
buf ( n1661 , n684 );
not ( n1662 , n1661 );
not ( n1663 , n1662 );
and ( n1664 , n1660 , n1663 );
not ( n1665 , n1628 );
buf ( n1666 , n619 );
and ( n1667 , n1665 , n1666 );
nor ( n1668 , n1664 , n1667 );
buf ( n1669 , n651 );
not ( n1670 , n1669 );
not ( n1671 , n1670 );
not ( n1672 , n1671 );
nor ( n1673 , n1294 , n1672 );
buf ( n1674 , n590 );
not ( n1675 , n1674 );
nor ( n1676 , n1276 , n1675 );
nor ( n1677 , n1673 , n1676 );
nand ( n1678 , n1668 , n1677 );
nand ( n1679 , n1658 , n1678 );
nor ( n1680 , n1647 , n1679 );
nand ( n1681 , n1598 , n1680 );
buf ( n1682 , n650 );
not ( n1683 , n1682 );
not ( n1684 , n1683 );
nand ( n1685 , n1415 , n1684 );
buf ( n1686 , n618 );
nand ( n1687 , n1665 , n1686 );
not ( n1688 , n1659 );
buf ( n1689 , n683 );
nand ( n1690 , n1688 , n1689 );
buf ( n1691 , n589 );
nand ( n1692 , n1277 , n1691 );
nand ( n1693 , n1685 , n1687 , n1690 , n1692 );
buf ( n1694 , n649 );
not ( n1695 , n1694 );
not ( n1696 , n1695 );
nand ( n1697 , n1415 , n1696 );
buf ( n1698 , n682 );
nand ( n1699 , n1688 , n1698 );
buf ( n1700 , n617 );
nand ( n1701 , n1291 , n1700 );
buf ( n1702 , n588 );
nand ( n1703 , n1277 , n1702 );
nand ( n1704 , n1697 , n1699 , n1701 , n1703 );
nand ( n1705 , n1693 , n1704 );
not ( n1706 , n1705 );
not ( n1707 , n1281 );
buf ( n1708 , n691 );
not ( n1709 , n1708 );
not ( n1710 , n1709 );
not ( n1711 , n1710 );
not ( n1712 , n1711 );
and ( n1713 , n1707 , n1712 );
buf ( n1714 , n626 );
not ( n1715 , n1714 );
not ( n1716 , n1715 );
and ( n1717 , n1515 , n1716 );
nor ( n1718 , n1713 , n1717 );
buf ( n1719 , n658 );
not ( n1720 , n1719 );
not ( n1721 , n1720 );
not ( n1722 , n1721 );
nor ( n1723 , n1399 , n1722 );
not ( n1724 , n1396 );
buf ( n1725 , n597 );
not ( n1726 , n1725 );
nor ( n1727 , n1724 , n1726 );
nor ( n1728 , n1723 , n1727 );
nand ( n1729 , n1718 , n1728 );
buf ( n1730 , n592 );
not ( n1731 , n1730 );
nor ( n1732 , n1276 , n1731 );
buf ( n1733 , n621 );
not ( n1734 , n1733 );
not ( n1735 , n1734 );
not ( n1736 , n1735 );
nor ( n1737 , n1290 , n1736 );
nor ( n1738 , n1732 , n1737 );
buf ( n1739 , n686 );
not ( n1740 , n1739 );
not ( n1741 , n1740 );
not ( n1742 , n1741 );
nor ( n1743 , n1281 , n1742 );
buf ( n1744 , n653 );
not ( n1745 , n1744 );
not ( n1746 , n1745 );
not ( n1747 , n1746 );
nor ( n1748 , n1294 , n1747 );
nor ( n1749 , n1743 , n1748 );
nand ( n1750 , n1738 , n1749 );
and ( n1751 , n1729 , n1750 );
not ( n1752 , n1281 );
buf ( n1753 , n687 );
not ( n1754 , n1753 );
not ( n1755 , n1754 );
not ( n1756 , n1755 );
not ( n1757 , n1756 );
and ( n1758 , n1752 , n1757 );
buf ( n1759 , n622 );
not ( n1760 , n1759 );
not ( n1761 , n1760 );
and ( n1762 , n1291 , n1761 );
nor ( n1763 , n1758 , n1762 );
buf ( n1764 , n593 );
not ( n1765 , n1764 );
not ( n1766 , n1765 );
not ( n1767 , n1766 );
nor ( n1768 , n1276 , n1767 );
buf ( n1769 , n654 );
not ( n1770 , n1769 );
not ( n1771 , n1770 );
not ( n1772 , n1771 );
nor ( n1773 , n1294 , n1772 );
nor ( n1774 , n1768 , n1773 );
nand ( n1775 , n1763 , n1774 );
buf ( n1776 , n631 );
not ( n1777 , n1776 );
not ( n1778 , n1777 );
nand ( n1779 , n1515 , n1778 );
buf ( n1780 , n696 );
nand ( n1781 , n1282 , n1780 );
buf ( n1782 , n663 );
not ( n1783 , n1782 );
not ( n1784 , n1783 );
nand ( n1785 , n1415 , n1784 );
nand ( n1786 , n1779 , n1781 , n1785 );
and ( n1787 , n1775 , n1786 );
buf ( n1788 , n625 );
not ( n1789 , n1788 );
not ( n1790 , n1789 );
and ( n1791 , n1587 , n1790 );
buf ( n1792 , n690 );
not ( n1793 , n1792 );
not ( n1794 , n1793 );
not ( n1795 , n1794 );
nor ( n1796 , n1520 , n1795 );
nor ( n1797 , n1791 , n1796 );
not ( n1798 , n1415 );
buf ( n1799 , n657 );
not ( n1800 , n1799 );
not ( n1801 , n1800 );
not ( n1802 , n1801 );
nor ( n1803 , n1798 , n1802 );
buf ( n1804 , n596 );
not ( n1805 , n1804 );
not ( n1806 , n1805 );
not ( n1807 , n1806 );
nor ( n1808 , n1276 , n1807 );
nor ( n1809 , n1803 , n1808 );
nand ( n1810 , n1797 , n1809 );
nand ( n1811 , n1706 , n1751 , n1787 , n1810 );
nor ( n1812 , n1681 , n1811 );
nand ( n1813 , n1514 , n1812 );
buf ( n1814 , n632 );
nand ( n1815 , n1587 , n1814 );
buf ( n1816 , n664 );
nand ( n1817 , n1415 , n1816 );
buf ( n1818 , n697 );
nand ( n1819 , n1407 , n1818 );
nand ( n1820 , n1815 , n1817 , n1819 );
not ( n1821 , n1820 );
and ( n1822 , n1813 , n1821 );
not ( n1823 , n1813 );
and ( n1824 , n1823 , n1820 );
nor ( n1825 , n1822 , n1824 );
nand ( n1826 , n1825 , n1302 );
not ( n1827 , n1826 );
buf ( n1828 , n573 );
nand ( n1829 , n1277 , n1828 );
buf ( n1830 , n634 );
not ( n1831 , n1830 );
not ( n1832 , n1831 );
nand ( n1833 , n1295 , n1832 );
buf ( n1834 , n602 );
not ( n1835 , n1834 );
not ( n1836 , n1835 );
nand ( n1837 , n1291 , n1836 );
buf ( n1838 , n667 );
nand ( n1839 , n1282 , n1838 );
nand ( n1840 , n1829 , n1833 , n1837 , n1839 );
nand ( n1841 , n1827 , n1840 );
not ( n1842 , n1841 );
or ( n1843 , n1325 , n1842 );
or ( n1844 , n1841 , n1324 );
nand ( n1845 , n1843 , n1844 );
and ( n1846 , n1304 , n1845 );
nor ( n1847 , n1303 , n1846 );
not ( n1848 , n1147 );
not ( n1849 , n1088 );
or ( n1850 , n1848 , n1849 );
not ( n1851 , n888 );
not ( n1852 , n1048 );
and ( n1853 , n1851 , n1852 );
nor ( n1854 , n1853 , n1089 );
nor ( n1855 , n1137 , n1089 );
nor ( n1856 , n1854 , n1855 );
nand ( n1857 , n1850 , n1856 );
nand ( n1858 , n1857 , n1169 );
not ( n1859 , n1858 );
not ( n1860 , n1156 );
and ( n1861 , n1859 , n1860 );
and ( n1862 , n1858 , n1156 );
nor ( n1863 , n1861 , n1862 );
not ( n1864 , n1863 );
not ( n1865 , n1864 );
buf ( n1866 , n665 );
not ( n1867 , n1866 );
nand ( n1868 , n1865 , n1867 );
not ( n1869 , n1868 );
not ( n1870 , n1156 );
nor ( n1871 , n1870 , n1858 );
xor ( n1872 , n1871 , n1182 );
not ( n1873 , n1872 );
or ( n1874 , n1869 , n1873 );
and ( n1875 , n1857 , n1169 );
not ( n1876 , n1857 );
not ( n1877 , n1169 );
and ( n1878 , n1876 , n1877 );
nor ( n1879 , n1875 , n1878 );
nand ( n1880 , n1874 , n1879 );
not ( n1881 , n1879 );
nand ( n1882 , n1881 , n1866 );
nor ( n1883 , n1864 , n1882 );
buf ( n1884 , n570 );
or ( n1885 , n1883 , n1884 );
nand ( n1886 , n1885 , n1872 );
nand ( n1887 , n1880 , n1886 );
not ( n1888 , n1864 );
not ( n1889 , n1872 );
not ( n1890 , n1889 );
or ( n1891 , n1888 , n1890 );
buf ( n1892 , n571 );
not ( n1893 , n1892 );
not ( n1894 , n1893 );
nand ( n1895 , n1879 , n1867 );
not ( n1896 , n1895 );
not ( n1897 , n1882 );
or ( n1898 , n1896 , n1897 );
nand ( n1899 , n1898 , n1865 );
not ( n1900 , n1899 );
or ( n1901 , n1894 , n1900 );
nand ( n1902 , n1901 , n1872 );
nand ( n1903 , n1891 , n1902 );
not ( n1904 , n1856 );
not ( n1905 , n1147 );
and ( n1906 , n1904 , n1905 );
and ( n1907 , n1856 , n1147 );
nor ( n1908 , n1906 , n1907 );
not ( n1909 , n1908 );
not ( n1910 , n1909 );
nand ( n1911 , n1887 , n1903 , n1910 );
not ( n1912 , n1879 );
nor ( n1913 , n1863 , n1912 );
nand ( n1914 , n1872 , n1913 );
not ( n1915 , n1099 );
nand ( n1916 , n1854 , n1915 );
nor ( n1917 , n1916 , n1115 );
nand ( n1918 , n1917 , n1123 );
xor ( n1919 , n1918 , n1136 );
not ( n1920 , n1123 );
nor ( n1921 , n1920 , n1917 );
not ( n1922 , n1921 );
not ( n1923 , n1123 );
nand ( n1924 , n1923 , n1917 );
nand ( n1925 , n1922 , n1924 );
nand ( n1926 , n1919 , n1925 );
not ( n1927 , n1926 );
not ( n1928 , n1115 );
not ( n1929 , n1928 );
not ( n1930 , n1916 );
or ( n1931 , n1929 , n1930 );
or ( n1932 , n1916 , n1928 );
nand ( n1933 , n1931 , n1932 );
and ( n1934 , n1854 , n1915 );
not ( n1935 , n1854 );
and ( n1936 , n1935 , n1099 );
nor ( n1937 , n1934 , n1936 );
nor ( n1938 , n1933 , n1937 );
buf ( n1939 , n537 );
not ( n1940 , n1939 );
not ( n1941 , n1940 );
and ( n1942 , n1938 , n1941 );
nand ( n1943 , n1914 , n1927 , n1942 );
nor ( n1944 , n1911 , n1943 );
not ( n1945 , n1944 );
or ( n1946 , n1847 , n1945 );
not ( n1947 , n1941 );
not ( n1948 , n1947 );
nand ( n1949 , n1914 , n1948 );
not ( n1950 , n1949 );
not ( n1951 , n1950 );
nor ( n1952 , n1951 , n1911 );
and ( n1953 , n1919 , n1937 );
not ( n1954 , n1919 );
and ( n1955 , n1954 , n1933 );
nor ( n1956 , n1953 , n1955 );
not ( n1957 , n1956 );
not ( n1958 , n1919 );
not ( n1959 , n1925 );
nand ( n1960 , n1958 , n1959 );
nand ( n1961 , n1960 , n1926 );
nor ( n1962 , n1957 , n1961 );
nand ( n1963 , n1952 , n1962 );
nor ( n1964 , n1961 , n1956 );
nand ( n1965 , n1952 , n1964 );
not ( n1966 , n1941 );
nor ( n1967 , n1944 , n1966 );
nand ( n1968 , n1963 , n1965 , n1967 );
not ( n1969 , n1968 );
not ( n1970 , n1925 );
not ( n1971 , n1933 );
nor ( n1972 , n1971 , n1919 );
nand ( n1973 , n1970 , n1972 );
not ( n1974 , n1973 );
not ( n1975 , n1974 );
not ( n1976 , n1952 );
or ( n1977 , n1975 , n1976 );
not ( n1978 , n1960 );
not ( n1979 , n1937 );
nor ( n1980 , n1933 , n1979 );
nand ( n1981 , n1980 , n1941 );
not ( n1982 , n1981 );
nand ( n1983 , n1914 , n1978 , n1982 , n1910 );
nand ( n1984 , n1977 , n1983 );
nand ( n1985 , n1914 , n1978 , n1942 );
nor ( n1986 , n1911 , n1985 );
nor ( n1987 , n1984 , n1986 );
nand ( n1988 , n1969 , n1987 );
not ( n1989 , n1947 );
nand ( n1990 , n1988 , n1989 );
and ( n1991 , n1990 , n1828 );
not ( n1992 , n1302 );
not ( n1993 , n1186 );
not ( n1994 , n1196 );
and ( n1995 , n1993 , n1994 );
and ( n1996 , n1186 , n1196 );
nor ( n1997 , n1995 , n1996 );
and ( n1998 , n1196 , n1211 );
not ( n1999 , n1196 );
and ( n2000 , n1999 , n1210 );
nor ( n2001 , n1998 , n2000 );
nand ( n2002 , n1997 , n2001 );
or ( n2003 , n2002 , n966 );
buf ( n2004 , n536 );
nand ( n2005 , n2002 , n2004 );
nand ( n2006 , n2003 , n2005 );
not ( n2007 , n2006 );
nand ( n2008 , n1992 , n2007 );
not ( n2009 , n2008 );
not ( n2010 , n2009 );
not ( n2011 , n2002 );
not ( n2012 , n965 );
and ( n2013 , n2011 , n2012 );
buf ( n2014 , n535 );
and ( n2015 , n2002 , n2014 );
nor ( n2016 , n2013 , n2015 );
not ( n2017 , n2016 );
or ( n2018 , n2017 , n1840 );
nand ( n2019 , n1840 , n2017 );
nand ( n2020 , n2018 , n2019 );
nor ( n2021 , n2020 , n1302 );
not ( n2022 , n2021 );
nand ( n2023 , n2020 , n1302 );
nand ( n2024 , n2022 , n2023 );
not ( n2025 , n2024 );
or ( n2026 , n2010 , n2025 );
or ( n2027 , n2024 , n2009 );
nand ( n2028 , n2026 , n2027 );
not ( n2029 , n1965 );
nand ( n2030 , n2028 , n2029 );
not ( n2031 , n1963 );
not ( n2032 , n2017 );
not ( n2033 , n1840 );
not ( n2034 , n2033 );
or ( n2035 , n2032 , n2034 );
not ( n2036 , n2017 );
nand ( n2037 , n1840 , n2036 );
nand ( n2038 , n2035 , n2037 );
not ( n2039 , n1302 );
not ( n2040 , n2006 );
nor ( n2041 , n2039 , n2040 );
xor ( n2042 , n2038 , n2041 );
nand ( n2043 , n2031 , n2042 );
nand ( n2044 , n1984 , n2017 );
not ( n2045 , n1986 );
not ( n2046 , n2045 );
not ( n2047 , n2017 );
not ( n2048 , n2047 );
not ( n2049 , n2006 );
or ( n2050 , n2048 , n2049 );
or ( n2051 , n2006 , n2047 );
nand ( n2052 , n2050 , n2051 );
nand ( n2053 , n2046 , n2052 );
nand ( n2054 , n2030 , n2043 , n2044 , n2053 );
nor ( n2055 , n1991 , n2054 );
nand ( n2056 , n1946 , n2055 );
buf ( n2057 , n2056 );
buf ( n2058 , n2057 );
buf ( n2059 , n531 );
not ( n2060 , n2059 );
not ( n2061 , n2060 );
buf ( n2062 , n2061 );
buf ( n2063 , n2062 );
buf ( n2064 , n698 );
and ( n2065 , n1217 , n1840 );
not ( n2066 , n1217 );
nand ( n2067 , n1498 , n1277 );
or ( n2068 , n1498 , n1277 );
and ( n2069 , n2067 , n2068 );
not ( n2070 , n1324 );
nor ( n2071 , n2070 , n1841 );
xor ( n2072 , n2069 , n2071 );
and ( n2073 , n2066 , n2072 );
nor ( n2074 , n2065 , n2073 );
or ( n2075 , n2074 , n1945 );
and ( n2076 , n1990 , n1305 );
not ( n2077 , n2045 );
not ( n2078 , n2002 );
not ( n2079 , n953 );
not ( n2080 , n2079 );
and ( n2081 , n2078 , n2080 );
buf ( n2082 , n534 );
and ( n2083 , n2002 , n2082 );
nor ( n2084 , n2081 , n2083 );
not ( n2085 , n2084 );
not ( n2086 , n2085 );
not ( n2087 , n2047 );
nor ( n2088 , n2087 , n2006 );
not ( n2089 , n2088 );
or ( n2090 , n2086 , n2089 );
or ( n2091 , n2088 , n2085 );
nand ( n2092 , n2090 , n2091 );
not ( n2093 , n2092 );
not ( n2094 , n2093 );
and ( n2095 , n2077 , n2094 );
not ( n2096 , n2085 );
not ( n2097 , n2096 );
not ( n2098 , n1324 );
not ( n2099 , n2098 );
or ( n2100 , n2097 , n2099 );
nand ( n2101 , n1324 , n2085 );
nand ( n2102 , n2100 , n2101 );
not ( n2103 , n1840 );
nor ( n2104 , n2103 , n2017 );
nor ( n2105 , n2102 , n2104 );
not ( n2106 , n2105 );
nand ( n2107 , n2102 , n2104 );
nand ( n2108 , n2106 , n2107 );
not ( n2109 , n2108 );
or ( n2110 , n2021 , n2008 );
nand ( n2111 , n2110 , n2023 );
not ( n2112 , n2111 );
or ( n2113 , n2109 , n2112 );
or ( n2114 , n2108 , n2111 );
nand ( n2115 , n2113 , n2114 );
and ( n2116 , n2115 , n2029 );
nor ( n2117 , n2095 , n2116 );
not ( n2118 , n1984 );
not ( n2119 , n2118 );
not ( n2120 , n2085 );
not ( n2121 , n2120 );
and ( n2122 , n2119 , n2121 );
nand ( n2123 , n2038 , n2041 );
not ( n2124 , n2123 );
not ( n2125 , n2124 );
not ( n2126 , n2085 );
not ( n2127 , n1324 );
not ( n2128 , n2127 );
or ( n2129 , n2126 , n2128 );
not ( n2130 , n2085 );
nand ( n2131 , n2130 , n1324 );
nand ( n2132 , n2129 , n2131 );
not ( n2133 , n2132 );
not ( n2134 , n1840 );
nor ( n2135 , n2134 , n2036 );
not ( n2136 , n2135 );
nand ( n2137 , n2133 , n2136 );
nand ( n2138 , n2132 , n2135 );
nand ( n2139 , n2137 , n2138 );
not ( n2140 , n2139 );
or ( n2141 , n2125 , n2140 );
or ( n2142 , n2139 , n2124 );
nand ( n2143 , n2141 , n2142 );
and ( n2144 , n2143 , n2031 );
nor ( n2145 , n2122 , n2144 );
nand ( n2146 , n2117 , n2145 );
nor ( n2147 , n2076 , n2146 );
nand ( n2148 , n2075 , n2147 );
buf ( n2149 , n2148 );
buf ( n2150 , n2149 );
not ( n2151 , n2060 );
buf ( n2152 , n2151 );
buf ( n2153 , n2152 );
buf ( n2154 , n698 );
not ( n2155 , n1216 );
and ( n2156 , n2155 , n1324 );
not ( n2157 , n2155 );
nand ( n2158 , n2071 , n2069 );
not ( n2159 , n1372 );
not ( n2160 , n2067 );
or ( n2161 , n2159 , n2160 );
or ( n2162 , n2067 , n1372 );
nand ( n2163 , n2161 , n2162 );
not ( n2164 , n2163 );
and ( n2165 , n2158 , n2164 );
not ( n2166 , n2158 );
and ( n2167 , n2166 , n2163 );
nor ( n2168 , n2165 , n2167 );
and ( n2169 , n2157 , n2168 );
nor ( n2170 , n2156 , n2169 );
or ( n2171 , n2170 , n1945 );
nor ( n2172 , n2021 , n2105 );
nand ( n2173 , n2023 , n2008 );
nand ( n2174 , n2172 , n2173 );
not ( n2175 , n2174 );
not ( n2176 , n2175 );
nand ( n2177 , n2176 , n2107 );
not ( n2178 , n1277 );
not ( n2179 , n1498 );
not ( n2180 , n2179 );
or ( n2181 , n2178 , n2180 );
not ( n2182 , n1277 );
nand ( n2183 , n1498 , n2182 );
nand ( n2184 , n2181 , n2183 );
not ( n2185 , n930 );
not ( n2186 , n2002 );
not ( n2187 , n2186 );
or ( n2188 , n2185 , n2187 );
buf ( n2189 , n533 );
nand ( n2190 , n2002 , n2189 );
nand ( n2191 , n2188 , n2190 );
not ( n2192 , n2191 );
and ( n2193 , n2184 , n2192 );
not ( n2194 , n2184 );
and ( n2195 , n2194 , n2191 );
nor ( n2196 , n2193 , n2195 );
and ( n2197 , n1324 , n2096 );
nor ( n2198 , n2196 , n2197 );
not ( n2199 , n2198 );
nand ( n2200 , n2196 , n2197 );
nand ( n2201 , n2199 , n2200 );
xnor ( n2202 , n2177 , n2201 );
and ( n2203 , n2202 , n2029 );
and ( n2204 , n1984 , n2191 );
nor ( n2205 , n2203 , n2204 );
nand ( n2206 , n2137 , n2124 );
not ( n2207 , n2206 );
not ( n2208 , n2207 );
nand ( n2209 , n2208 , n2138 );
not ( n2210 , n2209 );
xor ( n2211 , n1277 , n1498 );
xor ( n2212 , n2211 , n2191 );
and ( n2213 , n1324 , n2085 );
or ( n2214 , n2212 , n2213 );
nand ( n2215 , n2212 , n2213 );
nand ( n2216 , n2214 , n2215 );
not ( n2217 , n2216 );
or ( n2218 , n2210 , n2217 );
or ( n2219 , n2216 , n2209 );
nand ( n2220 , n2218 , n2219 );
and ( n2221 , n2220 , n2031 );
not ( n2222 , n2046 );
not ( n2223 , n2191 );
not ( n2224 , n2088 );
nor ( n2225 , n2224 , n2085 );
not ( n2226 , n2225 );
or ( n2227 , n2223 , n2226 );
or ( n2228 , n2225 , n2191 );
nand ( n2229 , n2227 , n2228 );
not ( n2230 , n2229 );
or ( n2231 , n2222 , n2230 );
not ( n2232 , n1491 );
nor ( n2233 , n2232 , n1989 );
not ( n2234 , n2233 );
nand ( n2235 , n2231 , n2234 );
nor ( n2236 , n2221 , n2235 );
not ( n2237 , n1988 );
nand ( n2238 , n2237 , n2232 );
and ( n2239 , n2205 , n2236 , n2238 );
nand ( n2240 , n2171 , n2239 );
buf ( n2241 , n2240 );
buf ( n2242 , n2241 );
not ( n2243 , n2060 );
buf ( n2244 , n2243 );
buf ( n2245 , n2244 );
buf ( n2246 , n698 );
not ( n2247 , n1216 );
nand ( n2248 , n1498 , n1277 );
not ( n2249 , n1372 );
or ( n2250 , n2248 , n2249 );
not ( n2251 , n1346 );
and ( n2252 , n2250 , n2251 );
not ( n2253 , n2250 );
and ( n2254 , n2253 , n1346 );
nor ( n2255 , n2252 , n2254 );
not ( n2256 , n2255 );
and ( n2257 , n1840 , n1324 );
nand ( n2258 , n2163 , n2069 , n2257 );
not ( n2259 , n2258 );
not ( n2260 , n1827 );
not ( n2261 , n2260 );
nand ( n2262 , n2259 , n2261 );
not ( n2263 , n2262 );
or ( n2264 , n2256 , n2263 );
or ( n2265 , n2262 , n2255 );
nand ( n2266 , n2264 , n2265 );
not ( n2267 , n2266 );
or ( n2268 , n2247 , n2267 );
nand ( n2269 , n2069 , n1217 );
nand ( n2270 , n2268 , n2269 );
not ( n2271 , n2270 );
or ( n2272 , n2271 , n1945 );
not ( n2273 , n2199 );
not ( n2274 , n2175 );
or ( n2275 , n2273 , n2274 );
not ( n2276 , n2107 );
and ( n2277 , n2199 , n2276 );
not ( n2278 , n2200 );
nor ( n2279 , n2277 , n2278 );
nand ( n2280 , n2275 , n2279 );
not ( n2281 , n1372 );
not ( n2282 , n2002 );
not ( n2283 , n942 );
and ( n2284 , n2282 , n2283 );
buf ( n2285 , n532 );
and ( n2286 , n2002 , n2285 );
nor ( n2287 , n2284 , n2286 );
not ( n2288 , n2287 );
not ( n2289 , n2288 );
or ( n2290 , n2281 , n2289 );
or ( n2291 , n2288 , n1372 );
nand ( n2292 , n2290 , n2291 );
not ( n2293 , n2182 );
not ( n2294 , n1498 );
not ( n2295 , n2294 );
or ( n2296 , n2293 , n2295 );
nand ( n2297 , n2296 , n2192 );
not ( n2298 , n2294 );
nand ( n2299 , n2298 , n1277 );
nand ( n2300 , n2297 , n2299 );
nor ( n2301 , n2292 , n2300 );
not ( n2302 , n2301 );
nand ( n2303 , n2300 , n2292 );
nand ( n2304 , n2302 , n2303 );
xnor ( n2305 , n2280 , n2304 );
nand ( n2306 , n2305 , n2029 );
xor ( n2307 , n1277 , n1498 );
and ( n2308 , n2307 , n2191 );
and ( n2309 , n1277 , n1498 );
or ( n2310 , n2308 , n2309 );
not ( n2311 , n2310 );
not ( n2312 , n1372 );
not ( n2313 , n2288 );
not ( n2314 , n2313 );
or ( n2315 , n2312 , n2314 );
not ( n2316 , n1372 );
nand ( n2317 , n2316 , n2288 );
nand ( n2318 , n2315 , n2317 );
not ( n2319 , n2318 );
nand ( n2320 , n2311 , n2319 );
and ( n2321 , n2310 , n2318 );
not ( n2322 , n2321 );
nand ( n2323 , n2320 , n2322 );
not ( n2324 , n2323 );
nand ( n2325 , n2207 , n2214 );
not ( n2326 , n2138 );
nand ( n2327 , n2214 , n2326 );
nand ( n2328 , n2325 , n2327 , n2215 );
not ( n2329 , n2328 );
or ( n2330 , n2324 , n2329 );
or ( n2331 , n2328 , n2323 );
nand ( n2332 , n2330 , n2331 );
nand ( n2333 , n2332 , n2031 );
not ( n2334 , n2288 );
not ( n2335 , n2334 );
and ( n2336 , n1984 , n2335 );
nor ( n2337 , n2191 , n2085 );
and ( n2338 , n2088 , n2337 );
not ( n2339 , n2334 );
not ( n2340 , n2339 );
and ( n2341 , n2338 , n2340 );
not ( n2342 , n2338 );
and ( n2343 , n2342 , n2339 );
nor ( n2344 , n2341 , n2343 );
not ( n2345 , n2344 );
not ( n2346 , n2046 );
or ( n2347 , n2345 , n2346 );
nand ( n2348 , n1367 , n1947 );
nand ( n2349 , n2347 , n2348 );
nor ( n2350 , n2336 , n2349 );
nand ( n2351 , n2306 , n2333 , n2350 );
not ( n2352 , n1367 );
and ( n2353 , n2352 , n1491 );
and ( n2354 , n2232 , n1367 );
nor ( n2355 , n2353 , n2354 );
nor ( n2356 , n1988 , n2355 );
nor ( n2357 , n2351 , n2356 );
nand ( n2358 , n2272 , n2357 );
buf ( n2359 , n2358 );
buf ( n2360 , n2359 );
endmodule
