module top( n19 , n24 , n29 , n32 , n36 , n49 , n52 , n58 , n59 ,
n60 , n69 , n73 , n76 , n96 , n97 , n100 , n108 , n117 , n123 ,
n143 , n149 , n151 , n152 , n158 , n167 , n189 , n194 , n196 , n197 ,
n198 , n206 , n209 , n210 , n217 , n218 , n222 , n224 , n226 , n233 ,
n242 , n245 , n248 , n258 );
    input n19 , n24 , n32 , n36 , n49 , n52 , n58 , n59 , n60 ,
n69 , n73 , n96 , n97 , n100 , n108 , n117 , n123 , n143 , n149 ,
n151 , n158 , n167 , n189 , n196 , n197 , n198 , n206 , n209 , n210 ,
n217 , n218 , n222 , n226 , n233 , n242 , n258 ;
    output n29 , n76 , n152 , n194 , n224 , n245 , n248 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 ,
n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 ,
n20 , n21 , n22 , n23 , n25 , n26 , n27 , n28 , n30 , n31 ,
n33 , n34 , n35 , n37 , n38 , n39 , n40 , n41 , n42 , n43 ,
n44 , n45 , n46 , n47 , n48 , n50 , n51 , n53 , n54 , n55 ,
n56 , n57 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 ,
n70 , n71 , n72 , n74 , n75 , n77 , n78 , n79 , n80 , n81 ,
n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 ,
n92 , n93 , n94 , n95 , n98 , n99 , n101 , n102 , n103 , n104 ,
n105 , n106 , n107 , n109 , n110 , n111 , n112 , n113 , n114 , n115 ,
n116 , n118 , n119 , n120 , n121 , n122 , n124 , n125 , n126 , n127 ,
n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 ,
n138 , n139 , n140 , n141 , n142 , n144 , n145 , n146 , n147 , n148 ,
n150 , n153 , n154 , n155 , n156 , n157 , n159 , n160 , n161 , n162 ,
n163 , n164 , n165 , n166 , n168 , n169 , n170 , n171 , n172 , n173 ,
n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 ,
n184 , n185 , n186 , n187 , n188 , n190 , n191 , n192 , n193 , n195 ,
n199 , n200 , n201 , n202 , n203 , n204 , n205 , n207 , n208 , n211 ,
n212 , n213 , n214 , n215 , n216 , n219 , n220 , n221 , n223 , n225 ,
n227 , n228 , n229 , n230 , n231 , n232 , n234 , n235 , n236 , n237 ,
n238 , n239 , n240 , n241 , n243 , n244 , n246 , n247 , n249 , n250 ,
n251 , n252 , n253 , n254 , n255 , n256 , n257 , n259 , n260 , n261 ,
n262 ;
    xnor g0 ( n95 , n29 , n40 );
    not g1 ( n43 , n218 );
    nor g2 ( n141 , n87 , n5 );
    and g3 ( n216 , n123 , n179 );
    or g4 ( n180 , n253 , n88 );
    xor g5 ( n2 , n245 , n190 );
    not g6 ( n88 , n213 );
    and g7 ( n191 , n185 , n114 );
    or g8 ( n199 , n250 , n157 );
    and g9 ( n129 , n109 , n214 );
    and g10 ( n236 , n21 , n10 );
    not g11 ( n40 , n184 );
    and g12 ( n168 , n117 , n137 );
    buf g13 ( n27 , n117 );
    nor g14 ( n9 , n220 , n42 );
    or g15 ( n7 , n129 , n34 );
    not g16 ( n41 , n168 );
    not g17 ( n257 , n210 );
    not g18 ( n70 , n197 );
    and g19 ( n156 , n150 , n141 );
    or g20 ( n173 , n68 , n11 );
    xnor g21 ( n223 , n29 , n35 );
    or g22 ( n219 , n120 , n131 );
    and g23 ( n262 , n70 , n55 );
    not g24 ( n28 , n149 );
    or g25 ( n122 , n243 , n238 );
    and g26 ( n120 , n69 , n29 );
    xor g27 ( n94 , n245 , n31 );
    not g28 ( n137 , n233 );
    not g29 ( n237 , n222 );
    and g30 ( n75 , n59 , n204 );
    or g31 ( n205 , n99 , n126 );
    xor g32 ( n215 , n245 , n154 );
    or g33 ( n155 , n70 , n88 );
    and g34 ( n99 , n12 , n33 );
    nor g35 ( n239 , n145 , n234 );
    or g36 ( n111 , n28 , n49 );
    and g37 ( n104 , n163 , n208 );
    or g38 ( n224 , n85 , n56 );
    not g39 ( n193 , n190 );
    or g40 ( n175 , n192 , n20 );
    or g41 ( n0 , n223 , n215 );
    or g42 ( n47 , n204 , n72 );
    not g43 ( n102 , n209 );
    and g44 ( n170 , n149 , n202 );
    or g45 ( n203 , n3 , n46 );
    nor g46 ( n183 , n166 , n223 );
    nor g47 ( n55 , n93 , n68 );
    nor g48 ( n246 , n102 , n225 );
    nor g49 ( n89 , n195 , n95 );
    and g50 ( n184 , n100 , n64 );
    not g51 ( n166 , n123 );
    not g52 ( n110 , n79 );
    not g53 ( n153 , n117 );
    and g54 ( n34 , n44 , n105 );
    not g55 ( n234 , n18 );
    buf g56 ( n61 , n65 );
    nor g57 ( n82 , n227 , n165 );
    not g58 ( n221 , n188 );
    or g59 ( n130 , n75 , n13 );
    and g60 ( n18 , n26 , n106 );
    or g61 ( n152 , n6 , n207 );
    and g62 ( n65 , n191 , n216 );
    xor g63 ( n144 , n245 , n241 );
    and g64 ( n12 , n47 , n155 );
    nor g65 ( n243 , n164 , n212 );
    or g66 ( n150 , n128 , n69 );
    or g67 ( n211 , n122 , n30 );
    or g68 ( n86 , n188 , n110 );
    or g69 ( n6 , n99 , n112 );
    and g70 ( n78 , n100 , n25 );
    or g71 ( n83 , n128 , n136 );
    not g72 ( n192 , n19 );
    or g73 ( n42 , n225 , n228 );
    and g74 ( n79 , n186 , n71 );
    nor g75 ( n53 , n61 , n86 );
    or g76 ( n62 , n251 , n135 );
    or g77 ( n164 , n50 , n32 );
    and g78 ( n71 , n149 , n54 );
    or g79 ( n163 , n64 , n72 );
    not g80 ( n169 , n49 );
    and g81 ( n3 , n258 , n43 );
    nor g82 ( n76 , n17 , n63 );
    or g83 ( n101 , n43 , n72 );
    and g84 ( n136 , n198 , n194 );
    xor g85 ( n4 , n245 , n178 );
    not g86 ( n20 , n194 );
    and g87 ( n67 , n77 , n180 );
    not g88 ( n204 , n151 );
    or g89 ( n85 , n99 , n188 );
    not g90 ( n35 , n46 );
    not g91 ( n29 , n156 );
    or g92 ( n248 , n171 , n205 );
    or g93 ( n148 , n188 , n236 );
    not g94 ( n107 , n170 );
    and g95 ( n31 , n237 , n51 );
    not g96 ( n252 , n194 );
    nor g97 ( n146 , n230 , n16 );
    nor g98 ( n51 , n28 , n200 );
    or g99 ( n1 , n257 , n45 );
    or g100 ( n244 , n80 , n146 );
    or g101 ( n124 , n202 , n45 );
    not g102 ( n250 , n158 );
    xor g103 ( n231 , n245 , n34 );
    not g104 ( n213 , n15 );
    not g105 ( n45 , n38 );
    nor g106 ( n17 , n148 , n62 );
    not g107 ( n38 , n156 );
    or g108 ( n121 , n166 , n226 );
    and g109 ( n15 , n193 , n82 );
    or g110 ( n139 , n237 , n88 );
    or g111 ( n177 , n260 , n244 );
    not g112 ( n253 , n52 );
    nor g113 ( n214 , n50 , n39 );
    not g114 ( n93 , n59 );
    and g115 ( n112 , n159 , n239 );
    not g116 ( n109 , n189 );
    and g117 ( n178 , n250 , n127 );
    and g118 ( n21 , n1 , n199 );
    or g119 ( n77 , n91 , n72 );
    not g120 ( n57 , n75 );
    and g121 ( n13 , n209 , n91 );
    xnor g122 ( n235 , n29 , n150 );
    or g123 ( n165 , n22 , n7 );
    not g124 ( n232 , n160 );
    xnor g125 ( n200 , n29 , n107 );
    nor g126 ( n174 , n236 , n240 );
    nor g127 ( n159 , n188 , n236 );
    not g128 ( n14 , n60 );
    not g129 ( n128 , n73 );
    not g130 ( n181 , n242 );
    not g131 ( n72 , n38 );
    or g132 ( n81 , n99 , n27 );
    not g133 ( n254 , n206 );
    not g134 ( n125 , n96 );
    xor g135 ( n256 , n245 , n129 );
    or g136 ( n5 , n203 , n116 );
    and g137 ( n132 , n209 , n8 );
    and g138 ( n154 , n254 , n183 );
    or g139 ( n176 , n128 , n198 );
    nor g140 ( n80 , n172 , n74 );
    or g141 ( n16 , n95 , n144 );
    not g142 ( n119 , n217 );
    or g143 ( n185 , n48 , n45 );
    not g144 ( n44 , n196 );
    or g145 ( n227 , n103 , n187 );
    or g146 ( n140 , n109 , n157 );
    xor g147 ( n228 , n245 , n255 );
    or g148 ( n54 , n169 , n20 );
    or g149 ( n201 , n177 , n211 );
    and g150 ( n145 , n104 , n78 );
    or g151 ( n74 , n142 , n4 );
    or g152 ( n8 , n125 , n20 );
    or g153 ( n207 , n126 , n53 );
    and g154 ( n10 , n217 , n175 );
    not g155 ( n229 , n167 );
    not g156 ( n133 , n143 );
    or g157 ( n212 , n39 , n256 );
    or g158 ( n230 , n195 , n167 );
    or g159 ( n25 , n229 , n20 );
    xnor g160 ( n98 , n29 , n41 );
    or g161 ( n171 , n188 , n145 );
    not g162 ( n247 , n65 );
    nor g163 ( n238 , n121 , n0 );
    nor g164 ( n105 , n153 , n98 );
    or g165 ( n113 , n261 , n252 );
    or g166 ( n103 , n255 , n178 );
    or g167 ( n249 , n160 , n184 );
    and g168 ( n106 , n258 , n113 );
    or g169 ( n179 , n134 , n252 );
    or g170 ( n116 , n170 , n168 );
    xnor g171 ( n225 , n29 , n138 );
    xnor g172 ( n142 , n29 , n232 );
    nor g173 ( n63 , n219 , n83 );
    not g174 ( n134 , n226 );
    not g175 ( n259 , n3 );
    not g176 ( n50 , n258 );
    or g177 ( n30 , n66 , n92 );
    or g178 ( n147 , n18 , n79 );
    not g179 ( n157 , n213 );
    xor g180 ( n11 , n245 , n262 );
    not g181 ( n64 , n24 );
    or g182 ( n37 , n93 , n143 );
    or g183 ( n240 , n145 , n247 );
    xnor g184 ( n39 , n29 , n259 );
    not g185 ( n245 , n15 );
    nor g186 ( n115 , n37 , n173 );
    or g187 ( n87 , n130 , n249 );
    not g188 ( n261 , n32 );
    or g189 ( n22 , n241 , n154 );
    or g190 ( n172 , n119 , n19 );
    and g191 ( n26 , n101 , n140 );
    not g192 ( n48 , n97 );
    or g193 ( n194 , n84 , n201 );
    and g194 ( n33 , n59 , n90 );
    and g195 ( n186 , n124 , n139 );
    or g196 ( n187 , n262 , n31 );
    and g197 ( n188 , n67 , n132 );
    not g198 ( n195 , n100 );
    and g199 ( n160 , n217 , n257 );
    or g200 ( n162 , n200 , n94 );
    or g201 ( n114 , n254 , n157 );
    nor g202 ( n182 , n128 , n235 );
    or g203 ( n220 , n102 , n96 );
    nor g204 ( n92 , n118 , n161 );
    or g205 ( n90 , n133 , n252 );
    nor g206 ( n66 , n111 , n162 );
    not g207 ( n91 , n108 );
    nor g208 ( n84 , n176 , n23 );
    or g209 ( n56 , n174 , n112 );
    and g210 ( n241 , n14 , n89 );
    not g211 ( n202 , n58 );
    and g212 ( n190 , n181 , n182 );
    and g213 ( n46 , n123 , n48 );
    or g214 ( n260 , n115 , n9 );
    or g215 ( n208 , n14 , n88 );
    or g216 ( n251 , n145 , n65 );
    or g217 ( n118 , n153 , n36 );
    and g218 ( n255 , n253 , n246 );
    or g219 ( n135 , n147 , n81 );
    xnor g220 ( n68 , n29 , n57 );
    or g221 ( n161 , n98 , n231 );
    not g222 ( n138 , n13 );
    or g223 ( n23 , n235 , n2 );
    and g224 ( n131 , n242 , n245 );
    and g225 ( n126 , n221 , n236 );
    nor g226 ( n127 , n119 , n142 );
endmodule
