module top( n7 , n9 , n12 , n18 , n19 , n33 , n38 , n39 , n56 ,
n60 , n61 , n64 , n66 , n67 , n75 , n77 , n83 , n84 , n92 ,
n101 , n107 , n112 , n117 , n119 , n123 , n128 , n129 , n130 , n132 ,
n157 , n158 , n165 , n168 , n173 , n179 , n186 , n187 , n190 , n193 ,
n211 , n222 , n228 , n235 , n236 , n238 , n239 , n245 , n249 , n257 ,
n259 , n261 , n262 , n264 , n270 , n288 , n297 , n307 , n315 , n319 ,
n320 , n321 , n326 , n335 , n337 , n342 , n357 , n361 , n370 , n371 ,
n375 , n377 , n378 , n379 , n380 , n381 , n384 , n386 , n387 , n389 ,
n403 , n413 , n417 , n448 , n454 , n456 , n457 , n476 , n482 , n487 ,
n488 , n495 , n504 , n516 , n520 , n530 , n541 , n542 , n544 , n547 ,
n560 , n564 , n565 , n566 , n567 , n574 , n579 , n591 , n596 , n600 ,
n601 , n606 , n611 , n617 , n623 , n627 , n635 , n636 , n643 , n649 ,
n661 , n668 , n673 , n676 , n697 , n708 , n714 , n715 , n721 , n722 ,
n754 , n758 , n760 , n765 , n776 , n779 , n786 , n793 , n801 , n807 ,
n813 , n824 , n830 , n840 , n841 , n845 , n849 , n850 , n860 , n878 ,
n882 , n887 , n889 , n894 , n912 , n917 , n918 , n937 , n944 , n946 ,
n951 , n955 , n961 , n962 , n964 , n966 , n967 , n971 , n974 , n984 ,
n999 , n1016 , n1027 , n1033 , n1039 , n1043 , n1044 , n1047 , n1050 , n1058 ,
n1065 , n1087 , n1088 , n1095 , n1096 , n1097 , n1100 , n1110 , n1119 , n1125 ,
n1135 , n1140 , n1150 , n1163 , n1172 , n1175 , n1177 , n1180 , n1181 , n1182 ,
n1186 , n1205 , n1207 , n1219 , n1224 , n1227 , n1233 , n1238 , n1269 , n1270 ,
n1279 , n1281 , n1288 , n1297 , n1299 , n1314 , n1322 , n1338 , n1346 , n1353 ,
n1355 , n1357 , n1361 , n1362 , n1363 , n1366 , n1370 , n1377 , n1378 , n1390 ,
n1391 , n1396 , n1402 , n1406 , n1408 , n1409 , n1414 , n1425 , n1426 , n1427 ,
n1435 , n1436 , n1454 , n1462 , n1463 , n1464 , n1471 , n1485 , n1491 , n1495 ,
n1498 , n1503 , n1510 , n1511 , n1515 , n1518 , n1519 , n1534 , n1540 , n1543 ,
n1553 , n1568 , n1575 , n1584 , n1587 , n1598 , n1613 , n1631 , n1632 , n1633 ,
n1649 , n1654 , n1655 , n1657 , n1660 , n1663 , n1674 , n1675 , n1676 , n1682 ,
n1697 , n1698 , n1700 , n1707 , n1708 , n1710 , n1721 , n1729 , n1733 , n1740 ,
n1743 , n1753 , n1755 , n1756 , n1761 , n1768 , n1780 , n1784 , n1788 , n1790 ,
n1793 , n1794 );
    input n7 , n9 , n12 , n19 , n33 , n38 , n39 , n60 , n64 ,
n77 , n84 , n92 , n119 , n128 , n132 , n157 , n179 , n186 , n187 ,
n190 , n228 , n236 , n238 , n239 , n257 , n261 , n270 , n288 , n297 ,
n307 , n319 , n321 , n326 , n335 , n342 , n371 , n377 , n378 , n380 ,
n384 , n386 , n387 , n389 , n403 , n448 , n457 , n482 , n488 , n495 ,
n504 , n516 , n520 , n530 , n541 , n544 , n560 , n564 , n565 , n566 ,
n579 , n591 , n600 , n601 , n606 , n617 , n627 , n636 , n643 , n668 ,
n676 , n697 , n708 , n714 , n715 , n721 , n754 , n758 , n760 , n779 ,
n801 , n807 , n813 , n830 , n841 , n850 , n887 , n894 , n912 , n917 ,
n918 , n937 , n946 , n955 , n961 , n962 , n966 , n971 , n984 , n999 ,
n1016 , n1033 , n1039 , n1043 , n1058 , n1088 , n1095 , n1097 , n1100 , n1119 ,
n1125 , n1135 , n1150 , n1172 , n1175 , n1177 , n1180 , n1181 , n1182 , n1205 ,
n1207 , n1219 , n1227 , n1238 , n1279 , n1281 , n1288 , n1299 , n1338 , n1353 ,
n1357 , n1361 , n1362 , n1363 , n1366 , n1391 , n1396 , n1402 , n1406 , n1408 ,
n1426 , n1427 , n1435 , n1436 , n1454 , n1463 , n1471 , n1485 , n1498 , n1503 ,
n1515 , n1518 , n1519 , n1534 , n1540 , n1553 , n1568 , n1575 , n1598 , n1613 ,
n1632 , n1633 , n1649 , n1655 , n1660 , n1663 , n1674 , n1675 , n1700 , n1707 ,
n1729 , n1740 , n1743 , n1753 , n1755 , n1756 , n1768 , n1788 , n1790 ;
    output n18 , n56 , n61 , n66 , n67 , n75 , n83 , n101 , n107 ,
n112 , n117 , n123 , n129 , n130 , n158 , n165 , n168 , n173 , n193 ,
n211 , n222 , n235 , n245 , n249 , n259 , n262 , n264 , n315 , n320 ,
n337 , n357 , n361 , n370 , n375 , n379 , n381 , n413 , n417 , n454 ,
n456 , n476 , n487 , n542 , n547 , n567 , n574 , n596 , n611 , n623 ,
n635 , n649 , n661 , n673 , n722 , n765 , n776 , n786 , n793 , n824 ,
n840 , n845 , n849 , n860 , n878 , n882 , n889 , n944 , n951 , n964 ,
n967 , n974 , n1027 , n1044 , n1047 , n1050 , n1065 , n1087 , n1096 , n1110 ,
n1140 , n1163 , n1186 , n1224 , n1233 , n1269 , n1270 , n1297 , n1314 , n1322 ,
n1346 , n1355 , n1370 , n1377 , n1378 , n1390 , n1409 , n1414 , n1425 , n1462 ,
n1464 , n1491 , n1495 , n1510 , n1511 , n1543 , n1584 , n1587 , n1631 , n1654 ,
n1657 , n1676 , n1682 , n1697 , n1698 , n1708 , n1710 , n1721 , n1733 , n1761 ,
n1780 , n1784 , n1793 , n1794 ;
    wire n0 , n1 , n2 , n3 , n4 , n5 , n6 , n8 , n10 ,
n11 , n13 , n14 , n15 , n16 , n17 , n20 , n21 , n22 , n23 ,
n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n34 ,
n35 , n36 , n37 , n40 , n41 , n42 , n43 , n44 , n45 , n46 ,
n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n57 ,
n58 , n59 , n62 , n63 , n65 , n68 , n69 , n70 , n71 , n72 ,
n73 , n74 , n76 , n78 , n79 , n80 , n81 , n82 , n85 , n86 ,
n87 , n88 , n89 , n90 , n91 , n93 , n94 , n95 , n96 , n97 ,
n98 , n99 , n100 , n102 , n103 , n104 , n105 , n106 , n108 , n109 ,
n110 , n111 , n113 , n114 , n115 , n116 , n118 , n120 , n121 , n122 ,
n124 , n125 , n126 , n127 , n131 , n133 , n134 , n135 , n136 , n137 ,
n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 ,
n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n159 ,
n160 , n161 , n162 , n163 , n164 , n166 , n167 , n169 , n170 , n171 ,
n172 , n174 , n175 , n176 , n177 , n178 , n180 , n181 , n182 , n183 ,
n184 , n185 , n188 , n189 , n191 , n192 , n194 , n195 , n196 , n197 ,
n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 ,
n208 , n209 , n210 , n212 , n213 , n214 , n215 , n216 , n217 , n218 ,
n219 , n220 , n221 , n223 , n224 , n225 , n226 , n227 , n229 , n230 ,
n231 , n232 , n233 , n234 , n237 , n240 , n241 , n242 , n243 , n244 ,
n246 , n247 , n248 , n250 , n251 , n252 , n253 , n254 , n255 , n256 ,
n258 , n260 , n263 , n265 , n266 , n267 , n268 , n269 , n271 , n272 ,
n273 , n274 , n275 , n276 , n277 , n278 , n279 , n280 , n281 , n282 ,
n283 , n284 , n285 , n286 , n287 , n289 , n290 , n291 , n292 , n293 ,
n294 , n295 , n296 , n298 , n299 , n300 , n301 , n302 , n303 , n304 ,
n305 , n306 , n308 , n309 , n310 , n311 , n312 , n313 , n314 , n316 ,
n317 , n318 , n322 , n323 , n324 , n325 , n327 , n328 , n329 , n330 ,
n331 , n332 , n333 , n334 , n336 , n338 , n339 , n340 , n341 , n343 ,
n344 , n345 , n346 , n347 , n348 , n349 , n350 , n351 , n352 , n353 ,
n354 , n355 , n356 , n358 , n359 , n360 , n362 , n363 , n364 , n365 ,
n366 , n367 , n368 , n369 , n372 , n373 , n374 , n376 , n382 , n383 ,
n385 , n388 , n390 , n391 , n392 , n393 , n394 , n395 , n396 , n397 ,
n398 , n399 , n400 , n401 , n402 , n404 , n405 , n406 , n407 , n408 ,
n409 , n410 , n411 , n412 , n414 , n415 , n416 , n418 , n419 , n420 ,
n421 , n422 , n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 ,
n431 , n432 , n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 ,
n441 , n442 , n443 , n444 , n445 , n446 , n447 , n449 , n450 , n451 ,
n452 , n453 , n455 , n458 , n459 , n460 , n461 , n462 , n463 , n464 ,
n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 , n473 , n474 ,
n475 , n477 , n478 , n479 , n480 , n481 , n483 , n484 , n485 , n486 ,
n489 , n490 , n491 , n492 , n493 , n494 , n496 , n497 , n498 , n499 ,
n500 , n501 , n502 , n503 , n505 , n506 , n507 , n508 , n509 , n510 ,
n511 , n512 , n513 , n514 , n515 , n517 , n518 , n519 , n521 , n522 ,
n523 , n524 , n525 , n526 , n527 , n528 , n529 , n531 , n532 , n533 ,
n534 , n535 , n536 , n537 , n538 , n539 , n540 , n543 , n545 , n546 ,
n548 , n549 , n550 , n551 , n552 , n553 , n554 , n555 , n556 , n557 ,
n558 , n559 , n561 , n562 , n563 , n568 , n569 , n570 , n571 , n572 ,
n573 , n575 , n576 , n577 , n578 , n580 , n581 , n582 , n583 , n584 ,
n585 , n586 , n587 , n588 , n589 , n590 , n592 , n593 , n594 , n595 ,
n597 , n598 , n599 , n602 , n603 , n604 , n605 , n607 , n608 , n609 ,
n610 , n612 , n613 , n614 , n615 , n616 , n618 , n619 , n620 , n621 ,
n622 , n624 , n625 , n626 , n628 , n629 , n630 , n631 , n632 , n633 ,
n634 , n637 , n638 , n639 , n640 , n641 , n642 , n644 , n645 , n646 ,
n647 , n648 , n650 , n651 , n652 , n653 , n654 , n655 , n656 , n657 ,
n658 , n659 , n660 , n662 , n663 , n664 , n665 , n666 , n667 , n669 ,
n670 , n671 , n672 , n674 , n675 , n677 , n678 , n679 , n680 , n681 ,
n682 , n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 ,
n692 , n693 , n694 , n695 , n696 , n698 , n699 , n700 , n701 , n702 ,
n703 , n704 , n705 , n706 , n707 , n709 , n710 , n711 , n712 , n713 ,
n716 , n717 , n718 , n719 , n720 , n723 , n724 , n725 , n726 , n727 ,
n728 , n729 , n730 , n731 , n732 , n733 , n734 , n735 , n736 , n737 ,
n738 , n739 , n740 , n741 , n742 , n743 , n744 , n745 , n746 , n747 ,
n748 , n749 , n750 , n751 , n752 , n753 , n755 , n756 , n757 , n759 ,
n761 , n762 , n763 , n764 , n766 , n767 , n768 , n769 , n770 , n771 ,
n772 , n773 , n774 , n775 , n777 , n778 , n780 , n781 , n782 , n783 ,
n784 , n785 , n787 , n788 , n789 , n790 , n791 , n792 , n794 , n795 ,
n796 , n797 , n798 , n799 , n800 , n802 , n803 , n804 , n805 , n806 ,
n808 , n809 , n810 , n811 , n812 , n814 , n815 , n816 , n817 , n818 ,
n819 , n820 , n821 , n822 , n823 , n825 , n826 , n827 , n828 , n829 ,
n831 , n832 , n833 , n834 , n835 , n836 , n837 , n838 , n839 , n842 ,
n843 , n844 , n846 , n847 , n848 , n851 , n852 , n853 , n854 , n855 ,
n856 , n857 , n858 , n859 , n861 , n862 , n863 , n864 , n865 , n866 ,
n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 , n875 , n876 ,
n877 , n879 , n880 , n881 , n883 , n884 , n885 , n886 , n888 , n890 ,
n891 , n892 , n893 , n895 , n896 , n897 , n898 , n899 , n900 , n901 ,
n902 , n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 ,
n913 , n914 , n915 , n916 , n919 , n920 , n921 , n922 , n923 , n924 ,
n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 ,
n935 , n936 , n938 , n939 , n940 , n941 , n942 , n943 , n945 , n947 ,
n948 , n949 , n950 , n952 , n953 , n954 , n956 , n957 , n958 , n959 ,
n960 , n963 , n965 , n968 , n969 , n970 , n972 , n973 , n975 , n976 ,
n977 , n978 , n979 , n980 , n981 , n982 , n983 , n985 , n986 , n987 ,
n988 , n989 , n990 , n991 , n992 , n993 , n994 , n995 , n996 , n997 ,
n998 , n1000 , n1001 , n1002 , n1003 , n1004 , n1005 , n1006 , n1007 , n1008 ,
n1009 , n1010 , n1011 , n1012 , n1013 , n1014 , n1015 , n1017 , n1018 , n1019 ,
n1020 , n1021 , n1022 , n1023 , n1024 , n1025 , n1026 , n1028 , n1029 , n1030 ,
n1031 , n1032 , n1034 , n1035 , n1036 , n1037 , n1038 , n1040 , n1041 , n1042 ,
n1045 , n1046 , n1048 , n1049 , n1051 , n1052 , n1053 , n1054 , n1055 , n1056 ,
n1057 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 , n1066 , n1067 , n1068 ,
n1069 , n1070 , n1071 , n1072 , n1073 , n1074 , n1075 , n1076 , n1077 , n1078 ,
n1079 , n1080 , n1081 , n1082 , n1083 , n1084 , n1085 , n1086 , n1089 , n1090 ,
n1091 , n1092 , n1093 , n1094 , n1098 , n1099 , n1101 , n1102 , n1103 , n1104 ,
n1105 , n1106 , n1107 , n1108 , n1109 , n1111 , n1112 , n1113 , n1114 , n1115 ,
n1116 , n1117 , n1118 , n1120 , n1121 , n1122 , n1123 , n1124 , n1126 , n1127 ,
n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 , n1136 , n1137 , n1138 ,
n1139 , n1141 , n1142 , n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 ,
n1151 , n1152 , n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 ,
n1161 , n1162 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 ,
n1173 , n1174 , n1176 , n1178 , n1179 , n1183 , n1184 , n1185 , n1187 , n1188 ,
n1189 , n1190 , n1191 , n1192 , n1193 , n1194 , n1195 , n1196 , n1197 , n1198 ,
n1199 , n1200 , n1201 , n1202 , n1203 , n1204 , n1206 , n1208 , n1209 , n1210 ,
n1211 , n1212 , n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1220 , n1221 ,
n1222 , n1223 , n1225 , n1226 , n1228 , n1229 , n1230 , n1231 , n1232 , n1234 ,
n1235 , n1236 , n1237 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 , n1245 ,
n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 , n1255 ,
n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 , n1265 ,
n1266 , n1267 , n1268 , n1271 , n1272 , n1273 , n1274 , n1275 , n1276 , n1277 ,
n1278 , n1280 , n1282 , n1283 , n1284 , n1285 , n1286 , n1287 , n1289 , n1290 ,
n1291 , n1292 , n1293 , n1294 , n1295 , n1296 , n1298 , n1300 , n1301 , n1302 ,
n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 ,
n1313 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1323 , n1324 ,
n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 ,
n1335 , n1336 , n1337 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 , n1345 ,
n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1354 , n1356 , n1358 , n1359 ,
n1360 , n1364 , n1365 , n1367 , n1368 , n1369 , n1371 , n1372 , n1373 , n1374 ,
n1375 , n1376 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 , n1385 , n1386 ,
n1387 , n1388 , n1389 , n1392 , n1393 , n1394 , n1395 , n1397 , n1398 , n1399 ,
n1400 , n1401 , n1403 , n1404 , n1405 , n1407 , n1410 , n1411 , n1412 , n1413 ,
n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 ,
n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 , n1437 , n1438 , n1439 ,
n1440 , n1441 , n1442 , n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 ,
n1450 , n1451 , n1452 , n1453 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 ,
n1461 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1472 , n1473 , n1474 ,
n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 ,
n1486 , n1487 , n1488 , n1489 , n1490 , n1492 , n1493 , n1494 , n1496 , n1497 ,
n1499 , n1500 , n1501 , n1502 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 ,
n1512 , n1513 , n1514 , n1516 , n1517 , n1520 , n1521 , n1522 , n1523 , n1524 ,
n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1535 ,
n1536 , n1537 , n1538 , n1539 , n1541 , n1542 , n1544 , n1545 , n1546 , n1547 ,
n1548 , n1549 , n1550 , n1551 , n1552 , n1554 , n1555 , n1556 , n1557 , n1558 ,
n1559 , n1560 , n1561 , n1562 , n1563 , n1564 , n1565 , n1566 , n1567 , n1569 ,
n1570 , n1571 , n1572 , n1573 , n1574 , n1576 , n1577 , n1578 , n1579 , n1580 ,
n1581 , n1582 , n1583 , n1585 , n1586 , n1588 , n1589 , n1590 , n1591 , n1592 ,
n1593 , n1594 , n1595 , n1596 , n1597 , n1599 , n1600 , n1601 , n1602 , n1603 ,
n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1614 ,
n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 ,
n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1634 , n1635 , n1636 , n1637 ,
n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 , n1645 , n1646 , n1647 ,
n1648 , n1650 , n1651 , n1652 , n1653 , n1656 , n1658 , n1659 , n1661 , n1662 ,
n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 ,
n1677 , n1678 , n1679 , n1680 , n1681 , n1683 , n1684 , n1685 , n1686 , n1687 ,
n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 , n1695 , n1696 , n1699 ,
n1701 , n1702 , n1703 , n1704 , n1705 , n1706 , n1709 , n1711 , n1712 , n1713 ,
n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1722 , n1723 , n1724 ,
n1725 , n1726 , n1727 , n1728 , n1730 , n1731 , n1732 , n1734 , n1735 , n1736 ,
n1737 , n1738 , n1739 , n1741 , n1742 , n1744 , n1745 , n1746 , n1747 , n1748 ,
n1749 , n1750 , n1751 , n1752 , n1754 , n1757 , n1758 , n1759 , n1760 , n1762 ,
n1763 , n1764 , n1765 , n1766 , n1767 , n1769 , n1770 , n1771 , n1772 , n1773 ,
n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1781 , n1782 , n1783 , n1785 ,
n1786 , n1787 , n1789 , n1791 , n1792 , n1795 , n1796 , n1797 ;
    nor g0 ( n1319 , n228 , n95 );
    not g1 ( n996 , n1457 );
    nor g2 ( n337 , n220 , n140 );
    nor g3 ( n1099 , n539 , n1022 );
    or g4 ( n464 , n24 , n465 );
    or g5 ( n1648 , n1081 , n1694 );
    or g6 ( n507 , n616 , n68 );
    xnor g7 ( n1741 , n1718 , n1332 );
    and g8 ( n586 , n1103 , n81 );
    nor g9 ( n1600 , n1618 , n807 );
    or g10 ( n1442 , n1439 , n1316 );
    or g11 ( n1011 , n186 , n1027 );
    or g12 ( n1782 , n1690 , n1694 );
    and g13 ( n1306 , n723 , n1251 );
    not g14 ( n491 , n1397 );
    xnor g15 ( n1677 , n525 , n578 );
    or g16 ( n1034 , n588 , n1497 );
    or g17 ( n1603 , n627 , n964 );
    or g18 ( n1090 , n1146 , n1407 );
    nor g19 ( n237 , n261 , n1028 );
    and g20 ( n562 , n842 , n356 );
    or g21 ( n840 , n452 , n421 );
    and g22 ( n218 , n1668 , n590 );
    nor g23 ( n1040 , n1395 , n354 );
    nor g24 ( n24 , n44 , n282 );
    or g25 ( n890 , n579 , n150 );
    and g26 ( n1171 , n99 , n1531 );
    xnor g27 ( n670 , n1435 , n1043 );
    nor g28 ( n1237 , n1788 , n1457 );
    or g29 ( n551 , n579 , n1189 );
    or g30 ( n1469 , n186 , n75 );
    nor g31 ( n932 , n261 , n281 );
    nor g32 ( n1221 , n378 , n1268 );
    or g33 ( n1548 , n186 , n370 );
    buf g34 ( n399 , n1326 );
    nor g35 ( n674 , n261 , n1746 );
    not g36 ( n1003 , n903 );
    not g37 ( n1720 , n240 );
    or g38 ( n48 , n669 , n77 );
    or g39 ( n1533 , n307 , n964 );
    and g40 ( n63 , n1391 , n713 );
    and g41 ( n1110 , n215 , n1764 );
    nor g42 ( n1679 , n473 , n1480 );
    nor g43 ( n166 , n1660 , n714 );
    or g44 ( n1480 , n1301 , n214 );
    nor g45 ( n1616 , n378 , n324 );
    not g46 ( n1597 , n884 );
    nor g47 ( n436 , n1765 , n219 );
    nor g48 ( n503 , n193 , n1662 );
    not g49 ( n1433 , n1039 );
    xnor g50 ( n557 , n1619 , n1555 );
    xnor g51 ( n1048 , n550 , n685 );
    xnor g52 ( n1035 , n778 , n1294 );
    not g53 ( n1766 , n1545 );
    buf g54 ( n1697 , n1414 );
    not g55 ( n1550 , n1085 );
    nor g56 ( n1614 , n1281 , n339 );
    nor g57 ( n1023 , n188 , n807 );
    not g58 ( n561 , n1506 );
    buf g59 ( n862 , n909 );
    and g60 ( n1046 , n1235 , n1636 );
    or g61 ( n1528 , n1295 , n947 );
    and g62 ( n518 , n302 , n1244 );
    and g63 ( n1437 , n396 , n55 );
    nor g64 ( n1179 , n44 , n881 );
    or g65 ( n1722 , n186 , n1314 );
    or g66 ( n891 , n627 , n1110 );
    not g67 ( n428 , n538 );
    or g68 ( n1318 , n307 , n1710 );
    not g69 ( n134 , n1172 );
    or g70 ( n1290 , n213 , n613 );
    not g71 ( n1750 , n1437 );
    nor g72 ( n1452 , n44 , n1563 );
    buf g73 ( n1355 , n288 );
    or g74 ( n700 , n307 , n905 );
    nor g75 ( n67 , n402 , n544 );
    or g76 ( n397 , n1106 , n1257 );
    or g77 ( n137 , n1205 , n964 );
    nor g78 ( n1458 , n377 , n701 );
    or g79 ( n175 , n764 , n1200 );
    or g80 ( n1060 , n462 , n1694 );
    nor g81 ( n202 , n669 , n504 );
    or g82 ( n1693 , n1205 , n1027 );
    or g83 ( n838 , n1072 , n1694 );
    nor g84 ( n770 , n862 , n355 );
    nor g85 ( n160 , n560 , n1018 );
    and g86 ( n242 , n139 , n436 );
    or g87 ( n286 , n1147 , n1749 );
    nor g88 ( n232 , n200 , n288 );
    or g89 ( n1761 , n1684 , n762 );
    nor g90 ( n133 , n1172 , n1519 );
    nor g91 ( n944 , n220 , n70 );
    or g92 ( n1460 , n1146 , n698 );
    nor g93 ( n1667 , n579 , n647 );
    or g94 ( n95 , n1205 , n168 );
    nor g95 ( n1520 , n1241 , n1585 );
    or g96 ( n1692 , n1113 , n998 );
    or g97 ( n1438 , n990 , n1200 );
    nor g98 ( n1158 , n704 , n144 );
    nor g99 ( n251 , n1681 , n479 );
    or g100 ( n805 , n1205 , n370 );
    and g101 ( n476 , n1613 , n1716 );
    nor g102 ( n746 , n560 , n1011 );
    xnor g103 ( n1051 , n428 , n916 );
    nor g104 ( n1670 , n560 , n1380 );
    nor g105 ( n1627 , n94 , n1215 );
    buf g106 ( n845 , n1613 );
    nor g107 ( n208 , n946 , n714 );
    and g108 ( n469 , n73 , n575 );
    or g109 ( n369 , n579 , n562 );
    and g110 ( n628 , n2 , n1204 );
    or g111 ( n1772 , n1744 , n229 );
    xnor g112 ( n266 , n654 , n1741 );
    or g113 ( n1285 , n694 , n227 );
    or g114 ( n1012 , n1295 , n1793 );
    or g115 ( n595 , n186 , n487 );
    or g116 ( n950 , n1295 , n1010 );
    or g117 ( n1508 , n651 , n942 );
    not g118 ( n1785 , n1598 );
    xnor g119 ( n1669 , n412 , n1108 );
    nor g120 ( n759 , n1580 , n1330 );
    nor g121 ( n366 , n853 , n1118 );
    or g122 ( n826 , n1280 , n394 );
    or g123 ( n1304 , n398 , n1694 );
    or g124 ( n735 , n1792 , n628 );
    and g125 ( n191 , n1585 , n1545 );
    nor g126 ( n429 , n378 , n1111 );
    or g127 ( n91 , n780 , n1440 );
    nor g128 ( n1403 , n1166 , n319 );
    not g129 ( n907 , n89 );
    or g130 ( n505 , n1349 , n1562 );
    or g131 ( n1145 , n63 , n176 );
    nor g132 ( n1291 , n1755 , n343 );
    and g133 ( n828 , n1660 , n1288 );
    not g134 ( n23 , n286 );
    nor g135 ( n110 , n1335 , n797 );
    not g136 ( n1676 , n1338 );
    or g137 ( n1297 , n203 , n349 );
    or g138 ( n842 , n298 , n1190 );
    not g139 ( n880 , n1226 );
    and g140 ( n741 , n147 , n1626 );
    or g141 ( n435 , n749 , n585 );
    and g142 ( n75 , n1453 , n241 );
    and g143 ( n1604 , n1235 , n252 );
    or g144 ( n1428 , n1374 , n1524 );
    or g145 ( n1546 , n1295 , n1422 );
    or g146 ( n1260 , n627 , n168 );
    or g147 ( n1410 , n206 , n879 );
    or g148 ( n361 , n1116 , n1692 );
    nor g149 ( n1541 , n377 , n1714 );
    or g150 ( n1341 , n1473 , n1211 );
    not g151 ( n345 , n1391 );
    not g152 ( n774 , n1663 );
    or g153 ( n215 , n1146 , n156 );
    and g154 ( n1369 , n703 , n243 );
    not g155 ( n669 , n617 );
    or g156 ( n130 , n1523 , n770 );
    xnor g157 ( n1647 , n517 , n1445 );
    nor g158 ( n1691 , n579 , n1145 );
    or g159 ( n1282 , n1298 , n579 );
    xnor g160 ( n666 , n526 , n1217 );
    or g161 ( n888 , n774 , n1694 );
    nor g162 ( n856 , n1032 , n1129 );
    and g163 ( n1244 , n777 , n185 );
    and g164 ( n259 , n732 , n858 );
    not g165 ( n1696 , n147 );
    or g166 ( n211 , n1602 , n605 );
    or g167 ( n1292 , n1618 , n1312 );
    or g168 ( n1066 , n1205 , n259 );
    or g169 ( n121 , n1384 , n1571 );
    or g170 ( n656 , n1482 , n480 );
    not g171 ( n1615 , n1097 );
    or g172 ( n1252 , n1054 , n268 );
    or g173 ( n1496 , n307 , n1346 );
    nor g174 ( n388 , n560 , n310 );
    or g175 ( n1524 , n348 , n283 );
    nor g176 ( n1622 , n1681 , n1363 );
    or g177 ( n698 , n1488 , n579 );
    or g178 ( n85 , n1419 , n1694 );
    and g179 ( n373 , n1037 , n65 );
    or g180 ( n223 , n982 , n1561 );
    nor g181 ( n1287 , n44 , n877 );
    nor g182 ( n1007 , n380 , n1227 );
    or g183 ( n784 , n271 , n1512 );
    or g184 ( n1412 , n857 , n809 );
    not g185 ( n332 , n758 );
    and g186 ( n168 , n74 , n712 );
    nor g187 ( n347 , n472 , n591 );
    not g188 ( n437 , n12 );
    not g189 ( n936 , n1171 );
    nor g190 ( n143 , n1162 , n1572 );
    nor g191 ( n647 , n353 , n1003 );
    not g192 ( n1681 , n1281 );
    nor g193 ( n1431 , n1600 , n1748 );
    or g194 ( n1509 , n1146 , n1282 );
    or g195 ( n975 , n338 , n1234 );
    or g196 ( n184 , n828 , n1398 );
    nor g197 ( n1141 , n545 , n1309 );
    or g198 ( n974 , n709 , n1290 );
    nor g199 ( n1202 , n832 , n708 );
    or g200 ( n1167 , n435 , n91 );
    and g201 ( n585 , n495 , n426 );
    or g202 ( n461 , n992 , n22 );
    nor g203 ( n1744 , n1162 , n908 );
    xnor g204 ( n1283 , n1249 , n1 );
    or g205 ( n1185 , n344 , n695 );
    nor g206 ( n330 , n1713 , n807 );
    and g207 ( n57 , n1146 , n1400 );
    or g208 ( n519 , n1295 , n1779 );
    not g209 ( n1661 , n1047 );
    nor g210 ( n512 , n228 , n1187 );
    nor g211 ( n443 , n1281 , n254 );
    and g212 ( n494 , n1125 , n76 );
    nor g213 ( n90 , n1162 , n874 );
    and g214 ( n295 , n1135 , n407 );
    not g215 ( n539 , n560 );
    nor g216 ( n1206 , n261 , n1494 );
    nor g217 ( n1745 , n261 , n1758 );
    or g218 ( n317 , n1536 , n276 );
    nor g219 ( n1731 , n1591 , n1642 );
    or g220 ( n691 , n1295 , n960 );
    or g221 ( n183 , n1670 , n533 );
    or g222 ( n49 , n675 , n1146 );
    or g223 ( n230 , n1375 , n1200 );
    or g224 ( n1718 , n930 , n232 );
    or g225 ( n82 , n1417 , n579 );
    not g226 ( n1429 , n708 );
    nor g227 ( n1711 , n1755 , n592 );
    not g228 ( n398 , n606 );
    or g229 ( n432 , n1334 , n1694 );
    and g230 ( n1087 , n1460 , n292 );
    nor g231 ( n1184 , n378 , n608 );
    or g232 ( n1333 , n1429 , n614 );
    xnor g233 ( n1415 , n438 , n825 );
    not g234 ( n1041 , n482 );
    nor g235 ( n1724 , n378 , n113 );
    not g236 ( n956 , n1279 );
    nor g237 ( n277 , n560 , n305 );
    not g238 ( n1147 , n1406 );
    nor g239 ( n930 , n710 , n614 );
    xnor g240 ( n903 , n1093 , n1329 );
    nor g241 ( n572 , n966 , n1227 );
    and g242 ( n1257 , n396 , n1795 );
    not g243 ( n61 , n1503 );
    nor g244 ( n511 , n560 , n1424 );
    or g245 ( n1188 , n1105 , n1043 );
    not g246 ( n1642 , n278 );
    nor g247 ( n1254 , n378 , n1603 );
    nor g248 ( n1153 , n832 , n1043 );
    nor g249 ( n1763 , n438 , n1569 );
    or g250 ( n768 , n821 , n268 );
    nor g251 ( n1082 , n579 , n1672 );
    or g252 ( n699 , n442 , n1589 );
    or g253 ( n679 , n50 , n903 );
    not g254 ( n1026 , n326 );
    and g255 ( n744 , n1426 , n600 );
    or g256 ( n194 , n781 , n1312 );
    and g257 ( n447 , n1515 , n591 );
    nor g258 ( n1739 , n1155 , n1594 );
    nor g259 ( n453 , n748 , n1288 );
    nor g260 ( n22 , n1166 , n1238 );
    not g261 ( n1264 , n19 );
    nor g262 ( n1261 , n1388 , n438 );
    or g263 ( n192 , n191 , n1566 );
    and g264 ( n570 , n895 , n1079 );
    or g265 ( n417 , n972 , n997 );
    and g266 ( n659 , n1402 , n929 );
    and g267 ( n671 , n60 , n1121 );
    not g268 ( n250 , n548 );
    or g269 ( n1064 , n1690 , n1200 );
    nor g270 ( n465 , n378 , n1036 );
    nor g271 ( n513 , n743 , n820 );
    or g272 ( n1726 , n311 , n763 );
    and g273 ( n649 , n1613 , n915 );
    nor g274 ( n906 , n523 , n504 );
    nor g275 ( n1209 , n1553 , n721 );
    nor g276 ( n1056 , n625 , n674 );
    xnor g277 ( n526 , n711 , n719 );
    and g278 ( n1160 , n909 , n280 );
    and g279 ( n1773 , n946 , n1118 );
    nor g280 ( n446 , n44 , n1154 );
    not g281 ( n532 , n403 );
    and g282 ( n485 , n996 , n1356 );
    or g283 ( n1246 , n1205 , n454 );
    or g284 ( n210 , n25 , n609 );
    not g285 ( n1358 , n1718 );
    not g286 ( n439 , n504 );
    nor g287 ( n1747 , n200 , n319 );
    or g288 ( n1268 , n957 , n1200 );
    or g289 ( n34 , n326 , n1590 );
    and g290 ( n176 , n1607 , n536 );
    xnor g291 ( n678 , n428 , n467 );
    xor g292 ( n878 , n1131 , n364 );
    or g293 ( n664 , n186 , n905 );
    or g294 ( n100 , n472 , n77 );
    or g295 ( n652 , n1466 , n359 );
    or g296 ( n1148 , n307 , n1087 );
    and g297 ( n1010 , n1446 , n317 );
    or g298 ( n374 , n1295 , n1002 );
    and g299 ( n552 , n342 , n1524 );
    and g300 ( n300 , n228 , n1078 );
    or g301 ( n1127 , n252 , n835 );
    or g302 ( n734 , n1295 , n1025 );
    or g303 ( n231 , n1089 , n667 );
    nor g304 ( n827 , n1162 , n873 );
    nor g305 ( n707 , n200 , n708 );
    nor g306 ( n515 , n228 , n289 );
    or g307 ( n783 , n602 , n1061 );
    buf g308 ( n235 , n1721 );
    or g309 ( n400 , n1574 , n1413 );
    not g310 ( n802 , n715 );
    nor g311 ( n1594 , n261 , n796 );
    or g312 ( n1053 , n627 , n75 );
    and g313 ( n456 , n1509 , n1539 );
    nor g314 ( n161 , n1146 , n1686 );
    or g315 ( n109 , n1295 , n427 );
    nor g316 ( n650 , n1681 , n437 );
    or g317 ( n127 , n1280 , n1208 );
    xnor g318 ( n578 , n1070 , n652 );
    and g319 ( n808 , n1244 , n645 );
    and g320 ( n1787 , n1045 , n484 );
    nor g321 ( n925 , n1435 , n714 );
    or g322 ( n1017 , n1464 , n1662 );
    xnor g323 ( n1143 , n719 , n1623 );
    nor g324 ( n340 , n539 , n1671 );
    nor g325 ( n1532 , n209 , n87 );
    or g326 ( n661 , n72 , n102 );
    nor g327 ( n1274 , n377 , n1601 );
    nor g328 ( n1599 , n378 , n180 );
    nor g329 ( n725 , n44 , n1005 );
    and g330 ( n124 , n1588 , n309 );
    or g331 ( n909 , n154 , n1226 );
    and g332 ( n213 , n1146 , n1628 );
    nor g333 ( n45 , n627 , n123 );
    or g334 ( n1037 , n523 , n1312 );
    xnor g335 ( n1130 , n1401 , n1391 );
    and g336 ( n1250 , n60 , n1070 );
    not g337 ( n1128 , n676 );
    and g338 ( n673 , n703 , n859 );
    or g339 ( n1447 , n1771 , n1184 );
    or g340 ( n52 , n1797 , n876 );
    and g341 ( n1107 , n1518 , n1662 );
    or g342 ( n290 , n1169 , n268 );
    nor g343 ( n1086 , n1166 , n1729 );
    not g344 ( n1013 , n1104 );
    or g345 ( n1571 , n825 , n548 );
    nor g346 ( n798 , n472 , n807 );
    or g347 ( n959 , n159 , n752 );
    or g348 ( n182 , n789 , n62 );
    nor g349 ( n773 , n539 , n1730 );
    xnor g350 ( n884 , n624 , n558 );
    nor g351 ( n214 , n1395 , n308 );
    not g352 ( n990 , n830 );
    not g353 ( n1527 , n1463 );
    xnor g354 ( n933 , n818 , n14 );
    nor g355 ( n199 , n378 , n1644 );
    not g356 ( n268 , n307 );
    or g357 ( n823 , n1191 , n814 );
    xnor g358 ( n1059 , n820 , n711 );
    or g359 ( n1247 , n1757 , n511 );
    not g360 ( n1654 , n457 );
    and g361 ( n1620 , n39 , n1508 );
    or g362 ( n817 , n1341 , n993 );
    not g363 ( n150 , n265 );
    not g364 ( n1451 , n342 );
    or g365 ( n607 , n1146 , n441 );
    nor g366 ( n1270 , n220 , n80 );
    or g367 ( n618 , n764 , n1694 );
    nor g368 ( n1301 , n228 , n1214 );
    nor g369 ( n249 , n220 , n1371 );
    not g370 ( n1775 , n1135 );
    or g371 ( n1607 , n748 , n77 );
    nor g372 ( n726 , n228 , n833 );
    not g373 ( n1307 , n1180 );
    or g374 ( n1154 , n627 , n259 );
    and g375 ( n94 , n1146 , n1691 );
    and g376 ( n255 , n1388 , n1569 );
    or g377 ( n816 , n1074 , n478 );
    and g378 ( n499 , n1436 , n504 );
    nor g379 ( n103 , n560 , n1469 );
    and g380 ( n383 , n961 , n504 );
    xnor g381 ( n1619 , n1226 , n154 );
    or g382 ( n555 , n450 , n579 );
    nor g383 ( n712 , n724 , n1529 );
    or g384 ( n1446 , n260 , n192 );
    and g385 ( n1047 , n92 , n457 );
    or g386 ( n655 , n1775 , n1086 );
    xnor g387 ( n1397 , n1241 , n1790 );
    or g388 ( n2 , n956 , n1774 );
    nor g389 ( n1634 , n954 , n869 );
    or g390 ( n1077 , n1241 , n1160 );
    or g391 ( n1063 , n117 , n53 );
    or g392 ( n152 , n307 , n454 );
    or g393 ( n1716 , n1490 , n40 );
    xnor g394 ( n1161 , n708 , n1660 );
    or g395 ( n421 , n1541 , n108 );
    and g396 ( n1473 , n851 , n1091 );
    nor g397 ( n1474 , n1238 , n1227 );
    nor g398 ( n794 , n228 , n279 );
    nor g399 ( n165 , n240 , n1389 );
    buf g400 ( n173 , n84 );
    or g401 ( n574 , n1703 , n117 );
    or g402 ( n98 , n1146 , n1340 );
    nor g403 ( n1539 , n1258 , n164 );
    nor g404 ( n25 , n1395 , n838 );
    nor g405 ( n42 , n560 , n1478 );
    or g406 ( n1737 , n1383 , n1542 );
    not g407 ( n1690 , n1033 );
    or g408 ( n372 , n579 , n1358 );
    not g409 ( n1152 , n747 );
    not g410 ( n920 , n485 );
    not g411 ( n41 , n984 );
    nor g412 ( n857 , n481 , n151 );
    nor g413 ( n1350 , n134 , n1288 );
    or g414 ( n474 , n626 , n791 );
    or g415 ( n812 , n583 , n1552 );
    buf g416 ( n430 , n1645 );
    nor g417 ( n1224 , n368 , n1537 );
    not g418 ( n227 , n186 );
    nor g419 ( n588 , n1395 , n1648 );
    or g420 ( n1157 , n388 , n376 );
    not g421 ( n1295 , n579 );
    or g422 ( n987 , n1146 , n1259 );
    xnor g423 ( n364 , n868 , n1161 );
    xnor g424 ( n271 , n1235 , n1231 );
    nor g425 ( n1651 , n1435 , n1227 );
    nor g426 ( n31 , n377 , n178 );
    not g427 ( n44 , n378 );
    or g428 ( n333 , n579 , n28 );
    xnor g429 ( n278 , n35 , n1386 );
    or g430 ( n1343 , n445 , n1725 );
    or g431 ( n65 , n1105 , n319 );
    nor g432 ( n577 , n656 , n198 );
    nor g433 ( n1529 , n261 , n931 );
    nor g434 ( n1000 , n1162 , n522 );
    or g435 ( n693 , n864 , n815 );
    or g436 ( n506 , n1350 , n731 );
    nor g437 ( n1784 , n220 , n1328 );
    xnor g438 ( n1093 , n1664 , n466 );
    or g439 ( n1481 , n11 , n160 );
    or g440 ( n958 , n847 , n1514 );
    not g441 ( n865 , n962 );
    xnor g442 ( n320 , n933 , n26 );
    or g443 ( n407 , n963 , n221 );
    nor g444 ( n1547 , n1166 , n1660 );
    or g445 ( n993 , n265 , n1347 );
    nor g446 ( n1717 , n261 , n519 );
    or g447 ( n685 , n499 , n906 );
    and g448 ( n1440 , n495 , n552 );
    and g449 ( n1321 , n966 , n1662 );
    nor g450 ( n391 , n748 , n591 );
    nor g451 ( n935 , n1618 , n591 );
    or g452 ( n385 , n1136 , n419 );
    or g453 ( n824 , n5 , n1759 );
    not g454 ( n395 , n1435 );
    and g455 ( n811 , n1135 , n550 );
    or g456 ( n790 , n1250 , n174 );
    xnor g457 ( n1085 , n667 , n273 );
    or g458 ( n1094 , n1476 , n1777 );
    and g459 ( n587 , n946 , n614 );
    or g460 ( n1630 , n1696 , n1571 );
    nor g461 ( n780 , n495 , n1174 );
    or g462 ( n1124 , n186 , n1710 );
    xnor g463 ( n1762 , n1293 , n1051 );
    or g464 ( n1407 , n1210 , n579 );
    or g465 ( n1065 , n220 , n242 );
    or g466 ( n1008 , n307 , n259 );
    nor g467 ( n785 , n377 , n1533 );
    xnor g468 ( n195 , n740 , n313 );
    or g469 ( n1430 , n844 , n1694 );
    nor g470 ( n536 , n1391 , n1526 );
    nor g471 ( n943 , n1700 , n1281 );
    nor g472 ( n344 , n228 , n137 );
    and g473 ( n810 , n1125 , n580 );
    or g474 ( n799 , n1477 , n655 );
    nor g475 ( n787 , n378 , n969 );
    nor g476 ( n138 , n756 , n1521 );
    and g477 ( n1061 , n100 , n1291 );
    not g478 ( n1286 , n1768 );
    or g479 ( n1401 , n589 , n425 );
    or g480 ( n1096 , n693 , n1410 );
    not g481 ( n234 , n711 );
    nor g482 ( n1323 , n200 , n1729 );
    nor g483 ( n1544 , n1713 , n591 );
    or g484 ( n701 , n307 , n1495 );
    not g485 ( n1190 , n1288 );
    not g486 ( n1081 , n335 );
    or g487 ( n1296 , n332 , n1694 );
    and g488 ( n1557 , n319 , n591 );
    or g489 ( n1116 , n148 , n1364 );
    or g490 ( n1273 , n251 , n1614 );
    not g491 ( n357 , n566 );
    xnor g492 ( n207 , n325 , n1582 );
    not g493 ( n1253 , n9 );
    or g494 ( n309 , n1004 , n1302 );
    nor g495 ( n224 , n377 , n1530 );
    nor g496 ( n902 , n44 , n1277 );
    or g497 ( n948 , n428 , n920 );
    or g498 ( n1265 , n1307 , n1200 );
    and g499 ( n1584 , n1613 , n912 );
    or g500 ( n1022 , n186 , n469 );
    not g501 ( n481 , n147 );
    or g502 ( n1475 , n1205 , n469 );
    or g503 ( n722 , n1772 , n1344 );
    nor g504 ( n1665 , n377 , n365 );
    or g505 ( n269 , n579 , n1196 );
    and g506 ( n620 , n904 , n822 );
    not g507 ( n1200 , n627 );
    or g508 ( n1457 , n733 , n848 );
    or g509 ( n1543 , n1343 , n834 );
    not g510 ( n1164 , n276 );
    or g511 ( n1220 , n718 , n726 );
    nor g512 ( n819 , n1570 , n1283 );
    or g513 ( n1656 , n186 , n259 );
    nor g514 ( n350 , n380 , n721 );
    nor g515 ( n406 , n1395 , n1709 );
    buf g516 ( n542 , n84 );
    or g517 ( n1348 , n1295 , n1578 );
    not g518 ( n710 , n288 );
    not g519 ( n632 , n510 );
    nor g520 ( n229 , n377 , n314 );
    and g521 ( n351 , n1292 , n17 );
    or g522 ( n875 , n111 , n227 );
    nor g523 ( n1309 , n1039 , n1223 );
    nor g524 ( n745 , n1669 , n390 );
    nor g525 ( n1186 , n220 , n1317 );
    or g526 ( n646 , n455 , n1567 );
    nor g527 ( n792 , n1281 , n1020 );
    xnor g528 ( n534 , n580 , n1125 );
    and g529 ( n43 , n1279 , n1289 );
    or g530 ( n1129 , n1599 , n1062 );
    not g531 ( n1280 , n1755 );
    or g532 ( n1390 , n78 , n1641 );
    nor g533 ( n325 , n540 , n1711 );
    not g534 ( n1591 , n266 );
    nor g535 ( n814 , n228 , n432 );
    nor g536 ( n533 , n539 , n336 );
    or g537 ( n524 , n1402 , n373 );
    or g538 ( n1316 , n169 , n1403 );
    or g539 ( n1684 , n1500 , n1556 );
    nor g540 ( n527 , n261 , n890 );
    nor g541 ( n1778 , n261 , n1348 );
    and g542 ( n941 , n643 , n1662 );
    not g543 ( n263 , n1125 );
    xnor g544 ( n1 , n940 , n122 );
    nor g545 ( n1421 , n1448 , n414 );
    nor g546 ( n114 , n745 , n167 );
    not g547 ( n1570 , n0 );
    or g548 ( n120 , n188 , n1312 );
    nor g549 ( n1420 , n472 , n1288 );
    or g550 ( n1491 , n1286 , n1574 );
    or g551 ( n929 , n1557 , n163 );
    not g552 ( n280 , n1236 );
    or g553 ( n873 , n307 , n1631 );
    xnor g554 ( n431 , n1342 , n1783 );
    nor g555 ( n20 , n272 , n1763 );
    or g556 ( n363 , n1573 , n1031 );
    or g557 ( n3 , n1126 , n268 );
    or g558 ( n594 , n1146 , n563 );
    or g559 ( n1174 , n1041 , n1451 );
    or g560 ( n1596 , n569 , n327 );
    and g561 ( n205 , n1017 , n1472 );
    nor g562 ( n1699 , n669 , n1288 );
    and g563 ( n886 , n1019 , n1188 );
    or g564 ( n416 , n512 , n181 );
    or g565 ( n73 , n1194 , n1146 );
    nor g566 ( n1345 , n261 , n622 );
    nor g567 ( n1552 , n706 , n867 );
    not g568 ( n486 , n850 );
    nor g569 ( n1497 , n228 , n153 );
    or g570 ( n1337 , n395 , n1312 );
    nor g571 ( n181 , n1395 , n1073 );
    and g572 ( n602 , n1755 , n69 );
    or g573 ( n204 , n1081 , n1200 );
    or g574 ( n747 , n529 , n54 );
    nor g575 ( n226 , n560 , n664 );
    nor g576 ( n56 , n220 , n1399 );
    nor g577 ( n898 , n617 , n1519 );
    or g578 ( n1272 , n23 , n106 );
    not g579 ( n549 , n1579 );
    not g580 ( n675 , n321 );
    and g581 ( n716 , n1435 , n1288 );
    nor g582 ( n1339 , n1175 , n644 );
    nor g583 ( n1794 , n220 , n1723 );
    or g584 ( n1537 , n1596 , n1467 );
    nor g585 ( n1611 , n378 , n1064 );
    buf g586 ( n1425 , n1534 );
    nor g587 ( n1639 , n1162 , n1148 );
    or g588 ( n1121 , n1549 , n1202 );
    xnor g589 ( n1131 , n1284 , n177 );
    nor g590 ( n592 , n798 , n672 );
    nor g591 ( n1723 , n210 , n1159 );
    or g592 ( n1695 , n23 , n880 );
    nor g593 ( n498 , n560 , n597 );
    not g594 ( n1118 , n591 );
    and g595 ( n148 , n579 , n261 );
    or g596 ( n393 , n988 , n820 );
    nor g597 ( n1441 , n378 , n1053 );
    xnor g598 ( n1386 , n1638 , n581 );
    or g599 ( n493 , n1585 , n1719 );
    nor g600 ( n1517 , n228 , n888 );
    or g601 ( n281 , n1295 , n870 );
    nor g602 ( n1617 , n377 , n1576 );
    not g603 ( n1736 , n1313 );
    nor g604 ( n1637 , n1162 , n290 );
    nor g605 ( n786 , n220 , n1505 );
    not g606 ( n1492 , n668 );
    nor g607 ( n1770 , n593 , n201 );
    nor g608 ( n970 , n377 , n1071 );
    xnor g609 ( n719 , n901 , n697 );
    nor g610 ( n426 , n342 , n491 );
    and g611 ( n626 , n1391 , n1401 );
    xnor g612 ( n654 , n1535 , n1423 );
    or g613 ( n1567 , n1423 , n1014 );
    xnor g614 ( n177 , n1729 , n319 );
    or g615 ( n1248 , n952 , n268 );
    or g616 ( n1183 , n458 , n43 );
    and g617 ( n1144 , n1143 , n820 );
    or g618 ( n1625 , n1205 , n1346 );
    or g619 ( n1601 , n1178 , n268 );
    or g620 ( n1641 , n1305 , n692 );
    or g621 ( n1042 , n197 , n268 );
    not g622 ( n853 , n1043 );
    or g623 ( n575 , n1564 , n299 );
    or g624 ( n1149 , n1286 , n1222 );
    nor g625 ( n1328 , n823 , n653 );
    or g626 ( n1530 , n307 , n1314 );
    nor g627 ( n475 , n1125 , n27 );
    xnor g628 ( n302 , n652 , n1575 );
    and g629 ( n743 , n159 , n752 );
    and g630 ( n1168 , n194 , n604 );
    or g631 ( n101 , n223 , n1030 );
    or g632 ( n1032 , n1404 , n1611 );
    and g633 ( n1234 , n1674 , n439 );
    not g634 ( n531 , n896 );
    or g635 ( n365 , n307 , n75 );
    or g636 ( n368 , n737 , n1144 );
    nor g637 ( n831 , n1498 , n1519 );
    or g638 ( n945 , n1046 , n1114 );
    xnor g639 ( n1029 , n1160 , n1695 );
    and g640 ( n1439 , n319 , n1288 );
    xnor g641 ( n1512 , n1130 , n945 );
    and g642 ( n483 , n600 , n541 );
    or g643 ( n301 , n1146 , n1057 );
    or g644 ( n623 , n1622 , n1063 );
    nor g645 ( n672 , n1553 , n714 );
    nor g646 ( n30 , n378 , n142 );
    or g647 ( n1735 , n900 , n227 );
    buf g648 ( n66 , n389 );
    or g649 ( n899 , n490 , n227 );
    nor g650 ( n1757 , n539 , n728 );
    nor g651 ( n651 , n669 , n1118 );
    not g652 ( n1044 , n918 );
    and g653 ( n546 , n1204 , n884 );
    not g654 ( n667 , n88 );
    or g655 ( n728 , n1522 , n227 );
    or g656 ( n795 , n295 , n346 );
    and g657 ( n848 , n1515 , n1662 );
    xnor g658 ( n1468 , n216 , n509 );
    nor g659 ( n1728 , n472 , n504 );
    xnor g660 ( n216 , n686 , n39 );
    xnor g661 ( n1294 , n288 , n1518 );
    or g662 ( n240 , n334 , n800 );
    and g663 ( n1376 , n48 , n727 );
    buf g664 ( n129 , n566 );
    not g665 ( n537 , n841 );
    or g666 ( n1769 , n1773 , n638 );
    or g667 ( n1236 , n493 , n430 );
    not g668 ( n155 , n1636 );
    xnor g669 ( n360 , n534 , n1457 );
    nor g670 ( n1191 , n1395 , n618 );
    or g671 ( n1389 , n415 , n855 );
    nor g672 ( n704 , n261 , n369 );
    or g673 ( n782 , n990 , n1694 );
    or g674 ( n1311 , n1295 , n1085 );
    or g675 ( n354 , n1205 , n456 );
    or g676 ( n522 , n1689 , n268 );
    not g677 ( n1370 , n92 );
    or g678 ( n136 , n610 , n293 );
    or g679 ( n1786 , n1628 , n131 );
    nor g680 ( n753 , n186 , n123 );
    or g681 ( n922 , n117 , n943 );
    or g682 ( n1228 , n503 , n444 );
    or g683 ( n72 , n96 , n1262 );
    and g684 ( n500 , n531 , n43 );
    nor g685 ( n53 , n257 , n1281 );
    nor g686 ( n253 , n1162 , n470 );
    or g687 ( n1036 , n1419 , n1200 );
    xnor g688 ( n468 , n1672 , n1770 );
    nor g689 ( n1112 , n1162 , n1248 );
    nor g690 ( n32 , n748 , n807 );
    or g691 ( n452 , n1637 , n1459 );
    nor g692 ( n316 , n1395 , n1683 );
    or g693 ( n115 , n1791 , n268 );
    not g694 ( n571 , n1175 );
    not g695 ( n382 , n195 );
    buf g696 ( n1504 , n1326 );
    not g697 ( n1417 , n813 );
    or g698 ( n803 , n340 , n911 );
    nor g699 ( n418 , n757 , n590 );
    not g700 ( n1713 , n1498 );
    not g701 ( n1793 , n1524 );
    or g702 ( n633 , n702 , n1200 );
    nor g703 ( n285 , n1395 , n4 );
    and g704 ( n1204 , n121 , n20 );
    and g705 ( n681 , n1485 , n504 );
    and g706 ( n291 , n1545 , n909 );
    or g707 ( n74 , n1146 , n1303 );
    and g708 ( n283 , n1256 , n1706 );
    nor g709 ( n629 , n377 , n1042 );
    nor g710 ( n348 , n1565 , n1566 );
    nor g711 ( n1797 , n560 , n1722 );
    or g712 ( n509 , n741 , n809 );
    not g713 ( n298 , n238 );
    nor g714 ( n1561 , n560 , n1285 );
    nor g715 ( n144 , n261 , n691 );
    not g716 ( n1049 , n663 );
    and g717 ( n1466 , n801 , n504 );
    or g718 ( n713 , n453 , n350 );
    not g719 ( n703 , n1327 );
    nor g720 ( n750 , n380 , n714 );
    and g721 ( n1314 , n987 , n861 );
    nor g722 ( n724 , n261 , n551 );
    and g723 ( n1708 , n562 , n46 );
    and g724 ( n267 , n1337 , n1434 );
    nor g725 ( n1365 , n560 , n968 );
    nor g726 ( n885 , n378 , n1006 );
    and g727 ( n401 , n209 , n1235 );
    not g728 ( n1235 , n149 );
    not g729 ( n254 , n1299 );
    and g730 ( n346 , n1137 , n410 );
    nor g731 ( n872 , n1175 , n546 );
    or g732 ( n1629 , n1054 , n227 );
    and g733 ( n1449 , n120 , n769 );
    or g734 ( n855 , n687 , n1428 );
    or g735 ( n331 , n669 , n614 );
    or g736 ( n1572 , n1128 , n268 );
    xnor g737 ( n818 , n1585 , n1241 );
    or g738 ( n605 , n103 , n1525 );
    or g739 ( n327 , n1550 , n1506 );
    xnor g740 ( n89 , n1226 , n1566 );
    nor g741 ( n1521 , n261 , n1193 );
    not g742 ( n112 , n448 );
    or g743 ( n324 , n462 , n1200 );
    and g744 ( n107 , n1672 , n1331 );
    xnor g745 ( n1217 , n243 , n1623 );
    nor g746 ( n459 , n233 , n1320 );
    and g747 ( n68 , n946 , n1662 );
    nor g748 ( n879 , n1162 , n1318 );
    or g749 ( n767 , n843 , n440 );
    nor g750 ( n1582 , n1727 , n977 );
    and g751 ( n1315 , n411 , n475 );
    nor g752 ( n1271 , n560 , n341 );
    not g753 ( n1694 , n1205 );
    or g754 ( n441 , n1041 , n579 );
    nor g755 ( n1245 , n579 , n1229 );
    nor g756 ( n1371 , n1102 , n816 );
    not g757 ( n1646 , n1088 );
    nor g758 ( n246 , n539 , n1656 );
    nor g759 ( n376 , n539 , n1548 );
    or g760 ( n308 , n1205 , n1087 );
    nor g761 ( n1156 , n1166 , n1435 );
    not g762 ( n1719 , n258 );
    or g763 ( n1381 , n342 , n1358 );
    and g764 ( n1021 , n184 , n1098 );
    or g765 ( n1303 , n1492 , n579 );
    not g766 ( n339 , n371 );
    not g767 ( n998 , n1083 );
    not g768 ( n489 , n1638 );
    buf g769 ( n40 , n792 );
    nor g770 ( n140 , n323 , n1176 );
    or g771 ( n1585 , n287 , n1107 );
    and g772 ( n409 , n579 , n195 );
    xnor g773 ( n637 , n1515 , n643 );
    or g774 ( n299 , n261 , n409 );
    or g775 ( n1006 , n1785 , n1200 );
    and g776 ( n1578 , n1132 , n735 );
    or g777 ( n1259 , n1170 , n579 );
    not g778 ( n947 , n1512 );
    nor g779 ( n756 , n261 , n269 );
    and g780 ( n905 , n49 , n1786 );
    and g781 ( n1113 , n1146 , n1564 );
    not g782 ( n1795 , n1244 );
    or g783 ( n118 , n186 , n1631 );
    or g784 ( n910 , n627 , n1495 );
    or g785 ( n1558 , n1441 , n1452 );
    or g786 ( n1752 , n483 , n941 );
    not g787 ( n763 , n231 );
    or g788 ( n1070 , n358 , n1310 );
    xnor g789 ( n558 , n526 , n949 );
    nor g790 ( n260 , n1585 , n1545 );
    nor g791 ( n241 , n1745 , n212 );
    nor g792 ( n1499 , n1162 , n141 );
    not g793 ( n490 , n1119 );
    and g794 ( n1501 , n147 , n1382 );
    nor g795 ( n1765 , n228 , n1266 );
    or g796 ( n5 , n1379 , n1617 );
    xnor g797 ( n1583 , n1619 , n1029 );
    and g798 ( n1721 , n1520 , n477 );
    or g799 ( n871 , n1604 , n1114 );
    or g800 ( n4 , n1205 , n1631 );
    and g801 ( n508 , n887 , n504 );
    nor g802 ( n219 , n1395 , n1475 );
    and g803 ( n123 , n471 , n51 );
    or g804 ( n424 , n134 , n77 );
    and g805 ( n1631 , n301 , n1444 );
    xnor g806 ( n1443 , n216 , n10 );
    nor g807 ( n1556 , n560 , n1629 );
    and g808 ( n414 , n238 , n1118 );
    or g809 ( n705 , n794 , n1040 );
    nor g810 ( n843 , n1395 , n782 );
    and g811 ( n1423 , n136 , n34 );
    or g812 ( n1216 , n398 , n1200 );
    nor g813 ( n478 , n44 , n303 );
    nor g814 ( n225 , n307 , n123 );
    and g815 ( n501 , n966 , n614 );
    nor g816 ( n545 , n1544 , n1324 );
    nor g817 ( n93 , n560 , n621 );
    nor g818 ( n739 , n391 , n892 );
    or g819 ( n599 , n1146 , n1483 );
    or g820 ( n1394 , n725 , n1221 );
    and g821 ( n1549 , n708 , n591 );
    and g822 ( n265 , n799 , n1487 );
    or g823 ( n1734 , n1112 , n1712 );
    not g824 ( n106 , n154 );
    nor g825 ( n895 , n1367 , n787 );
    nor g826 ( n449 , n377 , n700 );
    or g827 ( n1222 , n400 , n1593 );
    xnor g828 ( n644 , n927 , n126 );
    nor g829 ( n1764 , n1345 , n1608 );
    xnor g830 ( n35 , n1421 , n736 );
    or g831 ( n289 , n1205 , n487 );
    not g832 ( n1199 , n1645 );
    nor g833 ( n29 , n261 , n1479 );
    buf g834 ( n375 , n84 );
    nor g835 ( n206 , n377 , n1486 );
    or g836 ( n653 , n8 , n285 );
    not g837 ( n1673 , n1229 );
    xnor g838 ( n126 , n47 , n431 );
    or g839 ( n1104 , n896 , n216 );
    or g840 ( n914 , n720 , n268 );
    not g841 ( n1685 , n1089 );
    and g842 ( n963 , n1729 , n591 );
    nor g843 ( n1404 , n44 , n1438 );
    or g844 ( n1322 , n220 , n570 );
    not g845 ( n1069 , n1578 );
    or g846 ( n1593 , n547 , n976 );
    nor g847 ( n158 , n220 , n856 );
    or g848 ( n1434 , n1105 , n1435 );
    nor g849 ( n1239 , n228 , n1060 );
    nor g850 ( n444 , n395 , n600 );
    or g851 ( n1510 , n1732 , n1055 );
    nor g852 ( n736 , n739 , n1052 );
    nor g853 ( n201 , n1575 , n738 );
    xnor g854 ( n1680 , n438 , n1412 );
    or g855 ( n470 , n307 , n370 );
    and g856 ( n454 , n196 , n1455 );
    xnor g857 ( n1293 , n149 , n1668 );
    or g858 ( n466 , n1620 , n1373 );
    or g859 ( n1760 , n1791 , n227 );
    nor g860 ( n1001 , n377 , n1513 );
    xnor g861 ( n896 , n747 , n1039 );
    nor g862 ( n1215 , n261 , n1528 );
    not g863 ( n79 , n601 );
    nor g864 ( n942 , n832 , n617 );
    or g865 ( n1083 , n1295 , n382 );
    nor g866 ( n164 , n261 , n374 );
    not g867 ( n1054 , n760 );
    nor g868 ( n1379 , n1162 , n914 );
    or g869 ( n596 , n1481 , n183 );
    nor g870 ( n1139 , n1162 , n768 );
    or g871 ( n167 , n1366 , n772 );
    or g872 ( n1650 , n1287 , n885 );
    not g873 ( n450 , n1095 );
    or g874 ( n1193 , n1295 , n561 );
    xnor g875 ( n1327 , n1070 , n60 );
    xnor g876 ( n1605 , n1457 , n1752 );
    not g877 ( n1302 , n15 );
    not g878 ( n169 , n1402 );
    nor g879 ( n318 , n767 , n37 );
    nor g880 ( n1335 , n935 , n1278 );
    or g881 ( n203 , n1502 , n498 );
    not g882 ( n1166 , n721 );
    not g883 ( n1114 , n1255 );
    buf g884 ( n1385 , n1326 );
    or g885 ( n548 , n363 , n896 );
    xnor g886 ( n147 , n1308 , n1402 );
    or g887 ( n1324 , n1433 , n641 );
    not g888 ( n1210 , n1633 );
    nor g889 ( n1109 , n904 , n15 );
    or g890 ( n78 , n143 , n629 );
    or g891 ( n314 , n995 , n268 );
    or g892 ( n866 , n1369 , n97 );
    and g893 ( n1645 , n23 , n106 );
    nor g894 ( n125 , n539 , n118 );
    xnor g895 ( n145 , n408 , n1401 );
    or g896 ( n37 , n1754 , n300 );
    or g897 ( n217 , n307 , n1110 );
    nor g898 ( n727 , n39 , n898 );
    or g899 ( n1123 , n620 , n1109 );
    buf g900 ( n1698 , n673 );
    nor g901 ( n104 , n1162 , n991 );
    or g902 ( n131 , n261 , n1325 );
    nor g903 ( n6 , n781 , n504 );
    nor g904 ( n1399 , n573 , n1609 );
    nor g905 ( n256 , n560 , n1760 );
    or g906 ( n1671 , n720 , n227 );
    or g907 ( n1683 , n1205 , n1710 );
    not g908 ( n188 , n1660 );
    or g909 ( n1212 , n821 , n227 );
    or g910 ( n1359 , n913 , n1728 );
    and g911 ( n1636 , n538 , n1507 );
    nor g912 ( n1197 , n1612 , n1206 );
    nor g913 ( n683 , n57 , n306 );
    nor g914 ( n440 , n228 , n1782 );
    or g915 ( n1414 , n790 , n1450 );
    not g916 ( n402 , n1471 );
    or g917 ( n1103 , n1336 , n1230 );
    not g918 ( n1075 , n1361 );
    or g919 ( n877 , n1072 , n1200 );
    or g920 ( n852 , n1146 , n555 );
    or g921 ( n968 , n186 , n1495 );
    or g922 ( n638 , n1147 , n1405 );
    not g923 ( n832 , n1227 );
    and g924 ( n978 , n1235 , n87 );
    and g925 ( n1310 , n708 , n439 );
    not g926 ( n1375 , n128 );
    or g927 ( n1240 , n1742 , n612 );
    or g928 ( n769 , n1105 , n1660 );
    or g929 ( n928 , n1678 , n443 );
    nor g930 ( n8 , n228 , n742 );
    not g931 ( n1308 , n685 );
    nor g932 ( n535 , n395 , n807 );
    xnor g933 ( n1038 , n1228 , n580 );
    or g934 ( n274 , n275 , n248 );
    not g935 ( n995 , n384 );
    not g936 ( n1170 , n1740 );
    xnor g937 ( n404 , n761 , n380 );
    or g938 ( n1330 , n1789 , n1651 );
    xnor g939 ( n804 , n808 , n1470 );
    or g940 ( n1777 , n1726 , n1275 );
    not g941 ( n645 , n55 );
    or g942 ( n1453 , n1146 , n82 );
    nor g943 ( n480 , n378 , n230 );
    or g944 ( n392 , n428 , n854 );
    or g945 ( n99 , n716 , n362 );
    or g946 ( n1340 , n41 , n579 );
    nor g947 ( n86 , n832 , n1515 );
    nor g948 ( n749 , n495 , n1381 );
    or g949 ( n423 , n1610 , n227 );
    nor g950 ( n445 , n1162 , n775 );
    or g951 ( n1478 , n1178 , n227 );
    not g952 ( n689 , n678 );
    nor g953 ( n1514 , n1172 , n1227 );
    not g954 ( n523 , n319 );
    or g955 ( n233 , n1351 , n939 );
    not g956 ( n1419 , n530 );
    nor g957 ( n292 , n1781 , n1778 );
    and g958 ( n1476 , n88 , n500 );
    not g959 ( n809 , n10 );
    or g960 ( n355 , n1585 , n1004 );
    or g961 ( n597 , n197 , n227 );
    not g962 ( n752 , n719 );
    or g963 ( n1666 , n1724 , n446 );
    or g964 ( n367 , n1204 , n1643 );
    or g965 ( n1672 , n671 , n171 );
    or g966 ( n1057 , n1624 , n579 );
    not g967 ( n1162 , n377 );
    nor g968 ( n1482 , n44 , n965 );
    xor g969 ( n547 , n1203 , n1677 );
    or g970 ( n1418 , n1699 , n21 );
    or g971 ( n1225 , n266 , n278 );
    not g972 ( n1618 , n1238 );
    nor g973 ( n1352 , n966 , n714 );
    or g974 ( n156 , n1253 , n579 );
    or g975 ( n502 , n494 , n1315 );
    nor g976 ( n262 , n220 , n665 );
    not g977 ( n200 , n714 );
    or g978 ( n1523 , n1241 , n1236 );
    or g979 ( n329 , n571 , n170 );
    nor g980 ( n1484 , n134 , n807 );
    or g981 ( n1424 , n1126 , n227 );
    xnor g982 ( n1489 , n1293 , n1461 );
    or g983 ( n122 , n458 , n1289 );
    or g984 ( n608 , n658 , n1200 );
    or g985 ( n294 , n659 , n1787 );
    or g986 ( n419 , n284 , n948 );
    nor g987 ( n718 , n1395 , n598 );
    nor g988 ( n1243 , n134 , n591 );
    or g989 ( n1214 , n1205 , n75 );
    nor g990 ( n980 , n200 , n617 );
    not g991 ( n1395 , n228 );
    or g992 ( n1266 , n1205 , n905 );
    nor g993 ( n1117 , n1162 , n217 );
    and g994 ( n584 , n560 , n753 );
    not g995 ( n59 , n901 );
    not g996 ( n825 , n88 );
    xnor g997 ( n927 , n1443 , n576 );
    not g998 ( n1488 , n386 );
    nor g999 ( n858 , n1198 , n1717 );
    nor g1000 ( n1115 , n378 , n660 );
    and g1001 ( n1231 , n155 , n1108 );
    nor g1002 ( n1658 , n261 , n1267 );
    or g1003 ( n1080 , n1615 , n579 );
    or g1004 ( n634 , n825 , n1104 );
    or g1005 ( n1076 , n957 , n1694 );
    and g1006 ( n859 , n1437 , n1501 );
    or g1007 ( n569 , n1368 , n663 );
    xnor g1008 ( n994 , n1605 , n1038 );
    not g1009 ( n151 , n1476 );
    nor g1010 ( n797 , n1100 , n1431 );
    or g1011 ( n258 , n1026 , n434 );
    or g1012 ( n991 , n307 , n469 );
    not g1013 ( n658 , n270 );
    and g1014 ( n1151 , n872 , n367 );
    not g1015 ( n1122 , n190 );
    xnor g1016 ( n1555 , n1236 , n286 );
    nor g1017 ( n1526 , n380 , n1519 );
    not g1018 ( n1774 , n1501 );
    nor g1019 ( n27 , n200 , n1043 );
    xnor g1020 ( n988 , n703 , n397 );
    not g1021 ( n821 , n1150 );
    not g1022 ( n185 , n743 );
    not g1023 ( n1574 , n119 );
    or g1024 ( n1465 , n61 , n1661 );
    or g1025 ( n323 , n433 , n619 );
    and g1026 ( n358 , n1408 , n504 );
    nor g1027 ( n359 , n188 , n504 );
    or g1028 ( n1071 , n1432 , n268 );
    or g1029 ( n528 , n1139 , n970 );
    or g1030 ( n1091 , n1100 , n351 );
    and g1031 ( n529 , n1632 , n504 );
    not g1032 ( n1662 , n600 );
    nor g1033 ( n1263 , n1484 , n839 );
    or g1034 ( n189 , n865 , n1694 );
    or g1035 ( n972 , n1000 , n1001 );
    xnor g1036 ( n517 , n686 , n975 );
    not g1037 ( n252 , n948 );
    or g1038 ( n17 , n1105 , n1238 );
    or g1039 ( n1098 , n1575 , n1449 );
    nor g1040 ( n212 , n261 , n950 );
    nor g1041 ( n788 , n1034 , n705 );
    nor g1042 ( n612 , n1498 , n721 );
    or g1043 ( n81 , n1125 , n886 );
    and g1044 ( n379 , n1613 , n172 );
    nor g1045 ( n1262 , n560 , n875 );
    not g1046 ( n630 , n1575 );
    or g1047 ( n1659 , n953 , n1696 );
    not g1048 ( n28 , n1535 );
    nor g1049 ( n733 , n1676 , n1662 );
    and g1050 ( n1780 , n84 , n1058 );
    nor g1051 ( n36 , n587 , n208 );
    not g1052 ( n849 , n516 );
    not g1053 ( n311 , n953 );
    nor g1054 ( n108 , n1162 , n1496 );
    not g1055 ( n1002 , n368 );
    nor g1056 ( n343 , n1553 , n1519 );
    or g1057 ( n981 , n1384 , n634 );
    or g1058 ( n1486 , n307 , n487 );
    xnor g1059 ( n154 , n717 , n326 );
    or g1060 ( n83 , n1247 , n505 );
    xnor g1061 ( n1284 , n1024 , n863 );
    nor g1062 ( n926 , n579 , n274 );
    nor g1063 ( n1608 , n261 , n1311 );
    not g1064 ( n1689 , n754 );
    not g1065 ( n1136 , n1788 );
    nor g1066 ( n1317 , n1447 , n322 );
    and g1067 ( n1628 , n1225 , n1581 );
    and g1068 ( n1495 , n852 , n1627 );
    and g1069 ( n648 , n1396 , n504 );
    not g1070 ( n434 , n717 );
    not g1071 ( n1686 , n33 );
    or g1072 ( n1472 , n710 , n600 );
    or g1073 ( n854 , n996 , n534 );
    xnor g1074 ( n1643 , n804 , n666 );
    or g1075 ( n1313 , n1551 , n1376 );
    or g1076 ( n1377 , n553 , n730 );
    or g1077 ( n1102 , n554 , n199 );
    xnor g1078 ( n1445 , n747 , n1579 );
    or g1079 ( n1531 , n1016 , n267 );
    or g1080 ( n657 , n924 , n579 );
    xnor g1081 ( n1134 , n818 , n291 );
    or g1082 ( n1456 , n1522 , n268 );
    or g1083 ( n1730 , n1264 , n227 );
    xnor g1084 ( n328 , n642 , n557 );
    nor g1085 ( n1455 , n29 , n71 );
    nor g1086 ( n939 , n378 , n1265 );
    or g1087 ( n415 , n979 , n784 );
    nor g1088 ( n1559 , n134 , n504 );
    nor g1089 ( n883 , n44 , n891 );
    xnor g1090 ( n1536 , n1585 , n291 );
    not g1091 ( n1624 , n157 );
    or g1092 ( n1073 , n1205 , n1110 );
    buf g1093 ( n793 , n544 );
    and g1094 ( n589 , n1707 , n600 );
    buf g1095 ( n860 , n623 );
    and g1096 ( n583 , n706 , n1597 );
    nor g1097 ( n492 , n228 , n1246 );
    xnor g1098 ( n863 , n1238 , n1498 );
    or g1099 ( n1089 , n1433 , n1152 );
    not g1100 ( n1289 , n216 );
    and g1101 ( n174 , n1106 , n703 );
    not g1102 ( n1573 , n39 );
    or g1103 ( n1479 , n579 , n1638 );
    and g1104 ( n487 , n594 , n1158 );
    xnor g1105 ( n778 , n966 , n946 );
    and g1106 ( n1108 , n1532 , n392 );
    or g1107 ( n1137 , n781 , n614 );
    xnor g1108 ( n1249 , n1195 , n1415 );
    or g1109 ( n1388 , n169 , n1308 );
    or g1110 ( n1138 , n486 , n579 );
    xnor g1111 ( n1025 , n996 , n1788 );
    or g1112 ( n662 , n1406 , n36 );
    or g1113 ( n113 , n627 , n454 );
    or g1114 ( n455 , n1171 , n1535 );
    nor g1115 ( n916 , n485 , n412 );
    or g1116 ( n1398 , n630 , n1547 );
    or g1117 ( n102 , n226 , n1099 );
    or g1118 ( n305 , n186 , n454 );
    xnor g1119 ( n663 , n896 , n1183 );
    nor g1120 ( n695 , n1395 , n805 );
    nor g1121 ( n771 , n1660 , n1227 );
    xnor g1122 ( n761 , n637 , n670 );
    not g1123 ( n1332 , n1737 );
    nor g1124 ( n420 , n261 , n1012 );
    nor g1125 ( n1687 , n1650 , n1652 );
    or g1126 ( n413 , n528 , n1738 );
    xnor g1127 ( n47 , n1777 , n363 );
    or g1128 ( n1165 , n1662 , n1568 );
    or g1129 ( n1483 , n1372 , n579 );
    not g1130 ( n1334 , n1743 );
    or g1131 ( n834 , n785 , n253 );
    nor g1132 ( n1331 , n817 , n182 );
    nor g1133 ( n116 , n378 , n1260 );
    nor g1134 ( n1562 , n539 , n1124 );
    nor g1135 ( n1367 , n44 , n521 );
    not g1136 ( n451 , n1219 );
    or g1137 ( n1467 , n496 , n1387 );
    nor g1138 ( n876 , n539 , n985 );
    nor g1139 ( n1767 , n1395 , n1430 );
    or g1140 ( n901 , n681 , n1559 );
    and g1141 ( n1507 , n1788 , n485 );
    nor g1142 ( n1727 , n1243 , n958 );
    or g1143 ( n1019 , n853 , n1312 );
    or g1144 ( n117 , n79 , n537 );
    nor g1145 ( n1079 , n1115 , n1606 );
    not g1146 ( n1356 , n534 );
    or g1147 ( n687 , n146 , n89 );
    or g1148 ( n1187 , n1205 , n1314 );
    nor g1149 ( n940 , n1626 , n1777 );
    or g1150 ( n1586 , n186 , n1346 );
    or g1151 ( n953 , n992 , n549 );
    nor g1152 ( n135 , n1276 , n420 );
    nor g1153 ( n692 , n1162 , n1008 );
    nor g1154 ( n1078 , n1205 , n123 );
    or g1155 ( n954 , n897 , n1616 );
    xnor g1156 ( n1565 , n1236 , n205 );
    or g1157 ( n892 , n345 , n1007 );
    not g1158 ( n1275 , n1571 );
    or g1159 ( n573 , n406 , n1538 );
    nor g1160 ( n609 , n228 , n304 );
    nor g1161 ( n170 , n0 , n766 );
    not g1162 ( n1374 , n1010 );
    nor g1163 ( n861 , n237 , n1658 );
    or g1164 ( n1256 , n205 , n1360 );
    or g1165 ( n686 , n648 , n202 );
    or g1166 ( n639 , n1295 , n1776 );
    xnor g1167 ( n581 , n1702 , n502 );
    not g1168 ( n1169 , n179 );
    and g1169 ( n1062 , n378 , n45 );
    nor g1170 ( n665 , n1394 , n1666 );
    nor g1171 ( n772 , n296 , n1489 );
    or g1172 ( n1602 , n582 , n93 );
    nor g1173 ( n559 , n1645 , n1164 );
    nor g1174 ( n1354 , n1016 , n1516 );
    nor g1175 ( n1748 , n1238 , n714 );
    not g1176 ( n1626 , n634 );
    not g1177 ( n422 , n132 );
    and g1178 ( n1027 , n607 , n135 );
    or g1179 ( n313 , n1151 , n1705 );
    or g1180 ( n1111 , n627 , n882 );
    not g1181 ( n296 , n1669 );
    or g1182 ( n180 , n627 , n1027 );
    not g1183 ( n1020 , n1181 );
    xnor g1184 ( n1506 , n481 , n1094 );
    or g1185 ( n874 , n490 , n268 );
    nor g1186 ( n1733 , n220 , n1634 );
    or g1187 ( n247 , n627 , n487 );
    or g1188 ( n1267 , n1295 , n689 );
    or g1189 ( n1746 , n1295 , n1049 );
    not g1190 ( n427 , n1680 );
    xnor g1191 ( n624 , n1470 , n1795 );
    nor g1192 ( n1701 , n703 , n243 );
    and g1193 ( n800 , n1192 , n1566 );
    nor g1194 ( n839 , n1172 , n714 );
    or g1195 ( n983 , n1689 , n227 );
    not g1196 ( n1146 , n261 );
    xnor g1197 ( n1461 , n534 , n919 );
    or g1198 ( n1732 , n688 , n42 );
    nor g1199 ( n1052 , n1391 , n1009 );
    not g1200 ( n613 , n639 );
    not g1201 ( n50 , n353 );
    nor g1202 ( n982 , n539 , n983 );
    or g1203 ( n341 , n186 , n168 );
    or g1204 ( n640 , n1128 , n227 );
    nor g1205 ( n273 , n1342 , n500 );
    nor g1206 ( n46 , n699 , n646 );
    and g1207 ( n757 , n238 , n1165 );
    or g1208 ( n243 , n1437 , n397 );
    or g1209 ( n603 , n1133 , n755 );
    nor g1210 ( n1715 , n261 , n109 );
    not g1211 ( n957 , n1675 );
    and g1212 ( n275 , n697 , n506 );
    or g1213 ( n590 , n401 , n978 );
    not g1214 ( n720 , n564 );
    nor g1215 ( n1444 , n527 , n1715 );
    and g1216 ( n934 , n1146 , n1082 );
    and g1217 ( n276 , n385 , n1004 );
    or g1218 ( n1490 , n1326 , n650 );
    nor g1219 ( n425 , n748 , n600 );
    or g1220 ( n869 , n30 , n883 );
    nor g1221 ( n567 , n220 , n1687 );
    nor g1222 ( n582 , n539 , n423 );
    nor g1223 ( n977 , n697 , n1263 );
    nor g1224 ( n615 , n377 , n1068 );
    or g1225 ( n1230 , n263 , n1621 );
    or g1226 ( n965 , n802 , n1200 );
    nor g1227 ( n986 , n188 , n591 );
    and g1228 ( n610 , n966 , n1118 );
    nor g1229 ( n463 , n438 , n825 );
    and g1230 ( n1346 , n1090 , n1056 );
    and g1231 ( n1004 , n1173 , n682 );
    nor g1232 ( n738 , n1023 , n166 );
    not g1233 ( n1189 , n586 );
    and g1234 ( n791 , n757 , n1668 );
    and g1235 ( n1373 , n331 , n989 );
    nor g1236 ( n51 , n934 , n932 );
    and g1237 ( n1564 , n679 , n1667 );
    or g1238 ( n1387 , n1069 , n1595 );
    not g1239 ( n1610 , n297 );
    or g1240 ( n730 , n1458 , n827 );
    not g1241 ( n1595 , n870 );
    nor g1242 ( n677 , n514 , n1204 );
    and g1243 ( n87 , n810 , n538 );
    nor g1244 ( n1493 , n1395 , n1066 );
    not g1245 ( n867 , n1643 );
    nor g1246 ( n222 , n220 , n577 );
    or g1247 ( n322 , n429 , n1179 );
    or g1248 ( n1342 , n1685 , n250 );
    xnor g1249 ( n576 , n88 , n531 );
    or g1250 ( n69 , n1420 , n1209 );
    or g1251 ( n411 , n853 , n614 );
    and g1252 ( n1705 , n1175 , n812 );
    or g1253 ( n1045 , n523 , n614 );
    or g1254 ( n789 , n1021 , n497 );
    not g1255 ( n462 , n387 );
    or g1256 ( n172 , n1385 , n1273 );
    nor g1257 ( n1459 , n377 , n1252 );
    nor g1258 ( n631 , n1681 , n38 );
    or g1259 ( n1709 , n702 , n1694 );
    or g1260 ( n362 , n1789 , n1156 );
    or g1261 ( n969 , n774 , n1200 );
    nor g1262 ( n1581 , n579 , n1731 );
    nor g1263 ( n1704 , n1498 , n714 );
    nor g1264 ( n911 , n560 , n1735 );
    xnor g1265 ( n1664 , n1141 , n110 );
    or g1266 ( n777 , n847 , n59 );
    and g1267 ( n171 , n1333 , n1577 );
    or g1268 ( n915 , n399 , n928 );
    not g1269 ( n1464 , n389 );
    and g1270 ( n1545 , n258 , n1199 );
    nor g1271 ( n1502 , n539 , n640 );
    or g1272 ( n951 , n631 , n922 );
    or g1273 ( n1005 , n332 , n1200 );
    not g1274 ( n1014 , n1145 );
    nor g1275 ( n837 , n378 , n247 );
    or g1276 ( n851 , n105 , n461 );
    or g1277 ( n806 , n518 , n820 );
    not g1278 ( n960 , n271 );
    nor g1279 ( n1588 , n1366 , n690 );
    xnor g1280 ( n0 , n751 , n1468 );
    or g1281 ( n352 , n1307 , n1694 );
    or g1282 ( n1229 , n921 , n1306 );
    or g1283 ( n1163 , n1527 , n117 );
    not g1284 ( n844 , n1353 );
    and g1285 ( n870 , n393 , n866 );
    nor g1286 ( n315 , n220 , n788 );
    and g1287 ( n964 , n1392 , n1197 );
    or g1288 ( n729 , n186 , n1087 );
    not g1289 ( n244 , n1473 );
    and g1290 ( n1255 , n460 , n418 );
    xnor g1291 ( n1142 , n1127 , n871 );
    not g1292 ( n822 , n328 );
    or g1293 ( n1173 , n284 , n392 );
    or g1294 ( n833 , n1375 , n1694 );
    not g1295 ( n1566 , n276 );
    or g1296 ( n196 , n1146 , n657 );
    not g1297 ( n1360 , n1160 );
    nor g1298 ( n593 , n986 , n1592 );
    xnor g1299 ( n438 , n550 , n1135 );
    not g1300 ( n1372 , n999 );
    not g1301 ( n1211 , n274 );
    or g1302 ( n1623 , n159 , n234 );
    or g1303 ( n467 , n1507 , n412 );
    or g1304 ( n76 , n366 , n1153 );
    or g1305 ( n349 , n277 , n246 );
    or g1306 ( n563 , n1075 , n579 );
    nor g1307 ( n1050 , n220 , n459 );
    not g1308 ( n1298 , n779 );
    not g1309 ( n1031 , n686 );
    nor g1310 ( n1276 , n261 , n372 );
    or g1311 ( n635 , n1734 , n923 );
    or g1312 ( n709 , n148 , n161 );
    nor g1313 ( n1606 , n44 , n556 );
    and g1314 ( n1383 , n1518 , n591 );
    or g1315 ( n938 , n124 , n543 );
    or g1316 ( n997 , n615 , n973 );
    nor g1317 ( n1349 , n560 , n595 );
    xnor g1318 ( n405 , n1762 , n16 );
    nor g1319 ( n1305 , n377 , n152 );
    or g1320 ( n1092 , n1146 , n162 );
    or g1321 ( n622 , n579 , n244 );
    and g1322 ( n1269 , n1411 , n1167 );
    not g1323 ( n193 , n937 );
    nor g1324 ( n96 , n539 , n836 );
    and g1325 ( n625 , n1146 , n1245 );
    xnor g1326 ( n88 , n549 , n1100 );
    nor g1327 ( n1678 , n1681 , n532 );
    not g1328 ( n1178 , n239 );
    buf g1329 ( n1233 , n1044 );
    nor g1330 ( n1542 , n832 , n1518 );
    xnor g1331 ( n1792 , n302 , n808 );
    nor g1332 ( n1771 , n44 , n204 );
    nor g1333 ( n1587 , n220 , n1679 );
    nor g1334 ( n1500 , n539 , n58 );
    nor g1335 ( n1364 , n1146 , n422 );
    and g1336 ( n370 , n98 , n683 );
    or g1337 ( n1392 , n1146 , n1080 );
    not g1338 ( n1791 , n955 );
    not g1339 ( n111 , n1756 );
    or g1340 ( n412 , n810 , n696 );
    or g1341 ( n1494 , n1295 , n907 );
    or g1342 ( n1589 , n1718 , n586 );
    xnor g1343 ( n711 , n1359 , n1755 );
    nor g1344 ( n740 , n1339 , n1300 );
    nor g1345 ( n989 , n39 , n980 );
    or g1346 ( n1413 , n849 , n878 );
    and g1347 ( n1232 , n1366 , n405 );
    or g1348 ( n62 , n1673 , n1736 );
    nor g1349 ( n641 , n1498 , n1227 );
    or g1350 ( n1644 , n1334 , n1200 );
    or g1351 ( n1759 , n224 , n1117 );
    and g1352 ( n1710 , n599 , n138 );
    buf g1353 ( n1378 , n84 );
    and g1354 ( n1198 , n1146 , n1120 );
    nor g1355 ( n1635 , n1618 , n504 );
    xnor g1356 ( n15 , n1134 , n1583 );
    not g1357 ( n696 , n854 );
    xnor g1358 ( n1776 , n938 , n684 );
    nor g1359 ( n54 , n1713 , n504 );
    and g1360 ( n737 , n959 , n513 );
    not g1361 ( n1140 , n1568 );
    or g1362 ( n58 , n1169 , n227 );
    and g1363 ( n334 , n1272 , n559 );
    not g1364 ( n146 , n1025 );
    or g1365 ( n1176 , n492 , n1493 );
    not g1366 ( n766 , n1283 );
    or g1367 ( n153 , n658 , n1694 );
    xnor g1368 ( n751 , n147 , n531 );
    buf g1369 ( n765 , n1044 );
    and g1370 ( n1551 , n39 , n1418 );
    nor g1371 ( n1712 , n377 , n312 );
    and g1372 ( n904 , n419 , n1004 );
    or g1373 ( n1278 , n992 , n1474 );
    nor g1374 ( n1067 , n853 , n600 );
    or g1375 ( n604 , n1105 , n1729 );
    or g1376 ( n142 , n627 , n1314 );
    or g1377 ( n1592 , n630 , n771 );
    nor g1378 ( n1590 , n501 , n1352 );
    and g1379 ( n105 , n1238 , n1288 );
    nor g1380 ( n755 , n1281 , n451 );
    or g1381 ( n1416 , n481 , n231 );
    or g1382 ( n976 , n1511 , n320 );
    nor g1383 ( n1577 , n60 , n707 );
    or g1384 ( n1384 , n438 , n481 );
    or g1385 ( n514 , n1327 , n1750 );
    not g1386 ( n924 , n1753 );
    or g1387 ( n471 , n1146 , n1138 );
    or g1388 ( n284 , n149 , n1130 );
    nor g1389 ( n1084 , n1395 , n189 );
    xnor g1390 ( n1192 , n154 , n1695 );
    xnor g1391 ( n16 , n1142 , n360 );
    or g1392 ( n836 , n952 , n227 );
    or g1393 ( n553 , n90 , n1274 );
    and g1394 ( n10 , n1630 , n255 );
    or g1395 ( n556 , n627 , n469 );
    buf g1396 ( n1682 , n130 );
    and g1397 ( n1258 , n1146 , n926 );
    and g1398 ( n1706 , n1077 , n1164 );
    and g1399 ( n497 , n1442 , n524 );
    or g1400 ( n1638 , n447 , n86 );
    buf g1401 ( n776 , n1613 );
    nor g1402 ( n619 , n228 , n1076 );
    or g1403 ( n732 , n1146 , n1688 );
    nor g1404 ( n1505 , n1220 , n1185 );
    and g1405 ( n882 , n1092 , n1739 );
    nor g1406 ( n221 , n832 , n1729 );
    not g1407 ( n1072 , n1362 );
    xnor g1408 ( n949 , n397 , n826 );
    or g1409 ( n1068 , n307 , n1027 );
    not g1410 ( n396 , n302 );
    not g1411 ( n835 , n1108 );
    and g1412 ( n1796 , n703 , n1257 );
    not g1413 ( n1422 , n1059 );
    nor g1414 ( n1074 , n378 , n910 );
    not g1415 ( n408 , n1165 );
    not g1416 ( n479 , n636 );
    nor g1417 ( n1009 , n32 , n750 );
    nor g1418 ( n70 , n464 , n1558 );
    and g1419 ( n921 , n1039 , n1240 );
    not g1420 ( n197 , n1207 );
    or g1421 ( n1738 , n31 , n1499 );
    not g1422 ( n764 , n236 );
    or g1423 ( n1213 , n1504 , n603 );
    or g1424 ( n356 , n238 , n77 );
    nor g1425 ( n264 , n1465 , n1149 );
    not g1426 ( n1196 , n497 );
    or g1427 ( n1159 , n515 , n316 );
    or g1428 ( n1563 , n627 , n1087 );
    and g1429 ( n543 , n1366 , n1123 );
    or g1430 ( n272 , n811 , n1261 );
    nor g1431 ( n410 , n1135 , n1323 );
    nor g1432 ( n1251 , n1039 , n831 );
    or g1433 ( n442 , n1332 , n489 );
    not g1434 ( n1312 , n77 );
    nor g1435 ( n477 , n909 , n419 );
    xor g1436 ( n538 , n1228 , n1016 );
    xor g1437 ( n149 , n408 , n238 );
    not g1438 ( n390 , n1489 );
    or g1439 ( n985 , n186 , n1110 );
    nor g1440 ( n1325 , n1295 , n1776 );
    not g1441 ( n1703 , n1454 );
    not g1442 ( n702 , n7 );
    or g1443 ( n496 , n1680 , n1059 );
    nor g1444 ( n80 , n568 , n416 );
    or g1445 ( n598 , n802 , n1694 );
    or g1446 ( n1018 , n1432 , n227 );
    or g1447 ( n1242 , n627 , n1346 );
    or g1448 ( n680 , n627 , n1710 );
    or g1449 ( n568 , n1393 , n1239 );
    and g1450 ( n1382 , n463 , n1013 );
    or g1451 ( n796 , n1295 , n1720 );
    nor g1452 ( n682 , n474 , n218 );
    xor g1453 ( n1511 , n404 , n1035 );
    nor g1454 ( n1462 , n220 , n318 );
    or g1455 ( n923 , n449 , n104 );
    or g1456 ( n1277 , n627 , n370 );
    or g1457 ( n1513 , n694 , n268 );
    nor g1458 ( n1223 , n330 , n1704 );
    or g1459 ( n304 , n1785 , n1694 );
    xnor g1460 ( n1203 , n1647 , n1048 );
    nor g1461 ( n306 , n261 , n1546 );
    not g1462 ( n694 , n1177 );
    and g1463 ( n55 , n752 , n234 );
    not g1464 ( n820 , n628 );
    xnor g1465 ( n868 , n1172 , n1553 );
    or g1466 ( n18 , n1201 , n1157 );
    nor g1467 ( n139 , n1084 , n1517 );
    or g1468 ( n521 , n865 , n1200 );
    nor g1469 ( n163 , n832 , n319 );
    or g1470 ( n310 , n186 , n964 );
    not g1471 ( n900 , n1655 );
    or g1472 ( n908 , n1610 , n268 );
    or g1473 ( n580 , n1015 , n1067 );
    nor g1474 ( n1133 , n1681 , n1646 );
    xnor g1475 ( n510 , n534 , n1237 );
    or g1476 ( n1688 , n1122 , n579 );
    nor g1477 ( n1554 , n1395 , n1625 );
    xnor g1478 ( n642 , n818 , n1766 );
    or g1479 ( n717 , n744 , n1321 );
    nor g1480 ( n484 , n1402 , n1747 );
    buf g1481 ( n1326 , n117 );
    nor g1482 ( n1208 , n1553 , n1227 );
    nor g1483 ( n21 , n617 , n721 );
    xnor g1484 ( n1024 , n617 , n1674 );
    or g1485 ( n621 , n995 , n227 );
    or g1486 ( n460 , n149 , n392 );
    or g1487 ( n381 , n803 , n52 );
    or g1488 ( n1758 , n579 , n1737 );
    or g1489 ( n1028 , n579 , n936 );
    nor g1490 ( n688 , n539 , n899 );
    nor g1491 ( n731 , n1172 , n721 );
    not g1492 ( n1789 , n1016 );
    xnor g1493 ( n1226 , n507 , n1406 );
    nor g1494 ( n893 , n228 , n85 );
    buf g1495 ( n1657 , n389 );
    nor g1496 ( n1653 , n44 , n680 );
    nor g1497 ( n1405 , n946 , n1227 );
    and g1498 ( n1477 , n1729 , n1288 );
    not g1499 ( n472 , n1553 );
    or g1500 ( n1714 , n307 , n168 );
    nor g1501 ( n897 , n44 , n1216 );
    not g1502 ( n952 , n187 );
    not g1503 ( n1105 , n1519 );
    not g1504 ( n1126 , n1540 );
    nor g1505 ( n1015 , n112 , n1662 );
    nor g1506 ( n1621 , n1166 , n1043 );
    or g1507 ( n198 , n1254 , n902 );
    buf g1508 ( n967 , n357 );
    nor g1509 ( n1120 , n579 , n1313 );
    or g1510 ( n473 , n1767 , n893 );
    not g1511 ( n159 , n826 );
    and g1512 ( n1106 , n1575 , n652 );
    or g1513 ( n1201 , n773 , n256 );
    nor g1514 ( n1101 , n539 , n1586 );
    buf g1515 ( n611 , n84 );
    or g1516 ( n279 , n1205 , n882 );
    or g1517 ( n1380 , n186 , n882 );
    or g1518 ( n1579 , n383 , n1635 );
    not g1519 ( n846 , n1182 );
    not g1520 ( n1522 , n565 );
    or g1521 ( n762 , n1271 , n1101 );
    and g1522 ( n616 , n894 , n600 );
    or g1523 ( n1450 , n1796 , n677 );
    or g1524 ( n1132 , n1257 , n806 );
    nor g1525 ( n1195 , n1342 , n1013 );
    not g1526 ( n781 , n1729 );
    not g1527 ( n1749 , n507 );
    nor g1528 ( n1400 , n579 , n783 );
    or g1529 ( n1640 , n579 , n1218 );
    or g1530 ( n550 , n508 , n6 );
    and g1531 ( n1569 , n1659 , n1416 );
    not g1532 ( n1218 , n1423 );
    not g1533 ( n1779 , n1368 );
    not g1534 ( n829 , n1021 );
    nor g1535 ( n1725 , n377 , n115 );
    or g1536 ( n1652 , n837 , n1653 );
    nor g1537 ( n13 , n697 , n133 );
    and g1538 ( n973 , n377 , n225 );
    or g1539 ( n97 , n1701 , n628 );
    and g1540 ( n690 , n1004 , n328 );
    or g1541 ( n1609 , n1319 , n1554 );
    not g1542 ( n614 , n807 );
    or g1543 ( n723 , n1713 , n77 );
    and g1544 ( n209 , n1016 , n1228 );
    nor g1545 ( n1448 , n614 , n238 );
    or g1546 ( n312 , n111 , n268 );
    nor g1547 ( n1538 , n228 , n352 );
    not g1548 ( n992 , n1100 );
    not g1549 ( n458 , n363 );
    or g1550 ( n293 , n1026 , n572 );
    nor g1551 ( n554 , n44 , n175 );
    nor g1552 ( n1580 , n395 , n591 );
    nor g1553 ( n1393 , n1395 , n1304 );
    not g1554 ( n1194 , n520 );
    xnor g1555 ( n14 , n717 , n507 );
    and g1556 ( n706 , n981 , n1204 );
    nor g1557 ( n815 , n377 , n3 );
    xnor g1558 ( n1329 , n795 , n294 );
    or g1559 ( n660 , n627 , n905 );
    or g1560 ( n1344 , n1665 , n1639 );
    xnor g1561 ( n919 , n428 , n1255 );
    or g1562 ( n931 , n1295 , n510 );
    nor g1563 ( n1516 , n535 , n925 );
    or g1564 ( n1055 , n1365 , n125 );
    nor g1565 ( n1525 , n539 , n729 );
    and g1566 ( n287 , n971 , n600 );
    xnor g1567 ( n26 , n145 , n994 );
    not g1568 ( n847 , n697 );
    nor g1569 ( n1560 , n44 , n1242 );
    or g1570 ( n141 , n307 , n456 );
    not g1571 ( n394 , n1359 );
    nor g1572 ( n11 , n539 , n1212 );
    nor g1573 ( n1155 , n261 , n1640 );
    or g1574 ( n162 , n846 , n579 );
    not g1575 ( n1668 , n1130 );
    nor g1576 ( n1781 , n261 , n1751 );
    and g1577 ( n245 , n1613 , n1213 );
    and g1578 ( n338 , n504 , n64 );
    nor g1579 ( n1612 , n261 , n333 );
    xnor g1580 ( n1783 , n438 , n1696 );
    not g1581 ( n1347 , n783 );
    and g1582 ( n1535 , n1769 , n662 );
    or g1583 ( n1751 , n579 , n829 );
    and g1584 ( n1336 , n1043 , n1288 );
    or g1585 ( n303 , n627 , n1631 );
    nor g1586 ( n1300 , n819 , n329 );
    or g1587 ( n178 , n307 , n882 );
    or g1588 ( n1576 , n900 , n268 );
    or g1589 ( n282 , n844 , n1200 );
    nor g1590 ( n864 , n1162 , n1456 );
    not g1591 ( n748 , n380 );
    or g1592 ( n684 , n114 , n1232 );
    xnor g1593 ( n889 , n1793 , n1397 );
    and g1594 ( n913 , n917 , n504 );
    nor g1595 ( n540 , n347 , n127 );
    or g1596 ( n1030 , n746 , n584 );
    or g1597 ( n775 , n1264 , n268 );
    or g1598 ( n742 , n1205 , n1495 );
    nor g1599 ( n1742 , n1713 , n1288 );
    nor g1600 ( n1351 , n44 , n633 );
    xnor g1601 ( n1470 , n703 , n396 );
    or g1602 ( n336 , n186 , n456 );
    not g1603 ( n1432 , n488 );
    or g1604 ( n1487 , n1135 , n1168 );
    or g1605 ( n1409 , n537 , n1427 );
    xnor g1606 ( n1368 , n216 , n1279 );
    or g1607 ( n979 , n632 , n678 );
    nor g1608 ( n1754 , n228 , n1693 );
    not g1609 ( n220 , n1534 );
    or g1610 ( n881 , n627 , n456 );
    xnor g1611 ( n525 , n901 , n1359 );
    nand g1612 ( n1411 , n1357 , n1649 );
    xnor g1613 ( n353 , n468 , n207 );
    and g1614 ( n248 , n424 , n13 );
    nor g1615 ( n71 , n261 , n734 );
    not g1616 ( n1241 , n205 );
    nor g1617 ( n433 , n1395 , n1296 );
    nor g1618 ( n1702 , n759 , n1354 );
    or g1619 ( n1320 , n116 , n1560 );
endmodule
