//
// Conformal-LEC Version 15.20-d227 ( 10-Mar-2016) ( 64 bit executable)
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , PI_DFF_B_reg_Q , n9 , PI_DFF_rd_reg_Q , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , PI_DFF_wr_reg_Q , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , PI_PI_reset , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , PI_DFF_state_reg_Q , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , PI_PI_clock , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 , n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , PI_DFF_B_reg_Q , n9 , PI_DFF_rd_reg_Q , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , PI_DFF_wr_reg_Q , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , PI_PI_reset , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , PI_DFF_state_reg_Q , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 , n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 , n216 , n217 , n218 , n219 , n220 , n221 , n222 , n223 , n224 , n225 , n226 , n227 , n228 , n229 , n230 , n231 , n232 , n233 , PI_PI_clock , n234 , n235 , n236 , n237 , n238 , n239 , n240 , n241 , n242 ;
output n243 , n244 , n245 , n246 , n247 , n248 , n249 , n250 , n251 , n252 , n253 , n254 , n255 , n256 , n257 ;

wire n516 , n517 , n518 , n519 , n520 , n521 , n522 , n523 , n524 ,
     n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 , n533 , n534 ,
     n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 , n543 , n544 ,
     n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 , n553 , n554 ,
     n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 , n563 , n564 ,
     n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 , n573 , n574 ,
     n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 , n583 , n584 ,
     n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 , n593 , n594 ,
     n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 , n603 , n604 ,
     n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 , n613 , n614 ,
     n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 , n623 , n624 ,
     n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 , n633 , n634 ,
     n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 , n643 , n644 ,
     n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 , n653 , n654 ,
     n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 , n663 , n664 ,
     n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 , n673 , n674 ,
     n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 , n683 , n684 ,
     n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 , n693 , n694 ,
     n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 , n703 , n704 ,
     n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 , n713 , n714 ,
     n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 , n723 , n724 ,
     n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 , n733 , n734 ,
     n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 , n743 , n744 ,
     n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 , n753 , n754 ,
     n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 , n763 , n764 ,
     n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 , n773 , n774 ,
     n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 , n783 , n784 ,
     n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 , n793 , n794 ,
     n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 , n803 , n804 ,
     n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 , n813 , n814 ,
     n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 , n823 , n824 ,
     n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 , n833 , n834 ,
     n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 , n843 , n844 ,
     n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 , n853 , n854 ,
     n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 , n863 , n864 ,
     n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 , n873 , n874 ,
     n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 , n883 , n884 ,
     n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 , n893 , n894 ,
     n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 , n903 , n904 ,
     n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 , n913 , n914 ,
     n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 , n923 , n924 ,
     n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 , n933 , n934 ,
     n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 , n943 , n944 ,
     n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 , n953 , n954 ,
     n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 , n963 , n964 ,
     n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 , n973 , n974 ,
     n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 , n983 , n984 ,
     n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 , n993 , n994 ,
     n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 , n1003 , n1004 ,
     n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 , n1013 , n1014 ,
     n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 , n1023 , n1024 ,
     n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 , n1033 , n1034 ,
     n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 , n1043 , n1044 ,
     n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 , n1053 , n1054 ,
     n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 , n1063 , n1064 ,
     n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 , n1073 , n1074 ,
     n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 , n1083 , n1084 ,
     n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 , n1093 , n1094 ,
     n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 , n1103 , n1104 ,
     n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 , n1113 , n1114 ,
     n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 , n1123 , n1124 ,
     n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 , n1133 , n1134 ,
     n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 , n1143 , n1144 ,
     n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 , n1153 , n1154 ,
     n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 , n1163 , n1164 ,
     n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 , n1173 , n1174 ,
     n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 , n1183 , n1184 ,
     n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 , n1193 , n1194 ,
     n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 , n1203 , n1204 ,
     n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 , n1213 , n1214 ,
     n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 , n1223 , n1224 ,
     n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 , n1233 , n1234 ,
     n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 , n1243 , n1244 ,
     n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 , n1253 , n1254 ,
     n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 , n1263 , n1264 ,
     n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 , n1273 , n1274 ,
     n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 , n1283 , n1284 ,
     n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 , n1293 , n1294 ,
     n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 , n1303 , n1304 ,
     n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 , n1313 , n1314 ,
     n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 , n1323 , n1324 ,
     n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 , n1333 , n1334 ,
     n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 , n1343 , n1344 ,
     n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 , n1353 , n1354 ,
     n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 , n1363 , n1364 ,
     n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 , n1373 , n1374 ,
     n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 , n1383 , n1384 ,
     n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 , n1393 , n1394 ,
     n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 , n1403 , n1404 ,
     n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 , n1413 , n1414 ,
     n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 , n1423 , n1424 ,
     n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 , n1433 , n1434 ,
     n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 , n1443 , n1444 ,
     n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 , n1453 , n1454 ,
     n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 , n1463 , n1464 ,
     n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 , n1473 , n1474 ,
     n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 , n1483 , n1484 ,
     n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 , n1493 , n1494 ,
     n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 , n1503 , n1504 ,
     n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 , n1513 , n1514 ,
     n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 , n1523 , n1524 ,
     n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 , n1533 , n1534 ,
     n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 , n1543 , n1544 ,
     n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 , n1553 , n1554 ,
     n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 , n1563 , n1564 ,
     n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 , n1573 , n1574 ,
     n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 , n1583 , n1584 ,
     n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 , n1593 , n1594 ,
     n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 , n1603 , n1604 ,
     n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 , n1613 , n1614 ,
     n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 , n1623 , n1624 ,
     n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 , n1633 , n1634 ,
     n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 , n1643 , n1644 ,
     n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 , n1653 , n1654 ,
     n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 , n1663 , n1664 ,
     n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 , n1673 , n1674 ,
     n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 , n1683 , n1684 ,
     n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 , n1693 , n1694 ,
     n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 , n1703 , n1704 ,
     n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 , n1713 , n1714 ,
     n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 , n1723 , n1724 ,
     n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 , n1733 , n1734 ,
     n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 , n1743 , n1744 ,
     n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 , n1753 , n1754 ,
     n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 , n1763 , n1764 ,
     n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 , n1773 , n1774 ,
     n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 , n1783 , n1784 ,
     n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 , n1793 , n1794 ,
     n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 , n1803 , n1804 ,
     n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 , n1813 , n1814 ,
     n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 , n1823 , n1824 ,
     n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 , n1833 , n1834 ,
     n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 , n1843 , n1844 ,
     n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 , n1853 , n1854 ,
     n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 , n1863 , n1864 ,
     n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 , n1873 , n1874 ,
     n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 , n1883 , n1884 ,
     n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 , n1893 , n1894 ,
     n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 , n1903 , n1904 ,
     n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 , n1913 , n1914 ,
     n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 , n1923 , n1924 ,
     n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 , n1933 , n1934 ,
     n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 , n1943 , n1944 ,
     n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 , n1953 , n1954 ,
     n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 , n1963 , n1964 ,
     n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 , n1973 , n1974 ,
     n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 , n1983 , n1984 ,
     n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 , n1993 , n1994 ,
     n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 , n2003 , n2004 ,
     n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 , n2013 , n2014 ,
     n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 , n2023 , n2024 ,
     n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 , n2033 , n2034 ,
     n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 , n2043 , n2044 ,
     n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 , n2053 , n2054 ,
     n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 , n2063 , n2064 ,
     n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 , n2073 , n2074 ,
     n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 , n2083 , n2084 ,
     n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 , n2093 , n2094 ,
     n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 , n2103 , n2104 ,
     n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 , n2113 , n2114 ,
     n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 , n2123 , n2124 ,
     n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 , n2133 , n2134 ,
     n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 , n2143 , n2144 ,
     n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 , n2153 , n2154 ,
     n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 , n2163 , n2164 ,
     n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 , n2173 , n2174 ,
     n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 , n2183 , n2184 ,
     n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 , n2193 , n2194 ,
     n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 , n2203 , n2204 ,
     n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 , n2213 , n2214 ,
     n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 , n2223 , n2224 ,
     n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 , n2233 , n2234 ,
     n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 , n2243 , n2244 ,
     n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 , n2253 , n2254 ,
     n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 , n2263 , n2264 ,
     n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 , n2273 , n2274 ,
     n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 , n2283 , n2284 ,
     n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 , n2293 , n2294 ,
     n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 , n2303 , n2304 ,
     n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 , n2313 , n2314 ,
     n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 , n2323 , n2324 ,
     n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 , n2333 , n2334 ,
     n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 , n2343 , n2344 ,
     n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 , n2353 , n2354 ,
     n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 , n2363 , n2364 ,
     n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 , n2373 , n2374 ,
     n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 , n2383 , n2384 ,
     n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 , n2393 , n2394 ,
     n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 , n2403 , n2404 ,
     n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 , n2413 , n2414 ,
     n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 , n2423 , n2424 ,
     n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 , n2433 , n2434 ,
     n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 , n2443 , n2444 ,
     n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 , n2453 , n2454 ,
     n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 , n2463 , n2464 ,
     n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 , n2473 , n2474 ,
     n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 , n2483 , n2484 ,
     n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 , n2493 , n2494 ,
     n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 , n2503 , n2504 ,
     n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 , n2513 , n2514 ,
     n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 , n2523 , n2524 ,
     n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 , n2533 , n2534 ,
     n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 , n2543 , n2544 ,
     n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 , n2553 , n2554 ,
     n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 , n2563 , n2564 ,
     n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 , n2573 , n2574 ,
     n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 , n2583 , n2584 ,
     n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 , n2593 , n2594 ,
     n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 , n2603 , n2604 ,
     n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 , n2613 , n2614 ,
     n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 , n2623 , n2624 ,
     n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 , n2633 , n2634 ,
     n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 , n2643 , n2644 ,
     n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 , n2653 , n2654 ,
     n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 , n2663 , n2664 ,
     n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 , n2673 , n2674 ,
     n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 , n2683 , n2684 ,
     n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 , n2693 , n2694 ,
     n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 , n2703 , n2704 ,
     n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 , n2713 , n2714 ,
     n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 , n2723 , n2724 ,
     n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 , n2733 , n2734 ,
     n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 , n2743 , n2744 ,
     n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 , n2753 , n2754 ,
     n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 , n2763 , n2764 ,
     n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 , n2773 , n2774 ,
     n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 , n2783 , n2784 ,
     n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 , n2793 , n2794 ,
     n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 , n2803 , n2804 ,
     n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 , n2813 , n2814 ,
     n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 , n2823 , n2824 ,
     n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 , n2833 , n2834 ,
     n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 , n2843 , n2844 ,
     n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 , n2853 , n2854 ,
     n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 , n2863 , n2864 ,
     n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 , n2873 , n2874 ,
     n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 , n2883 , n2884 ,
     n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 , n2893 , n2894 ,
     n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 , n2903 , n2904 ,
     n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 , n2913 , n2914 ,
     n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 , n2923 , n2924 ,
     n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 , n2933 , n2934 ,
     n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 , n2943 , n2944 ,
     n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 , n2953 , n2954 ,
     n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 , n2963 , n2964 ,
     n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 , n2973 , n2974 ,
     n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 , n2983 , n2984 ,
     n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 , n2993 , n2994 ,
     n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 , n3003 , n3004 ,
     n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 , n3013 , n3014 ,
     n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 , n3023 , n3024 ,
     n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 , n3033 , n3034 ,
     n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 , n3043 , n3044 ,
     n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 , n3053 , n3054 ,
     n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 , n3063 , n3064 ,
     n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 , n3073 , n3074 ,
     n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 , n3083 , n3084 ,
     n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 , n3093 , n3094 ,
     n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 , n3103 , n3104 ,
     n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 , n3113 , n3114 ,
     n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 , n3123 , n3124 ,
     n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 , n3133 , n3134 ,
     n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 , n3143 , n3144 ,
     n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 , n3153 , n3154 ,
     n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 , n3163 , n3164 ,
     n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 , n3173 , n3174 ,
     n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 , n3183 , n3184 ,
     n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 , n3193 , n3194 ,
     n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 , n3203 , n3204 ,
     n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 , n3213 , n3214 ,
     n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 , n3223 , n3224 ,
     n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 , n3233 , n3234 ,
     n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 , n3243 , n3244 ,
     n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 , n3253 , n3254 ,
     n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 , n3263 , n3264 ,
     n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 , n3273 , n3274 ,
     n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 , n3283 , n3284 ,
     n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 , n3293 , n3294 ,
     n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 , n3303 , n3304 ,
     n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 , n3313 , n3314 ,
     n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 , n3323 , n3324 ,
     n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 , n3333 , n3334 ,
     n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 , n3343 , n3344 ,
     n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 , n3353 , n3354 ,
     n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 , n3363 , n3364 ,
     n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 , n3373 , n3374 ,
     n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 , n3383 , n3384 ,
     n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 , n3393 , n3394 ,
     n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 , n3403 , n3404 ,
     n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 , n3413 , n3414 ,
     n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 , n3423 , n3424 ,
     n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 , n3433 , n3434 ,
     n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 , n3443 , n3444 ,
     n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 , n3453 , n3454 ,
     n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 , n3463 , n3464 ,
     n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 , n3473 , n3474 ,
     n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 , n3483 , n3484 ,
     n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 , n3493 , n3494 ,
     n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 , n3503 , n3504 ,
     n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 , n3513 , n3514 ,
     n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 , n3523 , n3524 ,
     n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 , n3533 , n3534 ,
     n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 , n3543 , n3544 ,
     n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 , n3553 , n3554 ,
     n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 , n3563 , n3564 ,
     n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 , n3573 , n3574 ,
     n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 , n3583 , n3584 ,
     n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 , n3593 , n3594 ,
     n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 , n3603 , n3604 ,
     n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 , n3613 , n3614 ,
     n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 , n3623 , n3624 ,
     n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 , n3633 , n3634 ,
     n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 , n3643 , n3644 ,
     n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 , n3653 , n3654 ,
     n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 , n3663 , n3664 ,
     n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 , n3673 , n3674 ,
     n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 , n3683 , n3684 ,
     n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 , n3693 , n3694 ,
     n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 , n3703 , n3704 ,
     n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 , n3713 , n3714 ,
     n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 , n3723 , n3724 ,
     n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 , n3733 , n3734 ,
     n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 , n3743 , n3744 ,
     n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 , n3753 , n3754 ,
     n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 , n3763 , n3764 ,
     n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 , n3773 , n3774 ,
     n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 , n3783 , n3784 ,
     n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 , n3793 , n3794 ,
     n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 , n3803 , n3804 ,
     n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 , n3813 , n3814 ,
     n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 , n3823 , n3824 ,
     n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 , n3833 , n3834 ,
     n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 , n3843 , n3844 ,
     n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 , n3853 , n3854 ,
     n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 , n3863 , n3864 ,
     n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 , n3873 , n3874 ,
     n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 , n3883 , n3884 ,
     n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 , n3893 , n3894 ,
     n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 , n3903 , n3904 ,
     n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 , n3913 , n3914 ,
     n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 , n3923 , n3924 ,
     n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 , n3933 , n3934 ,
     n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 , n3943 , n3944 ,
     n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 , n3953 , n3954 ,
     n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 , n3963 , n3964 ,
     n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 , n3973 , n3974 ,
     n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 , n3983 , n3984 ,
     n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 , n3993 , n3994 ,
     n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 , n4003 , n4004 ,
     n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 , n4013 , n4014 ,
     n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 , n4023 , n4024 ,
     n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 , n4033 , n4034 ,
     n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 , n4043 , n4044 ,
     n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 , n4053 , n4054 ,
     n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 , n4063 , n4064 ,
     n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 , n4073 , n4074 ,
     n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 , n4083 , n4084 ,
     n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 , n4093 , n4094 ,
     n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 , n4103 , n4104 ,
     n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 , n4113 , n4114 ,
     n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 , n4123 , n4124 ,
     n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 , n4133 , n4134 ,
     n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 , n4143 , n4144 ,
     n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 , n4153 , n4154 ,
     n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 , n4163 , n4164 ,
     n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 , n4173 , n4174 ,
     n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 , n4183 , n4184 ,
     n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 , n4193 , n4194 ,
     n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 , n4203 , n4204 ,
     n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 , n4213 , n4214 ,
     n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 , n4223 , n4224 ,
     n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 , n4233 , n4234 ,
     n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 , n4243 , n4244 ,
     n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 , n4253 , n4254 ,
     n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 , n4263 , n4264 ,
     n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 , n4273 , n4274 ,
     n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 , n4283 , n4284 ,
     n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 , n4293 , n4294 ,
     n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 , n4303 , n4304 ,
     n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 , n4313 , n4314 ,
     n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 , n4323 , n4324 ,
     n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 , n4333 , n4334 ,
     n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 , n4343 , n4344 ,
     n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 , n4353 , n4354 ,
     n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 , n4363 , n4364 ,
     n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 , n4373 , n4374 ,
     n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 , n4383 , n4384 ,
     n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 , n4393 , n4394 ,
     n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 , n4403 , n4404 ,
     n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 , n4413 , n4414 ,
     n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 , n4423 , n4424 ,
     n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 , n4433 , n4434 ,
     n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 , n4443 , n4444 ,
     n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 , n4453 , n4454 ,
     n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 , n4463 , n4464 ,
     n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 , n4473 , n4474 ,
     n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 , n4483 , n4484 ,
     n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 , n4493 , n4494 ,
     n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 , n4503 , n4504 ,
     n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 , n4513 , n4514 ,
     n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 , n4523 , n4524 ,
     n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 , n4533 , n4534 ,
     n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 , n4543 , n4544 ,
     n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 , n4553 , n4554 ,
     n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 , n4563 , n4564 ,
     n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 , n4573 , n4574 ,
     n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 , n4583 , n4584 ,
     n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 , n4593 , n4594 ,
     n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 , n4603 , n4604 ,
     n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 , n4613 , n4614 ,
     n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 , n4623 , n4624 ,
     n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 , n4633 , n4634 ,
     n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 , n4643 , n4644 ,
     n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 , n4653 , n4654 ,
     n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 , n4663 , n4664 ,
     n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 , n4673 , n4674 ,
     n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 , n4683 , n4684 ,
     n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 , n4693 , n4694 ,
     n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 , n4703 , n4704 ,
     n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 , n4713 , n4714 ,
     n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 , n4723 , n4724 ,
     n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 , n4733 , n4734 ,
     n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 , n4743 , n4744 ,
     n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 , n4753 , n4754 ,
     n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 , n4763 , n4764 ,
     n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 , n4773 , n4774 ,
     n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 , n4783 , n4784 ,
     n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 , n4793 , n4794 ,
     n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 , n4803 , n4804 ,
     n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 , n4813 , n4814 ,
     n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 , n4823 , n4824 ,
     n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 , n4833 , n4834 ,
     n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 , n4843 , n4844 ,
     n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 , n4853 , n4854 ,
     n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 , n4863 , n4864 ,
     n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 , n4873 , n4874 ,
     n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 , n4883 , n4884 ,
     n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 , n4893 , n4894 ,
     n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 , n4903 , n4904 ,
     n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 , n4913 , n4914 ,
     n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 , n4923 , n4924 ,
     n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 , n4933 , n4934 ,
     n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 , n4943 , n4944 ,
     n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 , n4953 , n4954 ,
     n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 , n4963 , n4964 ,
     n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 , n4973 , n4974 ,
     n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 , n4983 , n4984 ,
     n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 , n4993 , n4994 ,
     n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 , n5003 , n5004 ,
     n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 , n5013 , n5014 ,
     n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 , n5023 , n5024 ,
     n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 , n5033 , n5034 ,
     n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 , n5043 , n5044 ,
     n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 , n5053 , n5054 ,
     n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 , n5063 , n5064 ,
     n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 , n5073 , n5074 ,
     n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 , n5083 , n5084 ,
     n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 , n5093 , n5094 ,
     n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 , n5103 , n5104 ,
     n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 , n5113 , n5114 ,
     n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 , n5123 , n5124 ,
     n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 , n5133 , n5134 ,
     n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 , n5143 , n5144 ,
     n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 , n5153 , n5154 ,
     n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 , n5163 , n5164 ,
     n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 , n5173 , n5174 ,
     n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 , n5183 , n5184 ,
     n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 , n5193 , n5194 ,
     n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 , n5203 , n5204 ,
     n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 , n5213 , n5214 ,
     n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 , n5223 , n5224 ,
     n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 , n5233 , n5234 ,
     n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 , n5243 , n5244 ,
     n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 , n5253 , n5254 ,
     n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 , n5263 , n5264 ,
     n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 , n5273 , n5274 ,
     n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 , n5283 , n5284 ,
     n5285 , n5286 , n5287 , n5288 , n5289 , n5290 ;
buf ( n256 , n848 );
buf ( n255 , n5067 );
buf ( n257 , 1'b0 );
buf ( n254 , n5069 );
buf ( n252 , n5070 );
buf ( n244 , n5142 );
buf ( n251 , 1'b0 );
buf ( n243 , n5143 );
buf ( n246 , n5144 );
buf ( n248 , n5216 );
buf ( n247 , 1'b0 );
buf ( n249 , n5217 );
buf ( n250 , n5218 );
buf ( n253 , n5290 );
buf ( n245 , 1'b0 );
buf ( n652 , PI_PI_clock);
buf ( n653 , PI_PI_reset);
buf ( n654 , n6 );
buf ( n655 , n50 );
buf ( n656 , n58 );
buf ( n657 , n76 );
buf ( n658 , n71 );
buf ( n659 , n163 );
buf ( n660 , n234 );
buf ( n661 , n39 );
buf ( n662 , n225 );
buf ( n663 , n144 );
buf ( n664 , n156 );
buf ( n665 , n217 );
buf ( n666 , n194 );
buf ( n667 , n114 );
buf ( n668 , n17 );
buf ( n669 , n160 );
buf ( n670 , n209 );
buf ( n671 , n137 );
buf ( n672 , n167 );
buf ( n673 , n140 );
buf ( n674 , n147 );
buf ( n675 , n195 );
buf ( n676 , n60 );
buf ( n677 , n73 );
buf ( n678 , n242 );
buf ( n679 , n25 );
buf ( n680 , n223 );
buf ( n681 , n150 );
buf ( n682 , n227 );
buf ( n683 , n92 );
buf ( n684 , n54 );
buf ( n685 , n123 );
buf ( n686 , PI_DFF_state_reg_Q);
buf ( n687 , n190 );
buf ( n688 , n237 );
buf ( n689 , n183 );
buf ( n690 , n161 );
buf ( n691 , n86 );
buf ( n692 , n91 );
buf ( n693 , n178 );
buf ( n694 , n119 );
buf ( n695 , n11 );
buf ( n696 , n218 );
buf ( n697 , n192 );
buf ( n698 , n166 );
buf ( n699 , n63 );
buf ( n700 , n145 );
buf ( n701 , n38 );
buf ( n702 , n1 );
buf ( n703 , n3 );
buf ( n704 , n122 );
buf ( n705 , n40 );
buf ( n706 , n230 );
buf ( n707 , n228 );
buf ( n708 , n138 );
buf ( n709 , n32 );
buf ( n710 , n168 );
buf ( n711 , n0 );
buf ( n712 , n61 );
buf ( n713 , n26 );
buf ( n714 , n191 );
buf ( n715 , n68 );
buf ( n716 , n204 );
buf ( n717 , n197 );
buf ( n718 , n128 );
buf ( n719 , n34 );
buf ( n720 , n141 );
buf ( n721 , n108 );
buf ( n722 , n42 );
buf ( n723 , n117 );
buf ( n724 , n151 );
buf ( n725 , n198 );
buf ( n726 , n74 );
buf ( n727 , n111 );
buf ( n728 , n16 );
buf ( n729 , n79 );
buf ( n730 , n15 );
buf ( n731 , n52 );
buf ( n732 , n72 );
buf ( n733 , n124 );
buf ( n734 , n19 );
buf ( n735 , n98 );
buf ( n736 , n31 );
buf ( n737 , n81 );
buf ( n738 , n14 );
buf ( n739 , n200 );
buf ( n740 , n220 );
buf ( n741 , n43 );
buf ( n742 , n224 );
buf ( n743 , n233 );
buf ( n744 , n196 );
buf ( n745 , n132 );
buf ( n746 , n184 );
buf ( n747 , n94 );
buf ( n748 , n109 );
buf ( n749 , n21 );
buf ( n750 , n10 );
buf ( n751 , n95 );
buf ( n752 , n110 );
buf ( n753 , n78 );
buf ( n754 , n29 );
buf ( n755 , n189 );
buf ( n756 , n212 );
buf ( n757 , n51 );
buf ( n758 , n49 );
buf ( n759 , n77 );
buf ( n760 , n90 );
buf ( n761 , n4 );
buf ( n762 , n148 );
buf ( n763 , n7 );
buf ( n764 , n181 );
buf ( n765 , n9 );
buf ( n766 , n87 );
buf ( n767 , n232 );
buf ( n768 , n177 );
buf ( n769 , n240 );
buf ( n770 , n105 );
buf ( n771 , n236 );
buf ( n772 , n45 );
buf ( n773 , n30 );
buf ( n774 , n57 );
buf ( n775 , n65 );
buf ( n776 , n241 );
buf ( n777 , n202 );
buf ( n778 , n18 );
buf ( n779 , n106 );
buf ( n780 , n149 );
buf ( n781 , n113 );
buf ( n782 , n23 );
buf ( n783 , n101 );
buf ( n784 , n206 );
buf ( n785 , n2 );
buf ( n786 , n231 );
buf ( n787 , n70 );
buf ( n788 , n59 );
buf ( n789 , n180 );
buf ( n790 , n12 );
buf ( n791 , n172 );
buf ( n792 , n219 );
buf ( n793 , n80 );
buf ( n794 , n121 );
buf ( n795 , n8 );
buf ( n796 , n36 );
buf ( n797 , n207 );
buf ( n798 , n53 );
buf ( n799 , n69 );
buf ( n800 , n107 );
buf ( n801 , n176 );
buf ( n802 , n64 );
buf ( n803 , n136 );
buf ( n804 , n55 );
buf ( n805 , n130 );
buf ( n806 , n125 );
buf ( n807 , n157 );
buf ( n808 , n100 );
buf ( n809 , n99 );
buf ( n810 , n187 );
buf ( n811 , n96 );
buf ( n812 , n154 );
buf ( n813 , n164 );
buf ( n814 , PI_DFF_B_reg_Q);
buf ( n815 , n214 );
buf ( n816 , n135 );
buf ( n817 , n46 );
buf ( n818 , n5 );
buf ( n819 , n24 );
buf ( n820 , n13 );
buf ( n821 , n222 );
buf ( n822 , n118 );
buf ( n823 , n97 );
buf ( n824 , n238 );
buf ( n825 , n169 );
buf ( n826 , n133 );
buf ( n827 , n89 );
buf ( n828 , n142 );
buf ( n829 , n146 );
buf ( n830 , n213 );
buf ( n831 , n188 );
buf ( n832 , n44 );
buf ( n833 , n28 );
buf ( n834 , n112 );
buf ( n835 , n22 );
buf ( n836 , n171 );
buf ( n837 , n179 );
buf ( n838 , n162 );
buf ( n839 , n102 );
buf ( n840 , n186 );
buf ( n841 , n175 );
buf ( n842 , n203 );
buf ( n843 , n83 );
buf ( n844 , n153 );
buf ( n845 , n67 );
buf ( n846 , n210 );
buf ( n847 , n652 );
buf ( n848 , n847 );
buf ( n849 , n718 );
not ( n850 , n849 );
buf ( n851 , n717 );
not ( n852 , n851 );
buf ( n853 , n716 );
not ( n854 , n853 );
buf ( n855 , n715 );
not ( n856 , n855 );
buf ( n857 , n714 );
not ( n858 , n857 );
buf ( n859 , n713 );
not ( n860 , n859 );
buf ( n861 , n712 );
not ( n862 , n861 );
buf ( n863 , n711 );
not ( n864 , n863 );
buf ( n865 , n710 );
not ( n866 , n865 );
buf ( n867 , n709 );
not ( n868 , n867 );
buf ( n869 , n708 );
not ( n870 , n869 );
buf ( n871 , n707 );
not ( n872 , n871 );
buf ( n873 , n706 );
not ( n874 , n873 );
buf ( n875 , n705 );
not ( n876 , n875 );
buf ( n877 , n704 );
not ( n878 , n877 );
buf ( n879 , n703 );
not ( n880 , n879 );
buf ( n881 , n702 );
not ( n882 , n881 );
buf ( n883 , n701 );
not ( n884 , n883 );
buf ( n885 , n700 );
not ( n886 , n885 );
buf ( n887 , n699 );
not ( n888 , n887 );
buf ( n889 , n698 );
not ( n890 , n889 );
buf ( n891 , n697 );
not ( n892 , n891 );
buf ( n893 , n696 );
not ( n894 , n893 );
buf ( n895 , n695 );
not ( n896 , n895 );
buf ( n897 , n694 );
not ( n898 , n897 );
buf ( n899 , n693 );
not ( n900 , n899 );
buf ( n901 , n692 );
not ( n902 , n901 );
buf ( n903 , n691 );
not ( n904 , n903 );
buf ( n905 , n690 );
not ( n906 , n905 );
buf ( n907 , n689 );
not ( n908 , n907 );
buf ( n909 , n688 );
not ( n910 , n909 );
buf ( n911 , n687 );
not ( n912 , n911 );
and ( n913 , n910 , n912 );
and ( n914 , n908 , n913 );
and ( n915 , n906 , n914 );
and ( n916 , n904 , n915 );
and ( n917 , n902 , n916 );
and ( n918 , n900 , n917 );
and ( n919 , n898 , n918 );
and ( n920 , n896 , n919 );
and ( n921 , n894 , n920 );
and ( n922 , n892 , n921 );
and ( n923 , n890 , n922 );
and ( n924 , n888 , n923 );
and ( n925 , n886 , n924 );
and ( n926 , n884 , n925 );
and ( n927 , n882 , n926 );
and ( n928 , n880 , n927 );
and ( n929 , n878 , n928 );
and ( n930 , n876 , n929 );
and ( n931 , n874 , n930 );
and ( n932 , n872 , n931 );
and ( n933 , n870 , n932 );
and ( n934 , n868 , n933 );
and ( n935 , n866 , n934 );
and ( n936 , n864 , n935 );
and ( n937 , n862 , n936 );
and ( n938 , n860 , n937 );
and ( n939 , n858 , n938 );
and ( n940 , n856 , n939 );
and ( n941 , n854 , n940 );
and ( n942 , n852 , n941 );
xor ( n943 , n850 , n942 );
buf ( n944 , n849 );
and ( n945 , n943 , n944 );
buf ( n946 , n945 );
not ( n947 , n946 );
not ( n948 , n849 );
and ( n949 , n948 , n865 );
xor ( n950 , n866 , n934 );
and ( n951 , n950 , n849 );
or ( n952 , n949 , n951 );
and ( n953 , n947 , n952 );
not ( n954 , n952 );
not ( n955 , n849 );
and ( n956 , n955 , n867 );
xor ( n957 , n868 , n933 );
and ( n958 , n957 , n849 );
or ( n959 , n956 , n958 );
not ( n960 , n959 );
not ( n961 , n849 );
and ( n962 , n961 , n869 );
xor ( n963 , n870 , n932 );
and ( n964 , n963 , n849 );
or ( n965 , n962 , n964 );
not ( n966 , n965 );
not ( n967 , n849 );
and ( n968 , n967 , n871 );
xor ( n969 , n872 , n931 );
and ( n970 , n969 , n849 );
or ( n971 , n968 , n970 );
not ( n972 , n971 );
not ( n973 , n849 );
and ( n974 , n973 , n873 );
xor ( n975 , n874 , n930 );
and ( n976 , n975 , n849 );
or ( n977 , n974 , n976 );
not ( n978 , n977 );
not ( n979 , n849 );
and ( n980 , n979 , n875 );
xor ( n981 , n876 , n929 );
and ( n982 , n981 , n849 );
or ( n983 , n980 , n982 );
not ( n984 , n983 );
not ( n985 , n849 );
and ( n986 , n985 , n877 );
xor ( n987 , n878 , n928 );
and ( n988 , n987 , n849 );
or ( n989 , n986 , n988 );
not ( n990 , n989 );
not ( n991 , n849 );
and ( n992 , n991 , n879 );
xor ( n993 , n880 , n927 );
and ( n994 , n993 , n849 );
or ( n995 , n992 , n994 );
not ( n996 , n995 );
not ( n997 , n849 );
and ( n998 , n997 , n881 );
xor ( n999 , n882 , n926 );
and ( n1000 , n999 , n849 );
or ( n1001 , n998 , n1000 );
not ( n1002 , n1001 );
not ( n1003 , n849 );
and ( n1004 , n1003 , n883 );
xor ( n1005 , n884 , n925 );
and ( n1006 , n1005 , n849 );
or ( n1007 , n1004 , n1006 );
not ( n1008 , n1007 );
not ( n1009 , n849 );
and ( n1010 , n1009 , n885 );
xor ( n1011 , n886 , n924 );
and ( n1012 , n1011 , n849 );
or ( n1013 , n1010 , n1012 );
not ( n1014 , n1013 );
not ( n1015 , n849 );
and ( n1016 , n1015 , n887 );
xor ( n1017 , n888 , n923 );
and ( n1018 , n1017 , n849 );
or ( n1019 , n1016 , n1018 );
not ( n1020 , n1019 );
not ( n1021 , n849 );
and ( n1022 , n1021 , n889 );
xor ( n1023 , n890 , n922 );
and ( n1024 , n1023 , n849 );
or ( n1025 , n1022 , n1024 );
not ( n1026 , n1025 );
not ( n1027 , n849 );
and ( n1028 , n1027 , n891 );
xor ( n1029 , n892 , n921 );
and ( n1030 , n1029 , n849 );
or ( n1031 , n1028 , n1030 );
not ( n1032 , n1031 );
not ( n1033 , n849 );
and ( n1034 , n1033 , n893 );
xor ( n1035 , n894 , n920 );
and ( n1036 , n1035 , n849 );
or ( n1037 , n1034 , n1036 );
not ( n1038 , n1037 );
not ( n1039 , n849 );
and ( n1040 , n1039 , n895 );
xor ( n1041 , n896 , n919 );
and ( n1042 , n1041 , n849 );
or ( n1043 , n1040 , n1042 );
not ( n1044 , n1043 );
not ( n1045 , n849 );
and ( n1046 , n1045 , n897 );
xor ( n1047 , n898 , n918 );
and ( n1048 , n1047 , n849 );
or ( n1049 , n1046 , n1048 );
not ( n1050 , n1049 );
not ( n1051 , n849 );
and ( n1052 , n1051 , n899 );
xor ( n1053 , n900 , n917 );
and ( n1054 , n1053 , n849 );
or ( n1055 , n1052 , n1054 );
not ( n1056 , n1055 );
not ( n1057 , n849 );
and ( n1058 , n1057 , n901 );
xor ( n1059 , n902 , n916 );
and ( n1060 , n1059 , n849 );
or ( n1061 , n1058 , n1060 );
not ( n1062 , n1061 );
not ( n1063 , n849 );
and ( n1064 , n1063 , n903 );
xor ( n1065 , n904 , n915 );
and ( n1066 , n1065 , n849 );
or ( n1067 , n1064 , n1066 );
not ( n1068 , n1067 );
not ( n1069 , n849 );
and ( n1070 , n1069 , n905 );
xor ( n1071 , n906 , n914 );
and ( n1072 , n1071 , n849 );
or ( n1073 , n1070 , n1072 );
not ( n1074 , n1073 );
not ( n1075 , n849 );
and ( n1076 , n1075 , n907 );
xor ( n1077 , n908 , n913 );
and ( n1078 , n1077 , n849 );
or ( n1079 , n1076 , n1078 );
not ( n1080 , n1079 );
not ( n1081 , n849 );
and ( n1082 , n1081 , n909 );
xor ( n1083 , n910 , n912 );
and ( n1084 , n1083 , n849 );
or ( n1085 , n1082 , n1084 );
not ( n1086 , n1085 );
not ( n1087 , n911 );
and ( n1088 , n1086 , n1087 );
and ( n1089 , n1080 , n1088 );
and ( n1090 , n1074 , n1089 );
and ( n1091 , n1068 , n1090 );
and ( n1092 , n1062 , n1091 );
and ( n1093 , n1056 , n1092 );
and ( n1094 , n1050 , n1093 );
and ( n1095 , n1044 , n1094 );
and ( n1096 , n1038 , n1095 );
and ( n1097 , n1032 , n1096 );
and ( n1098 , n1026 , n1097 );
and ( n1099 , n1020 , n1098 );
and ( n1100 , n1014 , n1099 );
and ( n1101 , n1008 , n1100 );
and ( n1102 , n1002 , n1101 );
and ( n1103 , n996 , n1102 );
and ( n1104 , n990 , n1103 );
and ( n1105 , n984 , n1104 );
and ( n1106 , n978 , n1105 );
and ( n1107 , n972 , n1106 );
and ( n1108 , n966 , n1107 );
and ( n1109 , n960 , n1108 );
xor ( n1110 , n954 , n1109 );
and ( n1111 , n1110 , n946 );
or ( n1112 , n953 , n1111 );
not ( n1113 , n1112 );
not ( n1114 , n1113 );
not ( n1115 , n1114 );
not ( n1116 , n1115 );
buf ( n1117 , n1116 );
buf ( n1118 , n1117 );
not ( n1119 , n946 );
not ( n1120 , n849 );
and ( n1121 , n1120 , n851 );
xor ( n1122 , n852 , n941 );
and ( n1123 , n1122 , n849 );
or ( n1124 , n1121 , n1123 );
not ( n1125 , n1124 );
not ( n1126 , n849 );
and ( n1127 , n1126 , n853 );
xor ( n1128 , n854 , n940 );
and ( n1129 , n1128 , n849 );
or ( n1130 , n1127 , n1129 );
not ( n1131 , n1130 );
not ( n1132 , n849 );
and ( n1133 , n1132 , n855 );
xor ( n1134 , n856 , n939 );
and ( n1135 , n1134 , n849 );
or ( n1136 , n1133 , n1135 );
not ( n1137 , n1136 );
not ( n1138 , n849 );
and ( n1139 , n1138 , n857 );
xor ( n1140 , n858 , n938 );
and ( n1141 , n1140 , n849 );
or ( n1142 , n1139 , n1141 );
not ( n1143 , n1142 );
not ( n1144 , n849 );
and ( n1145 , n1144 , n859 );
xor ( n1146 , n860 , n937 );
and ( n1147 , n1146 , n849 );
or ( n1148 , n1145 , n1147 );
not ( n1149 , n1148 );
not ( n1150 , n849 );
and ( n1151 , n1150 , n861 );
xor ( n1152 , n862 , n936 );
and ( n1153 , n1152 , n849 );
or ( n1154 , n1151 , n1153 );
not ( n1155 , n1154 );
not ( n1156 , n849 );
and ( n1157 , n1156 , n863 );
xor ( n1158 , n864 , n935 );
and ( n1159 , n1158 , n849 );
or ( n1160 , n1157 , n1159 );
not ( n1161 , n1160 );
and ( n1162 , n954 , n1109 );
and ( n1163 , n1161 , n1162 );
and ( n1164 , n1155 , n1163 );
and ( n1165 , n1149 , n1164 );
and ( n1166 , n1143 , n1165 );
and ( n1167 , n1137 , n1166 );
and ( n1168 , n1131 , n1167 );
and ( n1169 , n1125 , n1168 );
xor ( n1170 , n1119 , n1169 );
buf ( n1171 , n946 );
and ( n1172 , n1170 , n1171 );
buf ( n1173 , n1172 );
not ( n1174 , n1173 );
not ( n1175 , n1174 );
not ( n1176 , n1175 );
not ( n1177 , n946 );
and ( n1178 , n1177 , n1124 );
xor ( n1179 , n1125 , n1168 );
and ( n1180 , n1179 , n946 );
or ( n1181 , n1178 , n1180 );
not ( n1182 , n1181 );
not ( n1183 , n1182 );
not ( n1184 , n1183 );
not ( n1185 , n946 );
and ( n1186 , n1185 , n1130 );
xor ( n1187 , n1131 , n1167 );
and ( n1188 , n1187 , n946 );
or ( n1189 , n1186 , n1188 );
not ( n1190 , n1189 );
not ( n1191 , n1190 );
not ( n1192 , n1191 );
not ( n1193 , n946 );
and ( n1194 , n1193 , n1136 );
xor ( n1195 , n1137 , n1166 );
and ( n1196 , n1195 , n946 );
or ( n1197 , n1194 , n1196 );
not ( n1198 , n1197 );
not ( n1199 , n1198 );
not ( n1200 , n1199 );
not ( n1201 , n946 );
and ( n1202 , n1201 , n1142 );
xor ( n1203 , n1143 , n1165 );
and ( n1204 , n1203 , n946 );
or ( n1205 , n1202 , n1204 );
not ( n1206 , n1205 );
not ( n1207 , n1206 );
not ( n1208 , n1207 );
not ( n1209 , n946 );
and ( n1210 , n1209 , n1148 );
xor ( n1211 , n1149 , n1164 );
and ( n1212 , n1211 , n946 );
or ( n1213 , n1210 , n1212 );
not ( n1214 , n1213 );
not ( n1215 , n1214 );
not ( n1216 , n1215 );
not ( n1217 , n946 );
and ( n1218 , n1217 , n1154 );
xor ( n1219 , n1155 , n1163 );
and ( n1220 , n1219 , n946 );
or ( n1221 , n1218 , n1220 );
not ( n1222 , n1221 );
not ( n1223 , n1222 );
not ( n1224 , n1223 );
not ( n1225 , n946 );
and ( n1226 , n1225 , n1160 );
xor ( n1227 , n1161 , n1162 );
and ( n1228 , n1227 , n946 );
or ( n1229 , n1226 , n1228 );
not ( n1230 , n1229 );
not ( n1231 , n1230 );
not ( n1232 , n1231 );
not ( n1233 , n1114 );
and ( n1234 , n1232 , n1233 );
and ( n1235 , n1224 , n1234 );
and ( n1236 , n1216 , n1235 );
and ( n1237 , n1208 , n1236 );
and ( n1238 , n1200 , n1237 );
and ( n1239 , n1192 , n1238 );
and ( n1240 , n1184 , n1239 );
and ( n1241 , n1176 , n1240 );
not ( n1242 , n1241 );
and ( n1243 , n1242 , n946 );
buf ( n1244 , n1243 );
and ( n1245 , n1118 , n1244 );
not ( n1246 , n1245 );
and ( n1247 , n1246 , n1116 );
xor ( n1248 , n1116 , n1244 );
xor ( n1249 , n1248 , n1244 );
and ( n1250 , n1249 , n1245 );
or ( n1251 , n1247 , n1250 );
not ( n1252 , n946 );
and ( n1253 , n1252 , n1160 );
not ( n1254 , n1160 );
not ( n1255 , n952 );
not ( n1256 , n959 );
not ( n1257 , n965 );
not ( n1258 , n971 );
not ( n1259 , n977 );
not ( n1260 , n983 );
not ( n1261 , n989 );
not ( n1262 , n995 );
not ( n1263 , n1001 );
not ( n1264 , n1007 );
not ( n1265 , n1013 );
not ( n1266 , n1019 );
not ( n1267 , n1025 );
not ( n1268 , n1031 );
not ( n1269 , n1037 );
not ( n1270 , n1043 );
not ( n1271 , n1049 );
not ( n1272 , n1055 );
not ( n1273 , n1061 );
not ( n1274 , n1067 );
not ( n1275 , n1073 );
not ( n1276 , n1079 );
not ( n1277 , n1085 );
not ( n1278 , n911 );
and ( n1279 , n1277 , n1278 );
and ( n1280 , n1276 , n1279 );
and ( n1281 , n1275 , n1280 );
and ( n1282 , n1274 , n1281 );
and ( n1283 , n1273 , n1282 );
and ( n1284 , n1272 , n1283 );
and ( n1285 , n1271 , n1284 );
and ( n1286 , n1270 , n1285 );
and ( n1287 , n1269 , n1286 );
and ( n1288 , n1268 , n1287 );
and ( n1289 , n1267 , n1288 );
and ( n1290 , n1266 , n1289 );
and ( n1291 , n1265 , n1290 );
and ( n1292 , n1264 , n1291 );
and ( n1293 , n1263 , n1292 );
and ( n1294 , n1262 , n1293 );
and ( n1295 , n1261 , n1294 );
and ( n1296 , n1260 , n1295 );
and ( n1297 , n1259 , n1296 );
and ( n1298 , n1258 , n1297 );
and ( n1299 , n1257 , n1298 );
and ( n1300 , n1256 , n1299 );
and ( n1301 , n1255 , n1300 );
xor ( n1302 , n1254 , n1301 );
and ( n1303 , n1302 , n946 );
or ( n1304 , n1253 , n1303 );
not ( n1305 , n1304 );
not ( n1306 , n1305 );
not ( n1307 , n1306 );
not ( n1308 , n1307 );
not ( n1309 , n946 );
not ( n1310 , n1124 );
not ( n1311 , n1130 );
not ( n1312 , n1136 );
not ( n1313 , n1142 );
not ( n1314 , n1148 );
not ( n1315 , n1154 );
and ( n1316 , n1254 , n1301 );
and ( n1317 , n1315 , n1316 );
and ( n1318 , n1314 , n1317 );
and ( n1319 , n1313 , n1318 );
and ( n1320 , n1312 , n1319 );
and ( n1321 , n1311 , n1320 );
and ( n1322 , n1310 , n1321 );
xor ( n1323 , n1309 , n1322 );
buf ( n1324 , n946 );
and ( n1325 , n1323 , n1324 );
buf ( n1326 , n1325 );
not ( n1327 , n1326 );
not ( n1328 , n1327 );
not ( n1329 , n1328 );
not ( n1330 , n946 );
and ( n1331 , n1330 , n1124 );
xor ( n1332 , n1310 , n1321 );
and ( n1333 , n1332 , n946 );
or ( n1334 , n1331 , n1333 );
not ( n1335 , n1334 );
not ( n1336 , n1335 );
not ( n1337 , n1336 );
not ( n1338 , n946 );
and ( n1339 , n1338 , n1130 );
xor ( n1340 , n1311 , n1320 );
and ( n1341 , n1340 , n946 );
or ( n1342 , n1339 , n1341 );
not ( n1343 , n1342 );
not ( n1344 , n1343 );
not ( n1345 , n1344 );
not ( n1346 , n946 );
and ( n1347 , n1346 , n1136 );
xor ( n1348 , n1312 , n1319 );
and ( n1349 , n1348 , n946 );
or ( n1350 , n1347 , n1349 );
not ( n1351 , n1350 );
not ( n1352 , n1351 );
not ( n1353 , n1352 );
not ( n1354 , n946 );
and ( n1355 , n1354 , n1142 );
xor ( n1356 , n1313 , n1318 );
and ( n1357 , n1356 , n946 );
or ( n1358 , n1355 , n1357 );
not ( n1359 , n1358 );
not ( n1360 , n1359 );
not ( n1361 , n1360 );
not ( n1362 , n946 );
and ( n1363 , n1362 , n1148 );
xor ( n1364 , n1314 , n1317 );
and ( n1365 , n1364 , n946 );
or ( n1366 , n1363 , n1365 );
not ( n1367 , n1366 );
not ( n1368 , n1367 );
not ( n1369 , n1368 );
not ( n1370 , n946 );
and ( n1371 , n1370 , n1154 );
xor ( n1372 , n1315 , n1316 );
and ( n1373 , n1372 , n946 );
or ( n1374 , n1371 , n1373 );
not ( n1375 , n1374 );
not ( n1376 , n1375 );
not ( n1377 , n1376 );
not ( n1378 , n1306 );
and ( n1379 , n1377 , n1378 );
and ( n1380 , n1369 , n1379 );
and ( n1381 , n1361 , n1380 );
and ( n1382 , n1353 , n1381 );
and ( n1383 , n1345 , n1382 );
and ( n1384 , n1337 , n1383 );
and ( n1385 , n1329 , n1384 );
not ( n1386 , n1385 );
and ( n1387 , n1386 , n946 );
buf ( n1388 , n1387 );
not ( n1389 , n1388 );
not ( n1390 , n946 );
and ( n1391 , n1390 , n1376 );
xor ( n1392 , n1377 , n1378 );
and ( n1393 , n1392 , n946 );
or ( n1394 , n1391 , n1393 );
and ( n1395 , n1389 , n1394 );
not ( n1396 , n1394 );
not ( n1397 , n1306 );
xor ( n1398 , n1396 , n1397 );
and ( n1399 , n1398 , n1388 );
or ( n1400 , n1395 , n1399 );
not ( n1401 , n1400 );
not ( n1402 , n1401 );
or ( n1403 , n1308 , n1402 );
not ( n1404 , n1388 );
not ( n1405 , n946 );
and ( n1406 , n1405 , n1368 );
xor ( n1407 , n1369 , n1379 );
and ( n1408 , n1407 , n946 );
or ( n1409 , n1406 , n1408 );
and ( n1410 , n1404 , n1409 );
not ( n1411 , n1409 );
and ( n1412 , n1396 , n1397 );
xor ( n1413 , n1411 , n1412 );
and ( n1414 , n1413 , n1388 );
or ( n1415 , n1410 , n1414 );
not ( n1416 , n1415 );
not ( n1417 , n1416 );
or ( n1418 , n1403 , n1417 );
and ( n1419 , n1418 , n1388 );
not ( n1420 , n1419 );
and ( n1421 , n1420 , n1308 );
xor ( n1422 , n1308 , n1388 );
xor ( n1423 , n1422 , n1388 );
and ( n1424 , n1423 , n1419 );
or ( n1425 , n1421 , n1424 );
not ( n1426 , n1419 );
and ( n1427 , n1426 , n1402 );
xor ( n1428 , n1402 , n1388 );
and ( n1429 , n1422 , n1388 );
xor ( n1430 , n1428 , n1429 );
and ( n1431 , n1430 , n1419 );
or ( n1432 , n1427 , n1431 );
not ( n1433 , n1419 );
and ( n1434 , n1433 , n1417 );
xor ( n1435 , n1417 , n1388 );
and ( n1436 , n1428 , n1429 );
xor ( n1437 , n1435 , n1436 );
and ( n1438 , n1437 , n1419 );
or ( n1439 , n1434 , n1438 );
and ( n1440 , n1425 , n1432 , n1439 );
or ( n1441 , n1251 , n1440 );
not ( n1442 , n1441 );
buf ( n1443 , n722 );
buf ( n1444 , n1443 );
not ( n1445 , n1444 );
not ( n1446 , n1445 );
buf ( n1447 , n1446 );
not ( n1448 , n946 );
and ( n1449 , n1448 , n977 );
not ( n1450 , n977 );
not ( n1451 , n983 );
not ( n1452 , n989 );
not ( n1453 , n995 );
not ( n1454 , n1001 );
not ( n1455 , n1007 );
not ( n1456 , n1013 );
not ( n1457 , n1019 );
not ( n1458 , n1025 );
not ( n1459 , n1031 );
not ( n1460 , n1037 );
not ( n1461 , n1043 );
not ( n1462 , n1049 );
not ( n1463 , n1055 );
not ( n1464 , n1061 );
not ( n1465 , n1067 );
not ( n1466 , n1073 );
not ( n1467 , n1079 );
not ( n1468 , n1085 );
not ( n1469 , n911 );
and ( n1470 , n1468 , n1469 );
and ( n1471 , n1467 , n1470 );
and ( n1472 , n1466 , n1471 );
and ( n1473 , n1465 , n1472 );
and ( n1474 , n1464 , n1473 );
and ( n1475 , n1463 , n1474 );
and ( n1476 , n1462 , n1475 );
and ( n1477 , n1461 , n1476 );
and ( n1478 , n1460 , n1477 );
and ( n1479 , n1459 , n1478 );
and ( n1480 , n1458 , n1479 );
and ( n1481 , n1457 , n1480 );
and ( n1482 , n1456 , n1481 );
and ( n1483 , n1455 , n1482 );
and ( n1484 , n1454 , n1483 );
and ( n1485 , n1453 , n1484 );
and ( n1486 , n1452 , n1485 );
and ( n1487 , n1451 , n1486 );
xor ( n1488 , n1450 , n1487 );
and ( n1489 , n1488 , n946 );
or ( n1490 , n1449 , n1489 );
not ( n1491 , n1490 );
not ( n1492 , n1491 );
not ( n1493 , n1492 );
not ( n1494 , n1493 );
not ( n1495 , n946 );
not ( n1496 , n1124 );
not ( n1497 , n1130 );
not ( n1498 , n1136 );
not ( n1499 , n1142 );
not ( n1500 , n1148 );
not ( n1501 , n1154 );
not ( n1502 , n1160 );
not ( n1503 , n952 );
not ( n1504 , n959 );
not ( n1505 , n965 );
not ( n1506 , n971 );
and ( n1507 , n1450 , n1487 );
and ( n1508 , n1506 , n1507 );
and ( n1509 , n1505 , n1508 );
and ( n1510 , n1504 , n1509 );
and ( n1511 , n1503 , n1510 );
and ( n1512 , n1502 , n1511 );
and ( n1513 , n1501 , n1512 );
and ( n1514 , n1500 , n1513 );
and ( n1515 , n1499 , n1514 );
and ( n1516 , n1498 , n1515 );
and ( n1517 , n1497 , n1516 );
and ( n1518 , n1496 , n1517 );
xor ( n1519 , n1495 , n1518 );
buf ( n1520 , n946 );
and ( n1521 , n1519 , n1520 );
buf ( n1522 , n1521 );
not ( n1523 , n1522 );
not ( n1524 , n1523 );
not ( n1525 , n1524 );
not ( n1526 , n946 );
and ( n1527 , n1526 , n1124 );
xor ( n1528 , n1496 , n1517 );
and ( n1529 , n1528 , n946 );
or ( n1530 , n1527 , n1529 );
not ( n1531 , n1530 );
not ( n1532 , n1531 );
not ( n1533 , n1532 );
not ( n1534 , n946 );
and ( n1535 , n1534 , n1130 );
xor ( n1536 , n1497 , n1516 );
and ( n1537 , n1536 , n946 );
or ( n1538 , n1535 , n1537 );
not ( n1539 , n1538 );
not ( n1540 , n1539 );
not ( n1541 , n1540 );
not ( n1542 , n946 );
and ( n1543 , n1542 , n1136 );
xor ( n1544 , n1498 , n1515 );
and ( n1545 , n1544 , n946 );
or ( n1546 , n1543 , n1545 );
not ( n1547 , n1546 );
not ( n1548 , n1547 );
not ( n1549 , n1548 );
not ( n1550 , n946 );
and ( n1551 , n1550 , n1142 );
xor ( n1552 , n1499 , n1514 );
and ( n1553 , n1552 , n946 );
or ( n1554 , n1551 , n1553 );
not ( n1555 , n1554 );
not ( n1556 , n1555 );
not ( n1557 , n1556 );
not ( n1558 , n946 );
and ( n1559 , n1558 , n1148 );
xor ( n1560 , n1500 , n1513 );
and ( n1561 , n1560 , n946 );
or ( n1562 , n1559 , n1561 );
not ( n1563 , n1562 );
not ( n1564 , n1563 );
not ( n1565 , n1564 );
not ( n1566 , n946 );
and ( n1567 , n1566 , n1154 );
xor ( n1568 , n1501 , n1512 );
and ( n1569 , n1568 , n946 );
or ( n1570 , n1567 , n1569 );
not ( n1571 , n1570 );
not ( n1572 , n1571 );
not ( n1573 , n1572 );
not ( n1574 , n946 );
and ( n1575 , n1574 , n1160 );
xor ( n1576 , n1502 , n1511 );
and ( n1577 , n1576 , n946 );
or ( n1578 , n1575 , n1577 );
not ( n1579 , n1578 );
not ( n1580 , n1579 );
not ( n1581 , n1580 );
not ( n1582 , n946 );
and ( n1583 , n1582 , n952 );
xor ( n1584 , n1503 , n1510 );
and ( n1585 , n1584 , n946 );
or ( n1586 , n1583 , n1585 );
not ( n1587 , n1586 );
not ( n1588 , n1587 );
not ( n1589 , n1588 );
not ( n1590 , n946 );
and ( n1591 , n1590 , n959 );
xor ( n1592 , n1504 , n1509 );
and ( n1593 , n1592 , n946 );
or ( n1594 , n1591 , n1593 );
not ( n1595 , n1594 );
not ( n1596 , n1595 );
not ( n1597 , n1596 );
not ( n1598 , n946 );
and ( n1599 , n1598 , n965 );
xor ( n1600 , n1505 , n1508 );
and ( n1601 , n1600 , n946 );
or ( n1602 , n1599 , n1601 );
not ( n1603 , n1602 );
not ( n1604 , n1603 );
not ( n1605 , n1604 );
not ( n1606 , n946 );
and ( n1607 , n1606 , n971 );
xor ( n1608 , n1506 , n1507 );
and ( n1609 , n1608 , n946 );
or ( n1610 , n1607 , n1609 );
not ( n1611 , n1610 );
not ( n1612 , n1611 );
not ( n1613 , n1612 );
not ( n1614 , n1492 );
and ( n1615 , n1613 , n1614 );
and ( n1616 , n1605 , n1615 );
and ( n1617 , n1597 , n1616 );
and ( n1618 , n1589 , n1617 );
and ( n1619 , n1581 , n1618 );
and ( n1620 , n1573 , n1619 );
and ( n1621 , n1565 , n1620 );
and ( n1622 , n1557 , n1621 );
and ( n1623 , n1549 , n1622 );
and ( n1624 , n1541 , n1623 );
and ( n1625 , n1533 , n1624 );
and ( n1626 , n1525 , n1625 );
not ( n1627 , n1626 );
and ( n1628 , n1627 , n946 );
buf ( n1629 , n1628 );
not ( n1630 , n1629 );
not ( n1631 , n946 );
and ( n1632 , n1631 , n1612 );
xor ( n1633 , n1613 , n1614 );
and ( n1634 , n1633 , n946 );
or ( n1635 , n1632 , n1634 );
and ( n1636 , n1630 , n1635 );
not ( n1637 , n1635 );
not ( n1638 , n1492 );
xor ( n1639 , n1637 , n1638 );
and ( n1640 , n1639 , n1629 );
or ( n1641 , n1636 , n1640 );
not ( n1642 , n1641 );
not ( n1643 , n1642 );
or ( n1644 , n1494 , n1643 );
not ( n1645 , n1629 );
not ( n1646 , n946 );
and ( n1647 , n1646 , n1604 );
xor ( n1648 , n1605 , n1615 );
and ( n1649 , n1648 , n946 );
or ( n1650 , n1647 , n1649 );
and ( n1651 , n1645 , n1650 );
not ( n1652 , n1650 );
and ( n1653 , n1637 , n1638 );
xor ( n1654 , n1652 , n1653 );
and ( n1655 , n1654 , n1629 );
or ( n1656 , n1651 , n1655 );
not ( n1657 , n1656 );
not ( n1658 , n1657 );
or ( n1659 , n1644 , n1658 );
not ( n1660 , n1629 );
not ( n1661 , n946 );
and ( n1662 , n1661 , n1596 );
xor ( n1663 , n1597 , n1616 );
and ( n1664 , n1663 , n946 );
or ( n1665 , n1662 , n1664 );
and ( n1666 , n1660 , n1665 );
not ( n1667 , n1665 );
and ( n1668 , n1652 , n1653 );
xor ( n1669 , n1667 , n1668 );
and ( n1670 , n1669 , n1629 );
or ( n1671 , n1666 , n1670 );
not ( n1672 , n1671 );
not ( n1673 , n1672 );
or ( n1674 , n1659 , n1673 );
buf ( n1675 , n1674 );
buf ( n1676 , n1675 );
and ( n1677 , n1676 , n1629 );
not ( n1678 , n1677 );
and ( n1679 , n1678 , n1494 );
xor ( n1680 , n1494 , n1629 );
xor ( n1681 , n1680 , n1629 );
and ( n1682 , n1681 , n1677 );
or ( n1683 , n1679 , n1682 );
not ( n1684 , n1677 );
and ( n1685 , n1684 , n1643 );
xor ( n1686 , n1643 , n1629 );
and ( n1687 , n1680 , n1629 );
xor ( n1688 , n1686 , n1687 );
and ( n1689 , n1688 , n1677 );
or ( n1690 , n1685 , n1689 );
not ( n1691 , n1690 );
not ( n1692 , n1677 );
and ( n1693 , n1692 , n1658 );
xor ( n1694 , n1658 , n1629 );
and ( n1695 , n1686 , n1687 );
xor ( n1696 , n1694 , n1695 );
and ( n1697 , n1696 , n1677 );
or ( n1698 , n1693 , n1697 );
not ( n1699 , n1677 );
and ( n1700 , n1699 , n1673 );
xor ( n1701 , n1673 , n1629 );
and ( n1702 , n1694 , n1695 );
xor ( n1703 , n1701 , n1702 );
and ( n1704 , n1703 , n1677 );
or ( n1705 , n1700 , n1704 );
and ( n1706 , n1683 , n1691 , n1698 , n1705 );
not ( n1707 , n1683 );
and ( n1708 , n1707 , n1690 , n1698 , n1705 );
or ( n1709 , n1706 , n1708 );
and ( n1710 , n1683 , n1690 , n1698 , n1705 );
or ( n1711 , n1709 , n1710 );
and ( n1712 , n1447 , n1711 );
buf ( n1713 , n721 );
not ( n1714 , n1713 );
not ( n1715 , n1714 );
buf ( n1716 , n1715 );
not ( n1717 , n946 );
and ( n1718 , n1717 , n1130 );
not ( n1719 , n1130 );
not ( n1720 , n1136 );
not ( n1721 , n1142 );
not ( n1722 , n1148 );
not ( n1723 , n1154 );
not ( n1724 , n1160 );
not ( n1725 , n952 );
not ( n1726 , n959 );
not ( n1727 , n965 );
not ( n1728 , n971 );
not ( n1729 , n977 );
not ( n1730 , n983 );
not ( n1731 , n989 );
not ( n1732 , n995 );
not ( n1733 , n1001 );
not ( n1734 , n1007 );
not ( n1735 , n1013 );
not ( n1736 , n1019 );
not ( n1737 , n1025 );
not ( n1738 , n1031 );
not ( n1739 , n1037 );
not ( n1740 , n1043 );
not ( n1741 , n1049 );
not ( n1742 , n1055 );
not ( n1743 , n1061 );
not ( n1744 , n1067 );
not ( n1745 , n1073 );
not ( n1746 , n1079 );
not ( n1747 , n1085 );
not ( n1748 , n911 );
and ( n1749 , n1747 , n1748 );
and ( n1750 , n1746 , n1749 );
and ( n1751 , n1745 , n1750 );
and ( n1752 , n1744 , n1751 );
and ( n1753 , n1743 , n1752 );
and ( n1754 , n1742 , n1753 );
and ( n1755 , n1741 , n1754 );
and ( n1756 , n1740 , n1755 );
and ( n1757 , n1739 , n1756 );
and ( n1758 , n1738 , n1757 );
and ( n1759 , n1737 , n1758 );
and ( n1760 , n1736 , n1759 );
and ( n1761 , n1735 , n1760 );
and ( n1762 , n1734 , n1761 );
and ( n1763 , n1733 , n1762 );
and ( n1764 , n1732 , n1763 );
and ( n1765 , n1731 , n1764 );
and ( n1766 , n1730 , n1765 );
and ( n1767 , n1729 , n1766 );
and ( n1768 , n1728 , n1767 );
and ( n1769 , n1727 , n1768 );
and ( n1770 , n1726 , n1769 );
and ( n1771 , n1725 , n1770 );
and ( n1772 , n1724 , n1771 );
and ( n1773 , n1723 , n1772 );
and ( n1774 , n1722 , n1773 );
and ( n1775 , n1721 , n1774 );
and ( n1776 , n1720 , n1775 );
xor ( n1777 , n1719 , n1776 );
and ( n1778 , n1777 , n946 );
or ( n1779 , n1718 , n1778 );
not ( n1780 , n1779 );
not ( n1781 , n1780 );
not ( n1782 , n1781 );
not ( n1783 , n1782 );
not ( n1784 , n946 );
not ( n1785 , n1124 );
and ( n1786 , n1719 , n1776 );
and ( n1787 , n1785 , n1786 );
xor ( n1788 , n1784 , n1787 );
buf ( n1789 , n946 );
and ( n1790 , n1788 , n1789 );
buf ( n1791 , n1790 );
not ( n1792 , n1791 );
not ( n1793 , n1792 );
not ( n1794 , n1793 );
not ( n1795 , n946 );
and ( n1796 , n1795 , n1124 );
xor ( n1797 , n1785 , n1786 );
and ( n1798 , n1797 , n946 );
or ( n1799 , n1796 , n1798 );
not ( n1800 , n1799 );
not ( n1801 , n1800 );
not ( n1802 , n1801 );
not ( n1803 , n1781 );
and ( n1804 , n1802 , n1803 );
and ( n1805 , n1794 , n1804 );
not ( n1806 , n1805 );
and ( n1807 , n1806 , n946 );
buf ( n1808 , n1807 );
not ( n1809 , n1808 );
not ( n1810 , n946 );
and ( n1811 , n1810 , n1801 );
xor ( n1812 , n1802 , n1803 );
and ( n1813 , n1812 , n946 );
or ( n1814 , n1811 , n1813 );
and ( n1815 , n1809 , n1814 );
not ( n1816 , n1814 );
not ( n1817 , n1781 );
xor ( n1818 , n1816 , n1817 );
and ( n1819 , n1818 , n1808 );
or ( n1820 , n1815 , n1819 );
not ( n1821 , n1820 );
not ( n1822 , n1821 );
or ( n1823 , n1783 , n1822 );
and ( n1824 , n1823 , n1808 );
not ( n1825 , n1824 );
and ( n1826 , n1825 , n1783 );
xor ( n1827 , n1783 , n1808 );
xor ( n1828 , n1827 , n1808 );
and ( n1829 , n1828 , n1824 );
or ( n1830 , n1826 , n1829 );
not ( n1831 , n1824 );
and ( n1832 , n1831 , n1822 );
xor ( n1833 , n1822 , n1808 );
and ( n1834 , n1827 , n1808 );
xor ( n1835 , n1833 , n1834 );
and ( n1836 , n1835 , n1824 );
or ( n1837 , n1832 , n1836 );
and ( n1838 , n1830 , n1837 );
and ( n1839 , n1716 , n1838 );
buf ( n1840 , n815 );
not ( n1841 , n1830 );
and ( n1842 , n1841 , n1837 );
and ( n1843 , n1840 , n1842 );
buf ( n1844 , n750 );
nor ( n1845 , n1841 , n1837 );
and ( n1846 , n1844 , n1845 );
buf ( n1847 , n782 );
nor ( n1848 , n1830 , n1837 );
and ( n1849 , n1847 , n1848 );
or ( n1850 , n1839 , n1843 , n1846 , n1849 );
not ( n1851 , n1850 );
not ( n1852 , n1851 );
buf ( n1853 , n846 );
and ( n1854 , n1853 , n1842 );
buf ( n1855 , n781 );
and ( n1856 , n1855 , n1845 );
buf ( n1857 , n813 );
and ( n1858 , n1857 , n1848 );
or ( n1859 , 1'b0 , n1854 , n1856 , n1858 );
not ( n1860 , n1859 );
and ( n1861 , n1447 , n1838 );
buf ( n1862 , n816 );
and ( n1863 , n1862 , n1842 );
buf ( n1864 , n751 );
and ( n1865 , n1864 , n1845 );
buf ( n1866 , n783 );
and ( n1867 , n1866 , n1848 );
or ( n1868 , n1861 , n1863 , n1865 , n1867 );
and ( n1869 , n1860 , n1868 );
not ( n1870 , n1868 );
not ( n1871 , n1850 );
xor ( n1872 , n1870 , n1871 );
and ( n1873 , n1872 , n1859 );
or ( n1874 , n1869 , n1873 );
not ( n1875 , n1874 );
not ( n1876 , n1875 );
or ( n1877 , n1852 , n1876 );
not ( n1878 , n1859 );
buf ( n1879 , n723 );
buf ( n1880 , n1879 );
not ( n1881 , n1880 );
not ( n1882 , n1881 );
buf ( n1883 , n1882 );
and ( n1884 , n1883 , n1838 );
buf ( n1885 , n817 );
and ( n1886 , n1885 , n1842 );
buf ( n1887 , n752 );
and ( n1888 , n1887 , n1845 );
buf ( n1889 , n784 );
and ( n1890 , n1889 , n1848 );
or ( n1891 , n1884 , n1886 , n1888 , n1890 );
and ( n1892 , n1878 , n1891 );
not ( n1893 , n1891 );
and ( n1894 , n1870 , n1871 );
xor ( n1895 , n1893 , n1894 );
and ( n1896 , n1895 , n1859 );
or ( n1897 , n1892 , n1896 );
not ( n1898 , n1897 );
not ( n1899 , n1898 );
or ( n1900 , n1877 , n1899 );
not ( n1901 , n1859 );
buf ( n1902 , n724 );
buf ( n1903 , n1902 );
not ( n1904 , n1903 );
not ( n1905 , n1904 );
buf ( n1906 , n1905 );
not ( n1907 , n1906 );
and ( n1908 , n1907 , n1838 );
buf ( n1909 , n818 );
and ( n1910 , n1909 , n1842 );
buf ( n1911 , n753 );
and ( n1912 , n1911 , n1845 );
buf ( n1913 , n785 );
and ( n1914 , n1913 , n1848 );
or ( n1915 , n1908 , n1910 , n1912 , n1914 );
and ( n1916 , n1901 , n1915 );
not ( n1917 , n1915 );
and ( n1918 , n1893 , n1894 );
xor ( n1919 , n1917 , n1918 );
and ( n1920 , n1919 , n1859 );
or ( n1921 , n1916 , n1920 );
not ( n1922 , n1921 );
not ( n1923 , n1922 );
or ( n1924 , n1900 , n1923 );
not ( n1925 , n1859 );
buf ( n1926 , n725 );
buf ( n1927 , n1926 );
not ( n1928 , n1927 );
not ( n1929 , n1928 );
buf ( n1930 , n1929 );
xor ( n1931 , n1930 , n1906 );
and ( n1932 , n1931 , n1838 );
buf ( n1933 , n819 );
and ( n1934 , n1933 , n1842 );
buf ( n1935 , n754 );
and ( n1936 , n1935 , n1845 );
buf ( n1937 , n786 );
and ( n1938 , n1937 , n1848 );
or ( n1939 , n1932 , n1934 , n1936 , n1938 );
and ( n1940 , n1925 , n1939 );
not ( n1941 , n1939 );
and ( n1942 , n1917 , n1918 );
xor ( n1943 , n1941 , n1942 );
and ( n1944 , n1943 , n1859 );
or ( n1945 , n1940 , n1944 );
not ( n1946 , n1945 );
not ( n1947 , n1946 );
or ( n1948 , n1924 , n1947 );
not ( n1949 , n1859 );
buf ( n1950 , n726 );
not ( n1951 , n1950 );
not ( n1952 , n1951 );
buf ( n1953 , n1952 );
and ( n1954 , n1930 , n1906 );
xor ( n1955 , n1953 , n1954 );
and ( n1956 , n1955 , n1838 );
buf ( n1957 , n820 );
and ( n1958 , n1957 , n1842 );
buf ( n1959 , n755 );
and ( n1960 , n1959 , n1845 );
buf ( n1961 , n787 );
and ( n1962 , n1961 , n1848 );
or ( n1963 , n1956 , n1958 , n1960 , n1962 );
and ( n1964 , n1949 , n1963 );
not ( n1965 , n1963 );
and ( n1966 , n1941 , n1942 );
xor ( n1967 , n1965 , n1966 );
and ( n1968 , n1967 , n1859 );
or ( n1969 , n1964 , n1968 );
not ( n1970 , n1969 );
not ( n1971 , n1970 );
or ( n1972 , n1948 , n1971 );
not ( n1973 , n1859 );
buf ( n1974 , n727 );
not ( n1975 , n1974 );
not ( n1976 , n1975 );
buf ( n1977 , n1976 );
and ( n1978 , n1953 , n1954 );
xor ( n1979 , n1977 , n1978 );
and ( n1980 , n1979 , n1838 );
buf ( n1981 , n821 );
and ( n1982 , n1981 , n1842 );
buf ( n1983 , n756 );
and ( n1984 , n1983 , n1845 );
buf ( n1985 , n788 );
and ( n1986 , n1985 , n1848 );
or ( n1987 , n1980 , n1982 , n1984 , n1986 );
and ( n1988 , n1973 , n1987 );
not ( n1989 , n1987 );
and ( n1990 , n1965 , n1966 );
xor ( n1991 , n1989 , n1990 );
and ( n1992 , n1991 , n1859 );
or ( n1993 , n1988 , n1992 );
not ( n1994 , n1993 );
not ( n1995 , n1994 );
or ( n1996 , n1972 , n1995 );
not ( n1997 , n1859 );
buf ( n1998 , n728 );
not ( n1999 , n1998 );
not ( n2000 , n1999 );
buf ( n2001 , n2000 );
and ( n2002 , n1977 , n1978 );
xor ( n2003 , n2001 , n2002 );
and ( n2004 , n2003 , n1838 );
buf ( n2005 , n822 );
and ( n2006 , n2005 , n1842 );
buf ( n2007 , n757 );
and ( n2008 , n2007 , n1845 );
buf ( n2009 , n789 );
and ( n2010 , n2009 , n1848 );
or ( n2011 , n2004 , n2006 , n2008 , n2010 );
and ( n2012 , n1997 , n2011 );
not ( n2013 , n2011 );
and ( n2014 , n1989 , n1990 );
xor ( n2015 , n2013 , n2014 );
and ( n2016 , n2015 , n1859 );
or ( n2017 , n2012 , n2016 );
not ( n2018 , n2017 );
not ( n2019 , n2018 );
or ( n2020 , n1996 , n2019 );
not ( n2021 , n1859 );
buf ( n2022 , n729 );
not ( n2023 , n2022 );
not ( n2024 , n2023 );
buf ( n2025 , n2024 );
and ( n2026 , n2001 , n2002 );
xor ( n2027 , n2025 , n2026 );
and ( n2028 , n2027 , n1838 );
buf ( n2029 , n823 );
and ( n2030 , n2029 , n1842 );
buf ( n2031 , n758 );
and ( n2032 , n2031 , n1845 );
buf ( n2033 , n790 );
and ( n2034 , n2033 , n1848 );
or ( n2035 , n2028 , n2030 , n2032 , n2034 );
and ( n2036 , n2021 , n2035 );
not ( n2037 , n2035 );
and ( n2038 , n2013 , n2014 );
xor ( n2039 , n2037 , n2038 );
and ( n2040 , n2039 , n1859 );
or ( n2041 , n2036 , n2040 );
not ( n2042 , n2041 );
not ( n2043 , n2042 );
or ( n2044 , n2020 , n2043 );
not ( n2045 , n1859 );
buf ( n2046 , n730 );
not ( n2047 , n2046 );
not ( n2048 , n2047 );
buf ( n2049 , n2048 );
and ( n2050 , n2025 , n2026 );
xor ( n2051 , n2049 , n2050 );
and ( n2052 , n2051 , n1838 );
buf ( n2053 , n824 );
and ( n2054 , n2053 , n1842 );
buf ( n2055 , n759 );
and ( n2056 , n2055 , n1845 );
buf ( n2057 , n791 );
and ( n2058 , n2057 , n1848 );
or ( n2059 , n2052 , n2054 , n2056 , n2058 );
and ( n2060 , n2045 , n2059 );
not ( n2061 , n2059 );
and ( n2062 , n2037 , n2038 );
xor ( n2063 , n2061 , n2062 );
and ( n2064 , n2063 , n1859 );
or ( n2065 , n2060 , n2064 );
not ( n2066 , n2065 );
not ( n2067 , n2066 );
or ( n2068 , n2044 , n2067 );
not ( n2069 , n1859 );
buf ( n2070 , n731 );
not ( n2071 , n2070 );
not ( n2072 , n2071 );
buf ( n2073 , n2072 );
and ( n2074 , n2049 , n2050 );
xor ( n2075 , n2073 , n2074 );
and ( n2076 , n2075 , n1838 );
buf ( n2077 , n825 );
and ( n2078 , n2077 , n1842 );
buf ( n2079 , n760 );
and ( n2080 , n2079 , n1845 );
buf ( n2081 , n792 );
and ( n2082 , n2081 , n1848 );
or ( n2083 , n2076 , n2078 , n2080 , n2082 );
and ( n2084 , n2069 , n2083 );
not ( n2085 , n2083 );
and ( n2086 , n2061 , n2062 );
xor ( n2087 , n2085 , n2086 );
and ( n2088 , n2087 , n1859 );
or ( n2089 , n2084 , n2088 );
not ( n2090 , n2089 );
not ( n2091 , n2090 );
or ( n2092 , n2068 , n2091 );
not ( n2093 , n1859 );
buf ( n2094 , n732 );
not ( n2095 , n2094 );
not ( n2096 , n2095 );
buf ( n2097 , n2096 );
and ( n2098 , n2073 , n2074 );
xor ( n2099 , n2097 , n2098 );
and ( n2100 , n2099 , n1838 );
buf ( n2101 , n826 );
and ( n2102 , n2101 , n1842 );
buf ( n2103 , n761 );
and ( n2104 , n2103 , n1845 );
buf ( n2105 , n793 );
and ( n2106 , n2105 , n1848 );
or ( n2107 , n2100 , n2102 , n2104 , n2106 );
and ( n2108 , n2093 , n2107 );
not ( n2109 , n2107 );
and ( n2110 , n2085 , n2086 );
xor ( n2111 , n2109 , n2110 );
and ( n2112 , n2111 , n1859 );
or ( n2113 , n2108 , n2112 );
not ( n2114 , n2113 );
not ( n2115 , n2114 );
or ( n2116 , n2092 , n2115 );
not ( n2117 , n1859 );
buf ( n2118 , n733 );
not ( n2119 , n2118 );
not ( n2120 , n2119 );
buf ( n2121 , n2120 );
and ( n2122 , n2097 , n2098 );
xor ( n2123 , n2121 , n2122 );
and ( n2124 , n2123 , n1838 );
buf ( n2125 , n827 );
and ( n2126 , n2125 , n1842 );
buf ( n2127 , n762 );
and ( n2128 , n2127 , n1845 );
buf ( n2129 , n794 );
and ( n2130 , n2129 , n1848 );
or ( n2131 , n2124 , n2126 , n2128 , n2130 );
and ( n2132 , n2117 , n2131 );
not ( n2133 , n2131 );
and ( n2134 , n2109 , n2110 );
xor ( n2135 , n2133 , n2134 );
and ( n2136 , n2135 , n1859 );
or ( n2137 , n2132 , n2136 );
not ( n2138 , n2137 );
not ( n2139 , n2138 );
or ( n2140 , n2116 , n2139 );
not ( n2141 , n1859 );
buf ( n2142 , n734 );
not ( n2143 , n2142 );
not ( n2144 , n2143 );
buf ( n2145 , n2144 );
and ( n2146 , n2121 , n2122 );
xor ( n2147 , n2145 , n2146 );
and ( n2148 , n2147 , n1838 );
buf ( n2149 , n828 );
and ( n2150 , n2149 , n1842 );
buf ( n2151 , n763 );
and ( n2152 , n2151 , n1845 );
buf ( n2153 , n795 );
and ( n2154 , n2153 , n1848 );
or ( n2155 , n2148 , n2150 , n2152 , n2154 );
and ( n2156 , n2141 , n2155 );
not ( n2157 , n2155 );
and ( n2158 , n2133 , n2134 );
xor ( n2159 , n2157 , n2158 );
and ( n2160 , n2159 , n1859 );
or ( n2161 , n2156 , n2160 );
not ( n2162 , n2161 );
not ( n2163 , n2162 );
or ( n2164 , n2140 , n2163 );
not ( n2165 , n1859 );
buf ( n2166 , n735 );
not ( n2167 , n2166 );
not ( n2168 , n2167 );
buf ( n2169 , n2168 );
and ( n2170 , n2145 , n2146 );
xor ( n2171 , n2169 , n2170 );
and ( n2172 , n2171 , n1838 );
buf ( n2173 , n829 );
and ( n2174 , n2173 , n1842 );
buf ( n2175 , n764 );
and ( n2176 , n2175 , n1845 );
buf ( n2177 , n796 );
and ( n2178 , n2177 , n1848 );
or ( n2179 , n2172 , n2174 , n2176 , n2178 );
and ( n2180 , n2165 , n2179 );
not ( n2181 , n2179 );
and ( n2182 , n2157 , n2158 );
xor ( n2183 , n2181 , n2182 );
and ( n2184 , n2183 , n1859 );
or ( n2185 , n2180 , n2184 );
not ( n2186 , n2185 );
not ( n2187 , n2186 );
or ( n2188 , n2164 , n2187 );
not ( n2189 , n1859 );
buf ( n2190 , n736 );
not ( n2191 , n2190 );
not ( n2192 , n2191 );
buf ( n2193 , n2192 );
and ( n2194 , n2169 , n2170 );
xor ( n2195 , n2193 , n2194 );
and ( n2196 , n2195 , n1838 );
buf ( n2197 , n830 );
and ( n2198 , n2197 , n1842 );
buf ( n2199 , n765 );
and ( n2200 , n2199 , n1845 );
buf ( n2201 , n797 );
and ( n2202 , n2201 , n1848 );
or ( n2203 , n2196 , n2198 , n2200 , n2202 );
and ( n2204 , n2189 , n2203 );
not ( n2205 , n2203 );
and ( n2206 , n2181 , n2182 );
xor ( n2207 , n2205 , n2206 );
and ( n2208 , n2207 , n1859 );
or ( n2209 , n2204 , n2208 );
not ( n2210 , n2209 );
not ( n2211 , n2210 );
or ( n2212 , n2188 , n2211 );
not ( n2213 , n1859 );
buf ( n2214 , n737 );
not ( n2215 , n2214 );
not ( n2216 , n2215 );
buf ( n2217 , n2216 );
and ( n2218 , n2193 , n2194 );
xor ( n2219 , n2217 , n2218 );
and ( n2220 , n2219 , n1838 );
buf ( n2221 , n831 );
and ( n2222 , n2221 , n1842 );
buf ( n2223 , n766 );
and ( n2224 , n2223 , n1845 );
buf ( n2225 , n798 );
and ( n2226 , n2225 , n1848 );
or ( n2227 , n2220 , n2222 , n2224 , n2226 );
and ( n2228 , n2213 , n2227 );
not ( n2229 , n2227 );
and ( n2230 , n2205 , n2206 );
xor ( n2231 , n2229 , n2230 );
and ( n2232 , n2231 , n1859 );
or ( n2233 , n2228 , n2232 );
not ( n2234 , n2233 );
not ( n2235 , n2234 );
or ( n2236 , n2212 , n2235 );
not ( n2237 , n1859 );
buf ( n2238 , n738 );
not ( n2239 , n2238 );
not ( n2240 , n2239 );
buf ( n2241 , n2240 );
and ( n2242 , n2217 , n2218 );
xor ( n2243 , n2241 , n2242 );
and ( n2244 , n2243 , n1838 );
buf ( n2245 , n832 );
and ( n2246 , n2245 , n1842 );
buf ( n2247 , n767 );
and ( n2248 , n2247 , n1845 );
buf ( n2249 , n799 );
and ( n2250 , n2249 , n1848 );
or ( n2251 , n2244 , n2246 , n2248 , n2250 );
and ( n2252 , n2237 , n2251 );
not ( n2253 , n2251 );
and ( n2254 , n2229 , n2230 );
xor ( n2255 , n2253 , n2254 );
and ( n2256 , n2255 , n1859 );
or ( n2257 , n2252 , n2256 );
not ( n2258 , n2257 );
not ( n2259 , n2258 );
or ( n2260 , n2236 , n2259 );
not ( n2261 , n1859 );
buf ( n2262 , n739 );
not ( n2263 , n2262 );
not ( n2264 , n2263 );
buf ( n2265 , n2264 );
and ( n2266 , n2241 , n2242 );
xor ( n2267 , n2265 , n2266 );
and ( n2268 , n2267 , n1838 );
buf ( n2269 , n833 );
and ( n2270 , n2269 , n1842 );
buf ( n2271 , n768 );
and ( n2272 , n2271 , n1845 );
buf ( n2273 , n800 );
and ( n2274 , n2273 , n1848 );
or ( n2275 , n2268 , n2270 , n2272 , n2274 );
and ( n2276 , n2261 , n2275 );
not ( n2277 , n2275 );
and ( n2278 , n2253 , n2254 );
xor ( n2279 , n2277 , n2278 );
and ( n2280 , n2279 , n1859 );
or ( n2281 , n2276 , n2280 );
not ( n2282 , n2281 );
not ( n2283 , n2282 );
or ( n2284 , n2260 , n2283 );
not ( n2285 , n1859 );
buf ( n2286 , n740 );
not ( n2287 , n2286 );
not ( n2288 , n2287 );
buf ( n2289 , n2288 );
and ( n2290 , n2265 , n2266 );
xor ( n2291 , n2289 , n2290 );
and ( n2292 , n2291 , n1838 );
buf ( n2293 , n834 );
and ( n2294 , n2293 , n1842 );
buf ( n2295 , n769 );
and ( n2296 , n2295 , n1845 );
buf ( n2297 , n801 );
and ( n2298 , n2297 , n1848 );
or ( n2299 , n2292 , n2294 , n2296 , n2298 );
and ( n2300 , n2285 , n2299 );
not ( n2301 , n2299 );
and ( n2302 , n2277 , n2278 );
xor ( n2303 , n2301 , n2302 );
and ( n2304 , n2303 , n1859 );
or ( n2305 , n2300 , n2304 );
not ( n2306 , n2305 );
not ( n2307 , n2306 );
or ( n2308 , n2284 , n2307 );
not ( n2309 , n1859 );
buf ( n2310 , n741 );
not ( n2311 , n2310 );
not ( n2312 , n2311 );
buf ( n2313 , n2312 );
and ( n2314 , n2289 , n2290 );
xor ( n2315 , n2313 , n2314 );
and ( n2316 , n2315 , n1838 );
buf ( n2317 , n835 );
and ( n2318 , n2317 , n1842 );
buf ( n2319 , n770 );
and ( n2320 , n2319 , n1845 );
buf ( n2321 , n802 );
and ( n2322 , n2321 , n1848 );
or ( n2323 , n2316 , n2318 , n2320 , n2322 );
and ( n2324 , n2309 , n2323 );
not ( n2325 , n2323 );
and ( n2326 , n2301 , n2302 );
xor ( n2327 , n2325 , n2326 );
and ( n2328 , n2327 , n1859 );
or ( n2329 , n2324 , n2328 );
not ( n2330 , n2329 );
not ( n2331 , n2330 );
or ( n2332 , n2308 , n2331 );
not ( n2333 , n1859 );
buf ( n2334 , n742 );
not ( n2335 , n2334 );
not ( n2336 , n2335 );
buf ( n2337 , n2336 );
and ( n2338 , n2313 , n2314 );
xor ( n2339 , n2337 , n2338 );
and ( n2340 , n2339 , n1838 );
buf ( n2341 , n836 );
and ( n2342 , n2341 , n1842 );
buf ( n2343 , n771 );
and ( n2344 , n2343 , n1845 );
buf ( n2345 , n803 );
and ( n2346 , n2345 , n1848 );
or ( n2347 , n2340 , n2342 , n2344 , n2346 );
and ( n2348 , n2333 , n2347 );
not ( n2349 , n2347 );
and ( n2350 , n2325 , n2326 );
xor ( n2351 , n2349 , n2350 );
and ( n2352 , n2351 , n1859 );
or ( n2353 , n2348 , n2352 );
not ( n2354 , n2353 );
not ( n2355 , n2354 );
or ( n2356 , n2332 , n2355 );
not ( n2357 , n1859 );
buf ( n2358 , n743 );
not ( n2359 , n2358 );
not ( n2360 , n2359 );
buf ( n2361 , n2360 );
and ( n2362 , n2337 , n2338 );
xor ( n2363 , n2361 , n2362 );
and ( n2364 , n2363 , n1838 );
buf ( n2365 , n837 );
and ( n2366 , n2365 , n1842 );
buf ( n2367 , n772 );
and ( n2368 , n2367 , n1845 );
buf ( n2369 , n804 );
and ( n2370 , n2369 , n1848 );
or ( n2371 , n2364 , n2366 , n2368 , n2370 );
and ( n2372 , n2357 , n2371 );
not ( n2373 , n2371 );
and ( n2374 , n2349 , n2350 );
xor ( n2375 , n2373 , n2374 );
and ( n2376 , n2375 , n1859 );
or ( n2377 , n2372 , n2376 );
not ( n2378 , n2377 );
not ( n2379 , n2378 );
or ( n2380 , n2356 , n2379 );
not ( n2381 , n1859 );
buf ( n2382 , n744 );
not ( n2383 , n2382 );
not ( n2384 , n2383 );
buf ( n2385 , n2384 );
and ( n2386 , n2361 , n2362 );
xor ( n2387 , n2385 , n2386 );
and ( n2388 , n2387 , n1838 );
buf ( n2389 , n838 );
and ( n2390 , n2389 , n1842 );
buf ( n2391 , n773 );
and ( n2392 , n2391 , n1845 );
buf ( n2393 , n805 );
and ( n2394 , n2393 , n1848 );
or ( n2395 , n2388 , n2390 , n2392 , n2394 );
and ( n2396 , n2381 , n2395 );
not ( n2397 , n2395 );
and ( n2398 , n2373 , n2374 );
xor ( n2399 , n2397 , n2398 );
and ( n2400 , n2399 , n1859 );
or ( n2401 , n2396 , n2400 );
not ( n2402 , n2401 );
not ( n2403 , n2402 );
or ( n2404 , n2380 , n2403 );
not ( n2405 , n1859 );
buf ( n2406 , n745 );
not ( n2407 , n2406 );
not ( n2408 , n2407 );
buf ( n2409 , n2408 );
and ( n2410 , n2385 , n2386 );
xor ( n2411 , n2409 , n2410 );
and ( n2412 , n2411 , n1838 );
buf ( n2413 , n839 );
and ( n2414 , n2413 , n1842 );
buf ( n2415 , n774 );
and ( n2416 , n2415 , n1845 );
buf ( n2417 , n806 );
and ( n2418 , n2417 , n1848 );
or ( n2419 , n2412 , n2414 , n2416 , n2418 );
and ( n2420 , n2405 , n2419 );
not ( n2421 , n2419 );
and ( n2422 , n2397 , n2398 );
xor ( n2423 , n2421 , n2422 );
and ( n2424 , n2423 , n1859 );
or ( n2425 , n2420 , n2424 );
not ( n2426 , n2425 );
not ( n2427 , n2426 );
or ( n2428 , n2404 , n2427 );
not ( n2429 , n1859 );
buf ( n2430 , n746 );
not ( n2431 , n2430 );
not ( n2432 , n2431 );
buf ( n2433 , n2432 );
and ( n2434 , n2409 , n2410 );
xor ( n2435 , n2433 , n2434 );
and ( n2436 , n2435 , n1838 );
buf ( n2437 , n840 );
and ( n2438 , n2437 , n1842 );
buf ( n2439 , n775 );
and ( n2440 , n2439 , n1845 );
buf ( n2441 , n807 );
and ( n2442 , n2441 , n1848 );
or ( n2443 , n2436 , n2438 , n2440 , n2442 );
and ( n2444 , n2429 , n2443 );
not ( n2445 , n2443 );
and ( n2446 , n2421 , n2422 );
xor ( n2447 , n2445 , n2446 );
and ( n2448 , n2447 , n1859 );
or ( n2449 , n2444 , n2448 );
not ( n2450 , n2449 );
not ( n2451 , n2450 );
or ( n2452 , n2428 , n2451 );
not ( n2453 , n1859 );
buf ( n2454 , n747 );
not ( n2455 , n2454 );
not ( n2456 , n2455 );
buf ( n2457 , n2456 );
and ( n2458 , n2433 , n2434 );
xor ( n2459 , n2457 , n2458 );
and ( n2460 , n2459 , n1838 );
buf ( n2461 , n841 );
and ( n2462 , n2461 , n1842 );
buf ( n2463 , n776 );
and ( n2464 , n2463 , n1845 );
buf ( n2465 , n808 );
and ( n2466 , n2465 , n1848 );
or ( n2467 , n2460 , n2462 , n2464 , n2466 );
and ( n2468 , n2453 , n2467 );
not ( n2469 , n2467 );
and ( n2470 , n2445 , n2446 );
xor ( n2471 , n2469 , n2470 );
and ( n2472 , n2471 , n1859 );
or ( n2473 , n2468 , n2472 );
not ( n2474 , n2473 );
not ( n2475 , n2474 );
or ( n2476 , n2452 , n2475 );
not ( n2477 , n1859 );
buf ( n2478 , n748 );
not ( n2479 , n2478 );
not ( n2480 , n2479 );
buf ( n2481 , n2480 );
and ( n2482 , n2457 , n2458 );
xor ( n2483 , n2481 , n2482 );
and ( n2484 , n2483 , n1838 );
buf ( n2485 , n842 );
and ( n2486 , n2485 , n1842 );
buf ( n2487 , n777 );
and ( n2488 , n2487 , n1845 );
buf ( n2489 , n809 );
and ( n2490 , n2489 , n1848 );
or ( n2491 , n2484 , n2486 , n2488 , n2490 );
and ( n2492 , n2477 , n2491 );
not ( n2493 , n2491 );
and ( n2494 , n2469 , n2470 );
xor ( n2495 , n2493 , n2494 );
and ( n2496 , n2495 , n1859 );
or ( n2497 , n2492 , n2496 );
not ( n2498 , n2497 );
not ( n2499 , n2498 );
or ( n2500 , n2476 , n2499 );
not ( n2501 , n1859 );
buf ( n2502 , n749 );
not ( n2503 , n2502 );
not ( n2504 , n2503 );
buf ( n2505 , n2504 );
and ( n2506 , n2481 , n2482 );
xor ( n2507 , n2505 , n2506 );
and ( n2508 , n2507 , n1838 );
buf ( n2509 , n843 );
and ( n2510 , n2509 , n1842 );
buf ( n2511 , n778 );
and ( n2512 , n2511 , n1845 );
buf ( n2513 , n810 );
and ( n2514 , n2513 , n1848 );
or ( n2515 , n2508 , n2510 , n2512 , n2514 );
and ( n2516 , n2501 , n2515 );
not ( n2517 , n2515 );
and ( n2518 , n2493 , n2494 );
xor ( n2519 , n2517 , n2518 );
and ( n2520 , n2519 , n1859 );
or ( n2521 , n2516 , n2520 );
not ( n2522 , n2521 );
not ( n2523 , n2522 );
or ( n2524 , n2500 , n2523 );
and ( n2525 , n2524 , n1859 );
not ( n2526 , n2525 );
and ( n2527 , n2526 , n1852 );
xor ( n2528 , n1852 , n1859 );
xor ( n2529 , n2528 , n1859 );
and ( n2530 , n2529 , n2525 );
or ( n2531 , n2527 , n2530 );
not ( n2532 , n946 );
and ( n2533 , n2532 , n1142 );
not ( n2534 , n1142 );
not ( n2535 , n1148 );
not ( n2536 , n1154 );
not ( n2537 , n1160 );
not ( n2538 , n952 );
not ( n2539 , n959 );
not ( n2540 , n965 );
not ( n2541 , n971 );
not ( n2542 , n977 );
not ( n2543 , n983 );
not ( n2544 , n989 );
not ( n2545 , n995 );
not ( n2546 , n1001 );
not ( n2547 , n1007 );
not ( n2548 , n1013 );
not ( n2549 , n1019 );
not ( n2550 , n1025 );
not ( n2551 , n1031 );
not ( n2552 , n1037 );
not ( n2553 , n1043 );
not ( n2554 , n1049 );
not ( n2555 , n1055 );
not ( n2556 , n1061 );
not ( n2557 , n1067 );
not ( n2558 , n1073 );
not ( n2559 , n1079 );
not ( n2560 , n1085 );
not ( n2561 , n911 );
and ( n2562 , n2560 , n2561 );
and ( n2563 , n2559 , n2562 );
and ( n2564 , n2558 , n2563 );
and ( n2565 , n2557 , n2564 );
and ( n2566 , n2556 , n2565 );
and ( n2567 , n2555 , n2566 );
and ( n2568 , n2554 , n2567 );
and ( n2569 , n2553 , n2568 );
and ( n2570 , n2552 , n2569 );
and ( n2571 , n2551 , n2570 );
and ( n2572 , n2550 , n2571 );
and ( n2573 , n2549 , n2572 );
and ( n2574 , n2548 , n2573 );
and ( n2575 , n2547 , n2574 );
and ( n2576 , n2546 , n2575 );
and ( n2577 , n2545 , n2576 );
and ( n2578 , n2544 , n2577 );
and ( n2579 , n2543 , n2578 );
and ( n2580 , n2542 , n2579 );
and ( n2581 , n2541 , n2580 );
and ( n2582 , n2540 , n2581 );
and ( n2583 , n2539 , n2582 );
and ( n2584 , n2538 , n2583 );
and ( n2585 , n2537 , n2584 );
and ( n2586 , n2536 , n2585 );
and ( n2587 , n2535 , n2586 );
xor ( n2588 , n2534 , n2587 );
and ( n2589 , n2588 , n946 );
or ( n2590 , n2533 , n2589 );
not ( n2591 , n2590 );
not ( n2592 , n2591 );
not ( n2593 , n2592 );
not ( n2594 , n2593 );
not ( n2595 , n946 );
not ( n2596 , n1124 );
not ( n2597 , n1130 );
not ( n2598 , n1136 );
and ( n2599 , n2534 , n2587 );
and ( n2600 , n2598 , n2599 );
and ( n2601 , n2597 , n2600 );
and ( n2602 , n2596 , n2601 );
xor ( n2603 , n2595 , n2602 );
buf ( n2604 , n946 );
and ( n2605 , n2603 , n2604 );
buf ( n2606 , n2605 );
not ( n2607 , n2606 );
not ( n2608 , n2607 );
not ( n2609 , n2608 );
not ( n2610 , n946 );
and ( n2611 , n2610 , n1124 );
xor ( n2612 , n2596 , n2601 );
and ( n2613 , n2612 , n946 );
or ( n2614 , n2611 , n2613 );
not ( n2615 , n2614 );
not ( n2616 , n2615 );
not ( n2617 , n2616 );
not ( n2618 , n946 );
and ( n2619 , n2618 , n1130 );
xor ( n2620 , n2597 , n2600 );
and ( n2621 , n2620 , n946 );
or ( n2622 , n2619 , n2621 );
not ( n2623 , n2622 );
not ( n2624 , n2623 );
not ( n2625 , n2624 );
not ( n2626 , n946 );
and ( n2627 , n2626 , n1136 );
xor ( n2628 , n2598 , n2599 );
and ( n2629 , n2628 , n946 );
or ( n2630 , n2627 , n2629 );
not ( n2631 , n2630 );
not ( n2632 , n2631 );
not ( n2633 , n2632 );
not ( n2634 , n2592 );
and ( n2635 , n2633 , n2634 );
and ( n2636 , n2625 , n2635 );
and ( n2637 , n2617 , n2636 );
and ( n2638 , n2609 , n2637 );
not ( n2639 , n2638 );
and ( n2640 , n2639 , n946 );
buf ( n2641 , n2640 );
not ( n2642 , n2641 );
not ( n2643 , n946 );
and ( n2644 , n2643 , n2632 );
xor ( n2645 , n2633 , n2634 );
and ( n2646 , n2645 , n946 );
or ( n2647 , n2644 , n2646 );
and ( n2648 , n2642 , n2647 );
not ( n2649 , n2647 );
not ( n2650 , n2592 );
xor ( n2651 , n2649 , n2650 );
and ( n2652 , n2651 , n2641 );
or ( n2653 , n2648 , n2652 );
not ( n2654 , n2653 );
not ( n2655 , n2654 );
or ( n2656 , n2594 , n2655 );
and ( n2657 , n2656 , n2641 );
not ( n2658 , n2657 );
and ( n2659 , n2658 , n2594 );
xor ( n2660 , n2594 , n2641 );
xor ( n2661 , n2660 , n2641 );
and ( n2662 , n2661 , n2657 );
or ( n2663 , n2659 , n2662 );
not ( n2664 , n2657 );
and ( n2665 , n2664 , n2655 );
xor ( n2666 , n2655 , n2641 );
and ( n2667 , n2660 , n2641 );
xor ( n2668 , n2666 , n2667 );
and ( n2669 , n2668 , n2657 );
or ( n2670 , n2665 , n2669 );
and ( n2671 , n2663 , n2670 );
and ( n2672 , n2531 , n2671 );
not ( n2673 , n2663 );
and ( n2674 , n2673 , n2670 );
and ( n2675 , n2531 , n2674 );
buf ( n2676 , n814 );
not ( n2677 , n2676 );
not ( n2678 , n1859 );
not ( n2679 , n1859 );
and ( n2680 , n2679 , n1891 );
not ( n2681 , n1891 );
not ( n2682 , n1868 );
not ( n2683 , n1850 );
and ( n2684 , n2682 , n2683 );
xor ( n2685 , n2681 , n2684 );
and ( n2686 , n2685 , n1859 );
or ( n2687 , n2680 , n2686 );
not ( n2688 , n2687 );
buf ( n2689 , n2688 );
buf ( n2690 , n2689 );
not ( n2691 , n2690 );
and ( n2692 , n2678 , n2691 );
not ( n2693 , n2691 );
not ( n2694 , n1859 );
and ( n2695 , n2694 , n1868 );
xor ( n2696 , n2682 , n2683 );
and ( n2697 , n2696 , n1859 );
or ( n2698 , n2695 , n2697 );
not ( n2699 , n2698 );
buf ( n2700 , n2699 );
buf ( n2701 , n2700 );
not ( n2702 , n2701 );
not ( n2703 , n2702 );
xor ( n2704 , n2693 , n2703 );
and ( n2705 , n2704 , n1859 );
or ( n2706 , n2692 , n2705 );
and ( n2707 , n2677 , n2706 );
not ( n2708 , n2702 );
not ( n2709 , n2708 );
not ( n2710 , n1859 );
buf ( n2711 , n845 );
and ( n2712 , n2711 , n1842 );
buf ( n2713 , n780 );
and ( n2714 , n2713 , n1845 );
buf ( n2715 , n812 );
and ( n2716 , n2715 , n1848 );
or ( n2717 , 1'b0 , n2712 , n2714 , n2716 );
not ( n2718 , n2717 );
and ( n2719 , n2505 , n2506 );
buf ( n2720 , n2719 );
and ( n2721 , n2720 , n1838 );
buf ( n2722 , n844 );
and ( n2723 , n2722 , n1842 );
buf ( n2724 , n779 );
and ( n2725 , n2724 , n1845 );
buf ( n2726 , n811 );
and ( n2727 , n2726 , n1848 );
or ( n2728 , n2721 , n2723 , n2725 , n2727 );
not ( n2729 , n2728 );
not ( n2730 , n2515 );
not ( n2731 , n2491 );
not ( n2732 , n2467 );
not ( n2733 , n2443 );
not ( n2734 , n2419 );
not ( n2735 , n2395 );
not ( n2736 , n2371 );
not ( n2737 , n2347 );
not ( n2738 , n2323 );
not ( n2739 , n2299 );
not ( n2740 , n2275 );
not ( n2741 , n2251 );
not ( n2742 , n2227 );
not ( n2743 , n2203 );
not ( n2744 , n2179 );
not ( n2745 , n2155 );
not ( n2746 , n2131 );
not ( n2747 , n2107 );
not ( n2748 , n2083 );
not ( n2749 , n2059 );
not ( n2750 , n2035 );
not ( n2751 , n2011 );
not ( n2752 , n1987 );
not ( n2753 , n1963 );
not ( n2754 , n1939 );
not ( n2755 , n1915 );
and ( n2756 , n2681 , n2684 );
and ( n2757 , n2755 , n2756 );
and ( n2758 , n2754 , n2757 );
and ( n2759 , n2753 , n2758 );
and ( n2760 , n2752 , n2759 );
and ( n2761 , n2751 , n2760 );
and ( n2762 , n2750 , n2761 );
and ( n2763 , n2749 , n2762 );
and ( n2764 , n2748 , n2763 );
and ( n2765 , n2747 , n2764 );
and ( n2766 , n2746 , n2765 );
and ( n2767 , n2745 , n2766 );
and ( n2768 , n2744 , n2767 );
and ( n2769 , n2743 , n2768 );
and ( n2770 , n2742 , n2769 );
and ( n2771 , n2741 , n2770 );
and ( n2772 , n2740 , n2771 );
and ( n2773 , n2739 , n2772 );
and ( n2774 , n2738 , n2773 );
and ( n2775 , n2737 , n2774 );
and ( n2776 , n2736 , n2775 );
and ( n2777 , n2735 , n2776 );
and ( n2778 , n2734 , n2777 );
and ( n2779 , n2733 , n2778 );
and ( n2780 , n2732 , n2779 );
and ( n2781 , n2731 , n2780 );
and ( n2782 , n2730 , n2781 );
and ( n2783 , n2729 , n2782 );
and ( n2784 , n2718 , n2783 );
xor ( n2785 , n2710 , n2784 );
buf ( n2786 , n1859 );
and ( n2787 , n2785 , n2786 );
buf ( n2788 , n2787 );
not ( n2789 , n2788 );
not ( n2790 , n2789 );
not ( n2791 , n2790 );
not ( n2792 , n1859 );
and ( n2793 , n2792 , n2717 );
xor ( n2794 , n2718 , n2783 );
and ( n2795 , n2794 , n1859 );
or ( n2796 , n2793 , n2795 );
not ( n2797 , n2796 );
not ( n2798 , n2797 );
not ( n2799 , n2798 );
not ( n2800 , n1859 );
and ( n2801 , n2800 , n2728 );
xor ( n2802 , n2729 , n2782 );
and ( n2803 , n2802 , n1859 );
or ( n2804 , n2801 , n2803 );
not ( n2805 , n2804 );
not ( n2806 , n2805 );
not ( n2807 , n2806 );
not ( n2808 , n1859 );
and ( n2809 , n2808 , n2515 );
xor ( n2810 , n2730 , n2781 );
and ( n2811 , n2810 , n1859 );
or ( n2812 , n2809 , n2811 );
not ( n2813 , n2812 );
not ( n2814 , n2813 );
not ( n2815 , n2814 );
not ( n2816 , n1859 );
and ( n2817 , n2816 , n2491 );
xor ( n2818 , n2731 , n2780 );
and ( n2819 , n2818 , n1859 );
or ( n2820 , n2817 , n2819 );
not ( n2821 , n2820 );
not ( n2822 , n2821 );
not ( n2823 , n2822 );
not ( n2824 , n1859 );
and ( n2825 , n2824 , n2467 );
xor ( n2826 , n2732 , n2779 );
and ( n2827 , n2826 , n1859 );
or ( n2828 , n2825 , n2827 );
not ( n2829 , n2828 );
not ( n2830 , n2829 );
not ( n2831 , n2830 );
not ( n2832 , n1859 );
and ( n2833 , n2832 , n2443 );
xor ( n2834 , n2733 , n2778 );
and ( n2835 , n2834 , n1859 );
or ( n2836 , n2833 , n2835 );
not ( n2837 , n2836 );
not ( n2838 , n2837 );
not ( n2839 , n2838 );
not ( n2840 , n1859 );
and ( n2841 , n2840 , n2419 );
xor ( n2842 , n2734 , n2777 );
and ( n2843 , n2842 , n1859 );
or ( n2844 , n2841 , n2843 );
not ( n2845 , n2844 );
not ( n2846 , n2845 );
not ( n2847 , n2846 );
not ( n2848 , n1859 );
and ( n2849 , n2848 , n2395 );
xor ( n2850 , n2735 , n2776 );
and ( n2851 , n2850 , n1859 );
or ( n2852 , n2849 , n2851 );
not ( n2853 , n2852 );
not ( n2854 , n2853 );
not ( n2855 , n2854 );
not ( n2856 , n1859 );
and ( n2857 , n2856 , n2371 );
xor ( n2858 , n2736 , n2775 );
and ( n2859 , n2858 , n1859 );
or ( n2860 , n2857 , n2859 );
not ( n2861 , n2860 );
not ( n2862 , n2861 );
not ( n2863 , n2862 );
not ( n2864 , n1859 );
and ( n2865 , n2864 , n2347 );
xor ( n2866 , n2737 , n2774 );
and ( n2867 , n2866 , n1859 );
or ( n2868 , n2865 , n2867 );
not ( n2869 , n2868 );
not ( n2870 , n2869 );
not ( n2871 , n2870 );
not ( n2872 , n1859 );
and ( n2873 , n2872 , n2323 );
xor ( n2874 , n2738 , n2773 );
and ( n2875 , n2874 , n1859 );
or ( n2876 , n2873 , n2875 );
not ( n2877 , n2876 );
not ( n2878 , n2877 );
not ( n2879 , n2878 );
not ( n2880 , n1859 );
and ( n2881 , n2880 , n2299 );
xor ( n2882 , n2739 , n2772 );
and ( n2883 , n2882 , n1859 );
or ( n2884 , n2881 , n2883 );
not ( n2885 , n2884 );
not ( n2886 , n2885 );
not ( n2887 , n2886 );
not ( n2888 , n1859 );
and ( n2889 , n2888 , n2275 );
xor ( n2890 , n2740 , n2771 );
and ( n2891 , n2890 , n1859 );
or ( n2892 , n2889 , n2891 );
not ( n2893 , n2892 );
not ( n2894 , n2893 );
not ( n2895 , n2894 );
not ( n2896 , n1859 );
and ( n2897 , n2896 , n2251 );
xor ( n2898 , n2741 , n2770 );
and ( n2899 , n2898 , n1859 );
or ( n2900 , n2897 , n2899 );
not ( n2901 , n2900 );
not ( n2902 , n2901 );
not ( n2903 , n2902 );
not ( n2904 , n1859 );
and ( n2905 , n2904 , n2227 );
xor ( n2906 , n2742 , n2769 );
and ( n2907 , n2906 , n1859 );
or ( n2908 , n2905 , n2907 );
not ( n2909 , n2908 );
not ( n2910 , n2909 );
not ( n2911 , n2910 );
not ( n2912 , n1859 );
and ( n2913 , n2912 , n2203 );
xor ( n2914 , n2743 , n2768 );
and ( n2915 , n2914 , n1859 );
or ( n2916 , n2913 , n2915 );
not ( n2917 , n2916 );
not ( n2918 , n2917 );
not ( n2919 , n2918 );
not ( n2920 , n1859 );
and ( n2921 , n2920 , n2179 );
xor ( n2922 , n2744 , n2767 );
and ( n2923 , n2922 , n1859 );
or ( n2924 , n2921 , n2923 );
not ( n2925 , n2924 );
not ( n2926 , n2925 );
not ( n2927 , n2926 );
not ( n2928 , n1859 );
and ( n2929 , n2928 , n2155 );
xor ( n2930 , n2745 , n2766 );
and ( n2931 , n2930 , n1859 );
or ( n2932 , n2929 , n2931 );
not ( n2933 , n2932 );
not ( n2934 , n2933 );
not ( n2935 , n2934 );
not ( n2936 , n1859 );
and ( n2937 , n2936 , n2131 );
xor ( n2938 , n2746 , n2765 );
and ( n2939 , n2938 , n1859 );
or ( n2940 , n2937 , n2939 );
not ( n2941 , n2940 );
not ( n2942 , n2941 );
not ( n2943 , n2942 );
not ( n2944 , n1859 );
and ( n2945 , n2944 , n2107 );
xor ( n2946 , n2747 , n2764 );
and ( n2947 , n2946 , n1859 );
or ( n2948 , n2945 , n2947 );
not ( n2949 , n2948 );
not ( n2950 , n2949 );
not ( n2951 , n2950 );
not ( n2952 , n1859 );
and ( n2953 , n2952 , n2083 );
xor ( n2954 , n2748 , n2763 );
and ( n2955 , n2954 , n1859 );
or ( n2956 , n2953 , n2955 );
not ( n2957 , n2956 );
buf ( n2958 , n2957 );
buf ( n2959 , n2958 );
not ( n2960 , n2959 );
not ( n2961 , n2960 );
not ( n2962 , n1859 );
and ( n2963 , n2962 , n2059 );
xor ( n2964 , n2749 , n2762 );
and ( n2965 , n2964 , n1859 );
or ( n2966 , n2963 , n2965 );
not ( n2967 , n2966 );
buf ( n2968 , n2967 );
buf ( n2969 , n2968 );
not ( n2970 , n2969 );
not ( n2971 , n2970 );
not ( n2972 , n1859 );
and ( n2973 , n2972 , n2035 );
xor ( n2974 , n2750 , n2761 );
and ( n2975 , n2974 , n1859 );
or ( n2976 , n2973 , n2975 );
not ( n2977 , n2976 );
buf ( n2978 , n2977 );
buf ( n2979 , n2978 );
not ( n2980 , n2979 );
not ( n2981 , n2980 );
not ( n2982 , n1859 );
and ( n2983 , n2982 , n2011 );
xor ( n2984 , n2751 , n2760 );
and ( n2985 , n2984 , n1859 );
or ( n2986 , n2983 , n2985 );
not ( n2987 , n2986 );
buf ( n2988 , n2987 );
buf ( n2989 , n2988 );
not ( n2990 , n2989 );
not ( n2991 , n2990 );
not ( n2992 , n1859 );
and ( n2993 , n2992 , n1987 );
xor ( n2994 , n2752 , n2759 );
and ( n2995 , n2994 , n1859 );
or ( n2996 , n2993 , n2995 );
not ( n2997 , n2996 );
buf ( n2998 , n2997 );
buf ( n2999 , n2998 );
not ( n3000 , n2999 );
not ( n3001 , n3000 );
not ( n3002 , n1859 );
and ( n3003 , n3002 , n1963 );
xor ( n3004 , n2753 , n2758 );
and ( n3005 , n3004 , n1859 );
or ( n3006 , n3003 , n3005 );
not ( n3007 , n3006 );
buf ( n3008 , n3007 );
buf ( n3009 , n3008 );
not ( n3010 , n3009 );
not ( n3011 , n3010 );
not ( n3012 , n1859 );
and ( n3013 , n3012 , n1939 );
xor ( n3014 , n2754 , n2757 );
and ( n3015 , n3014 , n1859 );
or ( n3016 , n3013 , n3015 );
not ( n3017 , n3016 );
buf ( n3018 , n3017 );
buf ( n3019 , n3018 );
not ( n3020 , n3019 );
not ( n3021 , n3020 );
not ( n3022 , n1859 );
and ( n3023 , n3022 , n1915 );
xor ( n3024 , n2755 , n2756 );
and ( n3025 , n3024 , n1859 );
or ( n3026 , n3023 , n3025 );
not ( n3027 , n3026 );
buf ( n3028 , n3027 );
buf ( n3029 , n3028 );
not ( n3030 , n3029 );
not ( n3031 , n3030 );
and ( n3032 , n2693 , n2703 );
and ( n3033 , n3031 , n3032 );
and ( n3034 , n3021 , n3033 );
and ( n3035 , n3011 , n3034 );
and ( n3036 , n3001 , n3035 );
and ( n3037 , n2991 , n3036 );
and ( n3038 , n2981 , n3037 );
and ( n3039 , n2971 , n3038 );
and ( n3040 , n2961 , n3039 );
and ( n3041 , n2951 , n3040 );
and ( n3042 , n2943 , n3041 );
and ( n3043 , n2935 , n3042 );
and ( n3044 , n2927 , n3043 );
and ( n3045 , n2919 , n3044 );
and ( n3046 , n2911 , n3045 );
and ( n3047 , n2903 , n3046 );
and ( n3048 , n2895 , n3047 );
and ( n3049 , n2887 , n3048 );
and ( n3050 , n2879 , n3049 );
and ( n3051 , n2871 , n3050 );
and ( n3052 , n2863 , n3051 );
and ( n3053 , n2855 , n3052 );
and ( n3054 , n2847 , n3053 );
and ( n3055 , n2839 , n3054 );
and ( n3056 , n2831 , n3055 );
and ( n3057 , n2823 , n3056 );
and ( n3058 , n2815 , n3057 );
and ( n3059 , n2807 , n3058 );
and ( n3060 , n2799 , n3059 );
and ( n3061 , n2791 , n3060 );
not ( n3062 , n3061 );
and ( n3063 , n3062 , n1859 );
buf ( n3064 , n3063 );
not ( n3065 , n3064 );
and ( n3066 , n3065 , n2706 );
not ( n3067 , n2706 );
not ( n3068 , n2702 );
xor ( n3069 , n3067 , n3068 );
and ( n3070 , n3069 , n3064 );
or ( n3071 , n3066 , n3070 );
not ( n3072 , n3071 );
not ( n3073 , n3072 );
or ( n3074 , n2709 , n3073 );
not ( n3075 , n3064 );
not ( n3076 , n1859 );
and ( n3077 , n3076 , n3030 );
xor ( n3078 , n3031 , n3032 );
and ( n3079 , n3078 , n1859 );
or ( n3080 , n3077 , n3079 );
and ( n3081 , n3075 , n3080 );
not ( n3082 , n3080 );
and ( n3083 , n3067 , n3068 );
xor ( n3084 , n3082 , n3083 );
and ( n3085 , n3084 , n3064 );
or ( n3086 , n3081 , n3085 );
not ( n3087 , n3086 );
not ( n3088 , n3087 );
or ( n3089 , n3074 , n3088 );
not ( n3090 , n3064 );
not ( n3091 , n1859 );
and ( n3092 , n3091 , n3020 );
xor ( n3093 , n3021 , n3033 );
and ( n3094 , n3093 , n1859 );
or ( n3095 , n3092 , n3094 );
and ( n3096 , n3090 , n3095 );
not ( n3097 , n3095 );
and ( n3098 , n3082 , n3083 );
xor ( n3099 , n3097 , n3098 );
and ( n3100 , n3099 , n3064 );
or ( n3101 , n3096 , n3100 );
not ( n3102 , n3101 );
not ( n3103 , n3102 );
or ( n3104 , n3089 , n3103 );
not ( n3105 , n3064 );
not ( n3106 , n1859 );
and ( n3107 , n3106 , n3010 );
xor ( n3108 , n3011 , n3034 );
and ( n3109 , n3108 , n1859 );
or ( n3110 , n3107 , n3109 );
and ( n3111 , n3105 , n3110 );
not ( n3112 , n3110 );
and ( n3113 , n3097 , n3098 );
xor ( n3114 , n3112 , n3113 );
and ( n3115 , n3114 , n3064 );
or ( n3116 , n3111 , n3115 );
not ( n3117 , n3116 );
not ( n3118 , n3117 );
or ( n3119 , n3104 , n3118 );
not ( n3120 , n3064 );
not ( n3121 , n1859 );
and ( n3122 , n3121 , n3000 );
xor ( n3123 , n3001 , n3035 );
and ( n3124 , n3123 , n1859 );
or ( n3125 , n3122 , n3124 );
and ( n3126 , n3120 , n3125 );
not ( n3127 , n3125 );
and ( n3128 , n3112 , n3113 );
xor ( n3129 , n3127 , n3128 );
and ( n3130 , n3129 , n3064 );
or ( n3131 , n3126 , n3130 );
not ( n3132 , n3131 );
not ( n3133 , n3132 );
or ( n3134 , n3119 , n3133 );
not ( n3135 , n3064 );
not ( n3136 , n1859 );
and ( n3137 , n3136 , n2990 );
xor ( n3138 , n2991 , n3036 );
and ( n3139 , n3138 , n1859 );
or ( n3140 , n3137 , n3139 );
and ( n3141 , n3135 , n3140 );
not ( n3142 , n3140 );
and ( n3143 , n3127 , n3128 );
xor ( n3144 , n3142 , n3143 );
and ( n3145 , n3144 , n3064 );
or ( n3146 , n3141 , n3145 );
not ( n3147 , n3146 );
not ( n3148 , n3147 );
or ( n3149 , n3134 , n3148 );
not ( n3150 , n3064 );
not ( n3151 , n1859 );
and ( n3152 , n3151 , n2980 );
xor ( n3153 , n2981 , n3037 );
and ( n3154 , n3153 , n1859 );
or ( n3155 , n3152 , n3154 );
and ( n3156 , n3150 , n3155 );
not ( n3157 , n3155 );
and ( n3158 , n3142 , n3143 );
xor ( n3159 , n3157 , n3158 );
and ( n3160 , n3159 , n3064 );
or ( n3161 , n3156 , n3160 );
not ( n3162 , n3161 );
not ( n3163 , n3162 );
or ( n3164 , n3149 , n3163 );
not ( n3165 , n3064 );
not ( n3166 , n1859 );
and ( n3167 , n3166 , n2970 );
xor ( n3168 , n2971 , n3038 );
and ( n3169 , n3168 , n1859 );
or ( n3170 , n3167 , n3169 );
and ( n3171 , n3165 , n3170 );
not ( n3172 , n3170 );
and ( n3173 , n3157 , n3158 );
xor ( n3174 , n3172 , n3173 );
and ( n3175 , n3174 , n3064 );
or ( n3176 , n3171 , n3175 );
not ( n3177 , n3176 );
not ( n3178 , n3177 );
or ( n3179 , n3164 , n3178 );
not ( n3180 , n3064 );
not ( n3181 , n1859 );
and ( n3182 , n3181 , n2960 );
xor ( n3183 , n2961 , n3039 );
and ( n3184 , n3183 , n1859 );
or ( n3185 , n3182 , n3184 );
and ( n3186 , n3180 , n3185 );
not ( n3187 , n3185 );
and ( n3188 , n3172 , n3173 );
xor ( n3189 , n3187 , n3188 );
and ( n3190 , n3189 , n3064 );
or ( n3191 , n3186 , n3190 );
not ( n3192 , n3191 );
not ( n3193 , n3192 );
or ( n3194 , n3179 , n3193 );
not ( n3195 , n3064 );
not ( n3196 , n1859 );
and ( n3197 , n3196 , n2950 );
xor ( n3198 , n2951 , n3040 );
and ( n3199 , n3198 , n1859 );
or ( n3200 , n3197 , n3199 );
and ( n3201 , n3195 , n3200 );
not ( n3202 , n3200 );
and ( n3203 , n3187 , n3188 );
xor ( n3204 , n3202 , n3203 );
and ( n3205 , n3204 , n3064 );
or ( n3206 , n3201 , n3205 );
not ( n3207 , n3206 );
not ( n3208 , n3207 );
or ( n3209 , n3194 , n3208 );
not ( n3210 , n3064 );
not ( n3211 , n1859 );
and ( n3212 , n3211 , n2942 );
xor ( n3213 , n2943 , n3041 );
and ( n3214 , n3213 , n1859 );
or ( n3215 , n3212 , n3214 );
and ( n3216 , n3210 , n3215 );
not ( n3217 , n3215 );
and ( n3218 , n3202 , n3203 );
xor ( n3219 , n3217 , n3218 );
and ( n3220 , n3219 , n3064 );
or ( n3221 , n3216 , n3220 );
not ( n3222 , n3221 );
not ( n3223 , n3222 );
or ( n3224 , n3209 , n3223 );
not ( n3225 , n3064 );
not ( n3226 , n1859 );
and ( n3227 , n3226 , n2934 );
xor ( n3228 , n2935 , n3042 );
and ( n3229 , n3228 , n1859 );
or ( n3230 , n3227 , n3229 );
and ( n3231 , n3225 , n3230 );
not ( n3232 , n3230 );
and ( n3233 , n3217 , n3218 );
xor ( n3234 , n3232 , n3233 );
and ( n3235 , n3234 , n3064 );
or ( n3236 , n3231 , n3235 );
not ( n3237 , n3236 );
not ( n3238 , n3237 );
or ( n3239 , n3224 , n3238 );
not ( n3240 , n3064 );
not ( n3241 , n1859 );
and ( n3242 , n3241 , n2926 );
xor ( n3243 , n2927 , n3043 );
and ( n3244 , n3243 , n1859 );
or ( n3245 , n3242 , n3244 );
and ( n3246 , n3240 , n3245 );
not ( n3247 , n3245 );
and ( n3248 , n3232 , n3233 );
xor ( n3249 , n3247 , n3248 );
and ( n3250 , n3249 , n3064 );
or ( n3251 , n3246 , n3250 );
not ( n3252 , n3251 );
not ( n3253 , n3252 );
or ( n3254 , n3239 , n3253 );
not ( n3255 , n3064 );
not ( n3256 , n1859 );
and ( n3257 , n3256 , n2918 );
xor ( n3258 , n2919 , n3044 );
and ( n3259 , n3258 , n1859 );
or ( n3260 , n3257 , n3259 );
and ( n3261 , n3255 , n3260 );
not ( n3262 , n3260 );
and ( n3263 , n3247 , n3248 );
xor ( n3264 , n3262 , n3263 );
and ( n3265 , n3264 , n3064 );
or ( n3266 , n3261 , n3265 );
not ( n3267 , n3266 );
not ( n3268 , n3267 );
or ( n3269 , n3254 , n3268 );
not ( n3270 , n3064 );
not ( n3271 , n1859 );
and ( n3272 , n3271 , n2910 );
xor ( n3273 , n2911 , n3045 );
and ( n3274 , n3273 , n1859 );
or ( n3275 , n3272 , n3274 );
and ( n3276 , n3270 , n3275 );
not ( n3277 , n3275 );
and ( n3278 , n3262 , n3263 );
xor ( n3279 , n3277 , n3278 );
and ( n3280 , n3279 , n3064 );
or ( n3281 , n3276 , n3280 );
not ( n3282 , n3281 );
not ( n3283 , n3282 );
or ( n3284 , n3269 , n3283 );
not ( n3285 , n3064 );
not ( n3286 , n1859 );
and ( n3287 , n3286 , n2902 );
xor ( n3288 , n2903 , n3046 );
and ( n3289 , n3288 , n1859 );
or ( n3290 , n3287 , n3289 );
and ( n3291 , n3285 , n3290 );
not ( n3292 , n3290 );
and ( n3293 , n3277 , n3278 );
xor ( n3294 , n3292 , n3293 );
and ( n3295 , n3294 , n3064 );
or ( n3296 , n3291 , n3295 );
not ( n3297 , n3296 );
not ( n3298 , n3297 );
or ( n3299 , n3284 , n3298 );
not ( n3300 , n3064 );
not ( n3301 , n1859 );
and ( n3302 , n3301 , n2894 );
xor ( n3303 , n2895 , n3047 );
and ( n3304 , n3303 , n1859 );
or ( n3305 , n3302 , n3304 );
and ( n3306 , n3300 , n3305 );
not ( n3307 , n3305 );
and ( n3308 , n3292 , n3293 );
xor ( n3309 , n3307 , n3308 );
and ( n3310 , n3309 , n3064 );
or ( n3311 , n3306 , n3310 );
not ( n3312 , n3311 );
not ( n3313 , n3312 );
or ( n3314 , n3299 , n3313 );
not ( n3315 , n3064 );
not ( n3316 , n1859 );
and ( n3317 , n3316 , n2886 );
xor ( n3318 , n2887 , n3048 );
and ( n3319 , n3318 , n1859 );
or ( n3320 , n3317 , n3319 );
and ( n3321 , n3315 , n3320 );
not ( n3322 , n3320 );
and ( n3323 , n3307 , n3308 );
xor ( n3324 , n3322 , n3323 );
and ( n3325 , n3324 , n3064 );
or ( n3326 , n3321 , n3325 );
not ( n3327 , n3326 );
not ( n3328 , n3327 );
or ( n3329 , n3314 , n3328 );
not ( n3330 , n3064 );
not ( n3331 , n1859 );
and ( n3332 , n3331 , n2878 );
xor ( n3333 , n2879 , n3049 );
and ( n3334 , n3333 , n1859 );
or ( n3335 , n3332 , n3334 );
and ( n3336 , n3330 , n3335 );
not ( n3337 , n3335 );
and ( n3338 , n3322 , n3323 );
xor ( n3339 , n3337 , n3338 );
and ( n3340 , n3339 , n3064 );
or ( n3341 , n3336 , n3340 );
not ( n3342 , n3341 );
not ( n3343 , n3342 );
or ( n3344 , n3329 , n3343 );
not ( n3345 , n3064 );
not ( n3346 , n1859 );
and ( n3347 , n3346 , n2870 );
xor ( n3348 , n2871 , n3050 );
and ( n3349 , n3348 , n1859 );
or ( n3350 , n3347 , n3349 );
and ( n3351 , n3345 , n3350 );
not ( n3352 , n3350 );
and ( n3353 , n3337 , n3338 );
xor ( n3354 , n3352 , n3353 );
and ( n3355 , n3354 , n3064 );
or ( n3356 , n3351 , n3355 );
not ( n3357 , n3356 );
not ( n3358 , n3357 );
or ( n3359 , n3344 , n3358 );
not ( n3360 , n3064 );
not ( n3361 , n1859 );
and ( n3362 , n3361 , n2862 );
xor ( n3363 , n2863 , n3051 );
and ( n3364 , n3363 , n1859 );
or ( n3365 , n3362 , n3364 );
and ( n3366 , n3360 , n3365 );
not ( n3367 , n3365 );
and ( n3368 , n3352 , n3353 );
xor ( n3369 , n3367 , n3368 );
and ( n3370 , n3369 , n3064 );
or ( n3371 , n3366 , n3370 );
not ( n3372 , n3371 );
not ( n3373 , n3372 );
or ( n3374 , n3359 , n3373 );
not ( n3375 , n3064 );
not ( n3376 , n1859 );
and ( n3377 , n3376 , n2854 );
xor ( n3378 , n2855 , n3052 );
and ( n3379 , n3378 , n1859 );
or ( n3380 , n3377 , n3379 );
and ( n3381 , n3375 , n3380 );
not ( n3382 , n3380 );
and ( n3383 , n3367 , n3368 );
xor ( n3384 , n3382 , n3383 );
and ( n3385 , n3384 , n3064 );
or ( n3386 , n3381 , n3385 );
not ( n3387 , n3386 );
not ( n3388 , n3387 );
or ( n3389 , n3374 , n3388 );
not ( n3390 , n3064 );
not ( n3391 , n1859 );
and ( n3392 , n3391 , n2846 );
xor ( n3393 , n2847 , n3053 );
and ( n3394 , n3393 , n1859 );
or ( n3395 , n3392 , n3394 );
and ( n3396 , n3390 , n3395 );
not ( n3397 , n3395 );
and ( n3398 , n3382 , n3383 );
xor ( n3399 , n3397 , n3398 );
and ( n3400 , n3399 , n3064 );
or ( n3401 , n3396 , n3400 );
not ( n3402 , n3401 );
not ( n3403 , n3402 );
or ( n3404 , n3389 , n3403 );
not ( n3405 , n3064 );
not ( n3406 , n1859 );
and ( n3407 , n3406 , n2838 );
xor ( n3408 , n2839 , n3054 );
and ( n3409 , n3408 , n1859 );
or ( n3410 , n3407 , n3409 );
and ( n3411 , n3405 , n3410 );
not ( n3412 , n3410 );
and ( n3413 , n3397 , n3398 );
xor ( n3414 , n3412 , n3413 );
and ( n3415 , n3414 , n3064 );
or ( n3416 , n3411 , n3415 );
not ( n3417 , n3416 );
not ( n3418 , n3417 );
or ( n3419 , n3404 , n3418 );
not ( n3420 , n3064 );
not ( n3421 , n1859 );
and ( n3422 , n3421 , n2830 );
xor ( n3423 , n2831 , n3055 );
and ( n3424 , n3423 , n1859 );
or ( n3425 , n3422 , n3424 );
and ( n3426 , n3420 , n3425 );
not ( n3427 , n3425 );
and ( n3428 , n3412 , n3413 );
xor ( n3429 , n3427 , n3428 );
and ( n3430 , n3429 , n3064 );
or ( n3431 , n3426 , n3430 );
not ( n3432 , n3431 );
not ( n3433 , n3432 );
or ( n3434 , n3419 , n3433 );
not ( n3435 , n3064 );
not ( n3436 , n1859 );
and ( n3437 , n3436 , n2822 );
xor ( n3438 , n2823 , n3056 );
and ( n3439 , n3438 , n1859 );
or ( n3440 , n3437 , n3439 );
and ( n3441 , n3435 , n3440 );
not ( n3442 , n3440 );
and ( n3443 , n3427 , n3428 );
xor ( n3444 , n3442 , n3443 );
and ( n3445 , n3444 , n3064 );
or ( n3446 , n3441 , n3445 );
not ( n3447 , n3446 );
not ( n3448 , n3447 );
or ( n3449 , n3434 , n3448 );
not ( n3450 , n3064 );
not ( n3451 , n1859 );
and ( n3452 , n3451 , n2814 );
xor ( n3453 , n2815 , n3057 );
and ( n3454 , n3453 , n1859 );
or ( n3455 , n3452 , n3454 );
and ( n3456 , n3450 , n3455 );
not ( n3457 , n3455 );
and ( n3458 , n3442 , n3443 );
xor ( n3459 , n3457 , n3458 );
and ( n3460 , n3459 , n3064 );
or ( n3461 , n3456 , n3460 );
not ( n3462 , n3461 );
not ( n3463 , n3462 );
or ( n3464 , n3449 , n3463 );
not ( n3465 , n3064 );
not ( n3466 , n1859 );
and ( n3467 , n3466 , n2806 );
xor ( n3468 , n2807 , n3058 );
and ( n3469 , n3468 , n1859 );
or ( n3470 , n3467 , n3469 );
and ( n3471 , n3465 , n3470 );
not ( n3472 , n3470 );
and ( n3473 , n3457 , n3458 );
xor ( n3474 , n3472 , n3473 );
and ( n3475 , n3474 , n3064 );
or ( n3476 , n3471 , n3475 );
not ( n3477 , n3476 );
not ( n3478 , n3477 );
or ( n3479 , n3464 , n3478 );
and ( n3480 , n3479 , n3064 );
not ( n3481 , n3480 );
and ( n3482 , n3481 , n3073 );
xor ( n3483 , n3073 , n3064 );
xor ( n3484 , n2709 , n3064 );
and ( n3485 , n3484 , n3064 );
xor ( n3486 , n3483 , n3485 );
and ( n3487 , n3486 , n3480 );
or ( n3488 , n3482 , n3487 );
and ( n3489 , n3488 , n2676 );
or ( n3490 , n2707 , n3489 );
nor ( n3491 , n2673 , n2670 );
and ( n3492 , n3490 , n3491 );
nor ( n3493 , n2663 , n2670 );
and ( n3494 , n2706 , n3493 );
or ( n3495 , n2672 , n2675 , n3492 , n3494 );
not ( n3496 , n1425 );
not ( n3497 , n1439 );
nor ( n3498 , n3496 , n1432 , n3497 );
not ( n3499 , n3498 );
nor ( n3500 , n1425 , n1432 , n3497 );
not ( n3501 , n3500 );
and ( n3502 , n1425 , n1432 , n3497 );
not ( n3503 , n3502 );
and ( n3504 , n3496 , n1432 , n3497 );
not ( n3505 , n3504 );
nor ( n3506 , n3496 , n1432 , n1439 );
not ( n3507 , n3506 );
nor ( n3508 , n1425 , n1432 , n1439 );
not ( n3509 , n3508 );
buf ( n3510 , n719 );
and ( n3511 , n3509 , n3510 );
buf ( n3512 , n3511 );
and ( n3513 , n3507 , n3512 );
buf ( n3514 , n3506 );
or ( n3515 , n3513 , n3514 );
and ( n3516 , n3505 , n3515 );
buf ( n3517 , n3516 );
and ( n3518 , n3503 , n3517 );
buf ( n3519 , n3502 );
or ( n3520 , n3518 , n3519 );
and ( n3521 , n3501 , n3520 );
not ( n3522 , n2676 );
and ( n3523 , n3522 , n3510 );
buf ( n3524 , n2676 );
or ( n3525 , n3523 , n3524 );
and ( n3526 , n3525 , n3500 );
or ( n3527 , n3521 , n3526 );
and ( n3528 , n3499 , n3527 );
not ( n3529 , n2676 );
not ( n3530 , n3529 );
and ( n3531 , n3530 , n3510 );
buf ( n3532 , n3529 );
or ( n3533 , n3531 , n3532 );
and ( n3534 , n3533 , n3498 );
or ( n3535 , n3528 , n3534 );
not ( n3536 , n3535 );
not ( n3537 , n3498 );
not ( n3538 , n3500 );
not ( n3539 , n3502 );
not ( n3540 , n3504 );
not ( n3541 , n3506 );
not ( n3542 , n3508 );
buf ( n3543 , n720 );
and ( n3544 , n3542 , n3543 );
buf ( n3545 , n3544 );
and ( n3546 , n3541 , n3545 );
buf ( n3547 , n3546 );
and ( n3548 , n3540 , n3547 );
buf ( n3549 , n3504 );
or ( n3550 , n3548 , n3549 );
and ( n3551 , n3539 , n3550 );
buf ( n3552 , n3502 );
or ( n3553 , n3551 , n3552 );
and ( n3554 , n3538 , n3553 );
not ( n3555 , n2676 );
and ( n3556 , n3555 , n3543 );
buf ( n3557 , n2676 );
or ( n3558 , n3556 , n3557 );
and ( n3559 , n3558 , n3500 );
or ( n3560 , n3554 , n3559 );
and ( n3561 , n3537 , n3560 );
not ( n3562 , n3529 );
and ( n3563 , n3562 , n3543 );
buf ( n3564 , n3529 );
or ( n3565 , n3563 , n3564 );
and ( n3566 , n3565 , n3498 );
or ( n3567 , n3561 , n3566 );
not ( n3568 , n3567 );
nor ( n3569 , n3536 , n3568 );
and ( n3570 , n3495 , n3569 );
nor ( n3571 , n3536 , n3567 );
nor ( n3572 , n3535 , n3567 );
or ( n3573 , n3571 , n3572 );
nor ( n3574 , n3535 , n3568 );
or ( n3575 , n3573 , n3574 );
buf ( n3576 , n3575 );
and ( n3577 , n1447 , n3576 );
or ( n3578 , n3570 , n3577 );
and ( n3579 , n1707 , n1691 , n1698 , n1705 );
and ( n3580 , n3578 , n3579 );
buf ( n3581 , n685 );
or ( n3582 , n3491 , n2674 );
or ( n3583 , n3582 , n2671 );
and ( n3584 , n3581 , n3583 );
not ( n3585 , n911 );
not ( n3586 , n3585 );
not ( n3587 , n946 );
and ( n3588 , n3587 , n1085 );
not ( n3589 , n1085 );
not ( n3590 , n911 );
xor ( n3591 , n3589 , n3590 );
and ( n3592 , n3591 , n946 );
or ( n3593 , n3588 , n3592 );
not ( n3594 , n3593 );
not ( n3595 , n3594 );
or ( n3596 , n3586 , n3595 );
not ( n3597 , n946 );
and ( n3598 , n3597 , n1079 );
not ( n3599 , n1079 );
and ( n3600 , n3589 , n3590 );
xor ( n3601 , n3599 , n3600 );
and ( n3602 , n3601 , n946 );
or ( n3603 , n3598 , n3602 );
not ( n3604 , n3603 );
not ( n3605 , n3604 );
or ( n3606 , n3596 , n3605 );
not ( n3607 , n946 );
and ( n3608 , n3607 , n1073 );
not ( n3609 , n1073 );
and ( n3610 , n3599 , n3600 );
xor ( n3611 , n3609 , n3610 );
and ( n3612 , n3611 , n946 );
or ( n3613 , n3608 , n3612 );
not ( n3614 , n3613 );
not ( n3615 , n3614 );
or ( n3616 , n3606 , n3615 );
not ( n3617 , n946 );
and ( n3618 , n3617 , n1067 );
not ( n3619 , n1067 );
and ( n3620 , n3609 , n3610 );
xor ( n3621 , n3619 , n3620 );
and ( n3622 , n3621 , n946 );
or ( n3623 , n3618 , n3622 );
not ( n3624 , n3623 );
not ( n3625 , n3624 );
or ( n3626 , n3616 , n3625 );
not ( n3627 , n946 );
and ( n3628 , n3627 , n1061 );
not ( n3629 , n1061 );
and ( n3630 , n3619 , n3620 );
xor ( n3631 , n3629 , n3630 );
and ( n3632 , n3631 , n946 );
or ( n3633 , n3628 , n3632 );
not ( n3634 , n3633 );
not ( n3635 , n3634 );
or ( n3636 , n3626 , n3635 );
not ( n3637 , n946 );
and ( n3638 , n3637 , n1055 );
not ( n3639 , n1055 );
and ( n3640 , n3629 , n3630 );
xor ( n3641 , n3639 , n3640 );
and ( n3642 , n3641 , n946 );
or ( n3643 , n3638 , n3642 );
not ( n3644 , n3643 );
not ( n3645 , n3644 );
or ( n3646 , n3636 , n3645 );
not ( n3647 , n946 );
and ( n3648 , n3647 , n1049 );
not ( n3649 , n1049 );
and ( n3650 , n3639 , n3640 );
xor ( n3651 , n3649 , n3650 );
and ( n3652 , n3651 , n946 );
or ( n3653 , n3648 , n3652 );
not ( n3654 , n3653 );
not ( n3655 , n3654 );
or ( n3656 , n3646 , n3655 );
not ( n3657 , n946 );
and ( n3658 , n3657 , n1043 );
not ( n3659 , n1043 );
and ( n3660 , n3649 , n3650 );
xor ( n3661 , n3659 , n3660 );
and ( n3662 , n3661 , n946 );
or ( n3663 , n3658 , n3662 );
not ( n3664 , n3663 );
not ( n3665 , n3664 );
or ( n3666 , n3656 , n3665 );
not ( n3667 , n946 );
and ( n3668 , n3667 , n1037 );
not ( n3669 , n1037 );
and ( n3670 , n3659 , n3660 );
xor ( n3671 , n3669 , n3670 );
and ( n3672 , n3671 , n946 );
or ( n3673 , n3668 , n3672 );
not ( n3674 , n3673 );
not ( n3675 , n3674 );
or ( n3676 , n3666 , n3675 );
not ( n3677 , n946 );
and ( n3678 , n3677 , n1031 );
not ( n3679 , n1031 );
and ( n3680 , n3669 , n3670 );
xor ( n3681 , n3679 , n3680 );
and ( n3682 , n3681 , n946 );
or ( n3683 , n3678 , n3682 );
not ( n3684 , n3683 );
not ( n3685 , n3684 );
or ( n3686 , n3676 , n3685 );
not ( n3687 , n946 );
and ( n3688 , n3687 , n1025 );
not ( n3689 , n1025 );
and ( n3690 , n3679 , n3680 );
xor ( n3691 , n3689 , n3690 );
and ( n3692 , n3691 , n946 );
or ( n3693 , n3688 , n3692 );
not ( n3694 , n3693 );
not ( n3695 , n3694 );
or ( n3696 , n3686 , n3695 );
not ( n3697 , n946 );
and ( n3698 , n3697 , n1019 );
not ( n3699 , n1019 );
and ( n3700 , n3689 , n3690 );
xor ( n3701 , n3699 , n3700 );
and ( n3702 , n3701 , n946 );
or ( n3703 , n3698 , n3702 );
not ( n3704 , n3703 );
not ( n3705 , n3704 );
or ( n3706 , n3696 , n3705 );
not ( n3707 , n946 );
and ( n3708 , n3707 , n1013 );
not ( n3709 , n1013 );
and ( n3710 , n3699 , n3700 );
xor ( n3711 , n3709 , n3710 );
and ( n3712 , n3711 , n946 );
or ( n3713 , n3708 , n3712 );
not ( n3714 , n3713 );
not ( n3715 , n3714 );
or ( n3716 , n3706 , n3715 );
not ( n3717 , n946 );
and ( n3718 , n3717 , n1007 );
not ( n3719 , n1007 );
and ( n3720 , n3709 , n3710 );
xor ( n3721 , n3719 , n3720 );
and ( n3722 , n3721 , n946 );
or ( n3723 , n3718 , n3722 );
not ( n3724 , n3723 );
not ( n3725 , n3724 );
or ( n3726 , n3716 , n3725 );
not ( n3727 , n946 );
and ( n3728 , n3727 , n1001 );
not ( n3729 , n1001 );
and ( n3730 , n3719 , n3720 );
xor ( n3731 , n3729 , n3730 );
and ( n3732 , n3731 , n946 );
or ( n3733 , n3728 , n3732 );
not ( n3734 , n3733 );
not ( n3735 , n3734 );
or ( n3736 , n3726 , n3735 );
not ( n3737 , n946 );
and ( n3738 , n3737 , n995 );
not ( n3739 , n995 );
and ( n3740 , n3729 , n3730 );
xor ( n3741 , n3739 , n3740 );
and ( n3742 , n3741 , n946 );
or ( n3743 , n3738 , n3742 );
not ( n3744 , n3743 );
not ( n3745 , n3744 );
or ( n3746 , n3736 , n3745 );
not ( n3747 , n946 );
and ( n3748 , n3747 , n989 );
not ( n3749 , n989 );
and ( n3750 , n3739 , n3740 );
xor ( n3751 , n3749 , n3750 );
and ( n3752 , n3751 , n946 );
or ( n3753 , n3748 , n3752 );
not ( n3754 , n3753 );
not ( n3755 , n3754 );
or ( n3756 , n3746 , n3755 );
not ( n3757 , n946 );
and ( n3758 , n3757 , n983 );
not ( n3759 , n983 );
and ( n3760 , n3749 , n3750 );
xor ( n3761 , n3759 , n3760 );
and ( n3762 , n3761 , n946 );
or ( n3763 , n3758 , n3762 );
not ( n3764 , n3763 );
not ( n3765 , n3764 );
or ( n3766 , n3756 , n3765 );
not ( n3767 , n946 );
and ( n3768 , n3767 , n977 );
not ( n3769 , n977 );
and ( n3770 , n3759 , n3760 );
xor ( n3771 , n3769 , n3770 );
and ( n3772 , n3771 , n946 );
or ( n3773 , n3768 , n3772 );
not ( n3774 , n3773 );
not ( n3775 , n3774 );
or ( n3776 , n3766 , n3775 );
and ( n3777 , n3776 , n946 );
not ( n3778 , n3777 );
and ( n3779 , n3778 , n3586 );
xor ( n3780 , n3586 , n946 );
xor ( n3781 , n3780 , n946 );
and ( n3782 , n3781 , n3777 );
or ( n3783 , n3779 , n3782 );
and ( n3784 , n3783 , n3493 );
or ( n3785 , n3584 , n3784 );
xor ( n3786 , n1850 , n3785 );
not ( n3787 , n3786 );
not ( n3788 , n3787 );
buf ( n3789 , n654 );
and ( n3790 , n3789 , n3583 );
not ( n3791 , n3790 );
xor ( n3792 , n1859 , n3791 );
buf ( n3793 , n655 );
and ( n3794 , n3793 , n3583 );
not ( n3795 , n3794 );
and ( n3796 , n2717 , n3795 );
buf ( n3797 , n656 );
and ( n3798 , n3797 , n3583 );
not ( n3799 , n3798 );
and ( n3800 , n2728 , n3799 );
buf ( n3801 , n657 );
and ( n3802 , n3801 , n3583 );
not ( n3803 , n3802 );
and ( n3804 , n2515 , n3803 );
buf ( n3805 , n658 );
and ( n3806 , n3805 , n3583 );
not ( n3807 , n3806 );
and ( n3808 , n2491 , n3807 );
buf ( n3809 , n659 );
and ( n3810 , n3809 , n3583 );
not ( n3811 , n3810 );
and ( n3812 , n2467 , n3811 );
buf ( n3813 , n660 );
and ( n3814 , n3813 , n3583 );
not ( n3815 , n3814 );
and ( n3816 , n2443 , n3815 );
buf ( n3817 , n661 );
and ( n3818 , n3817 , n3583 );
not ( n3819 , n3818 );
and ( n3820 , n2419 , n3819 );
buf ( n3821 , n662 );
and ( n3822 , n3821 , n3583 );
not ( n3823 , n3822 );
and ( n3824 , n2395 , n3823 );
buf ( n3825 , n663 );
and ( n3826 , n3825 , n3583 );
not ( n3827 , n3826 );
and ( n3828 , n2371 , n3827 );
buf ( n3829 , n664 );
and ( n3830 , n3829 , n3583 );
not ( n3831 , n3830 );
and ( n3832 , n2347 , n3831 );
buf ( n3833 , n665 );
and ( n3834 , n3833 , n3583 );
not ( n3835 , n3834 );
and ( n3836 , n2323 , n3835 );
buf ( n3837 , n666 );
and ( n3838 , n3837 , n3583 );
not ( n3839 , n3777 );
and ( n3840 , n3839 , n3775 );
xor ( n3841 , n3775 , n946 );
xor ( n3842 , n3765 , n946 );
xor ( n3843 , n3755 , n946 );
xor ( n3844 , n3745 , n946 );
xor ( n3845 , n3735 , n946 );
xor ( n3846 , n3725 , n946 );
xor ( n3847 , n3715 , n946 );
xor ( n3848 , n3705 , n946 );
xor ( n3849 , n3695 , n946 );
xor ( n3850 , n3685 , n946 );
xor ( n3851 , n3675 , n946 );
xor ( n3852 , n3665 , n946 );
xor ( n3853 , n3655 , n946 );
xor ( n3854 , n3645 , n946 );
xor ( n3855 , n3635 , n946 );
xor ( n3856 , n3625 , n946 );
xor ( n3857 , n3615 , n946 );
xor ( n3858 , n3605 , n946 );
xor ( n3859 , n3595 , n946 );
and ( n3860 , n3780 , n946 );
and ( n3861 , n3859 , n3860 );
and ( n3862 , n3858 , n3861 );
and ( n3863 , n3857 , n3862 );
and ( n3864 , n3856 , n3863 );
and ( n3865 , n3855 , n3864 );
and ( n3866 , n3854 , n3865 );
and ( n3867 , n3853 , n3866 );
and ( n3868 , n3852 , n3867 );
and ( n3869 , n3851 , n3868 );
and ( n3870 , n3850 , n3869 );
and ( n3871 , n3849 , n3870 );
and ( n3872 , n3848 , n3871 );
and ( n3873 , n3847 , n3872 );
and ( n3874 , n3846 , n3873 );
and ( n3875 , n3845 , n3874 );
and ( n3876 , n3844 , n3875 );
and ( n3877 , n3843 , n3876 );
and ( n3878 , n3842 , n3877 );
xor ( n3879 , n3841 , n3878 );
and ( n3880 , n3879 , n3777 );
or ( n3881 , n3840 , n3880 );
and ( n3882 , n3881 , n3493 );
or ( n3883 , n3838 , n3882 );
not ( n3884 , n3883 );
and ( n3885 , n2299 , n3884 );
buf ( n3886 , n667 );
and ( n3887 , n3886 , n3583 );
not ( n3888 , n3777 );
and ( n3889 , n3888 , n3765 );
xor ( n3890 , n3842 , n3877 );
and ( n3891 , n3890 , n3777 );
or ( n3892 , n3889 , n3891 );
and ( n3893 , n3892 , n3493 );
or ( n3894 , n3887 , n3893 );
not ( n3895 , n3894 );
and ( n3896 , n2275 , n3895 );
buf ( n3897 , n668 );
and ( n3898 , n3897 , n3583 );
not ( n3899 , n3777 );
and ( n3900 , n3899 , n3755 );
xor ( n3901 , n3843 , n3876 );
and ( n3902 , n3901 , n3777 );
or ( n3903 , n3900 , n3902 );
and ( n3904 , n3903 , n3493 );
or ( n3905 , n3898 , n3904 );
not ( n3906 , n3905 );
and ( n3907 , n2251 , n3906 );
buf ( n3908 , n669 );
and ( n3909 , n3908 , n3583 );
not ( n3910 , n3777 );
and ( n3911 , n3910 , n3745 );
xor ( n3912 , n3844 , n3875 );
and ( n3913 , n3912 , n3777 );
or ( n3914 , n3911 , n3913 );
and ( n3915 , n3914 , n3493 );
or ( n3916 , n3909 , n3915 );
not ( n3917 , n3916 );
and ( n3918 , n2227 , n3917 );
buf ( n3919 , n670 );
and ( n3920 , n3919 , n3583 );
not ( n3921 , n3777 );
and ( n3922 , n3921 , n3735 );
xor ( n3923 , n3845 , n3874 );
and ( n3924 , n3923 , n3777 );
or ( n3925 , n3922 , n3924 );
and ( n3926 , n3925 , n3493 );
or ( n3927 , n3920 , n3926 );
not ( n3928 , n3927 );
and ( n3929 , n2203 , n3928 );
buf ( n3930 , n671 );
and ( n3931 , n3930 , n3583 );
not ( n3932 , n3777 );
and ( n3933 , n3932 , n3725 );
xor ( n3934 , n3846 , n3873 );
and ( n3935 , n3934 , n3777 );
or ( n3936 , n3933 , n3935 );
and ( n3937 , n3936 , n3493 );
or ( n3938 , n3931 , n3937 );
not ( n3939 , n3938 );
and ( n3940 , n2179 , n3939 );
buf ( n3941 , n672 );
and ( n3942 , n3941 , n3583 );
not ( n3943 , n3777 );
and ( n3944 , n3943 , n3715 );
xor ( n3945 , n3847 , n3872 );
and ( n3946 , n3945 , n3777 );
or ( n3947 , n3944 , n3946 );
and ( n3948 , n3947 , n3493 );
or ( n3949 , n3942 , n3948 );
not ( n3950 , n3949 );
and ( n3951 , n2155 , n3950 );
buf ( n3952 , n673 );
and ( n3953 , n3952 , n3583 );
not ( n3954 , n3777 );
and ( n3955 , n3954 , n3705 );
xor ( n3956 , n3848 , n3871 );
and ( n3957 , n3956 , n3777 );
or ( n3958 , n3955 , n3957 );
and ( n3959 , n3958 , n3493 );
or ( n3960 , n3953 , n3959 );
not ( n3961 , n3960 );
and ( n3962 , n2131 , n3961 );
buf ( n3963 , n674 );
and ( n3964 , n3963 , n3583 );
not ( n3965 , n3777 );
and ( n3966 , n3965 , n3695 );
xor ( n3967 , n3849 , n3870 );
and ( n3968 , n3967 , n3777 );
or ( n3969 , n3966 , n3968 );
and ( n3970 , n3969 , n3493 );
or ( n3971 , n3964 , n3970 );
not ( n3972 , n3971 );
and ( n3973 , n2107 , n3972 );
buf ( n3974 , n675 );
and ( n3975 , n3974 , n3583 );
not ( n3976 , n3777 );
and ( n3977 , n3976 , n3685 );
xor ( n3978 , n3850 , n3869 );
and ( n3979 , n3978 , n3777 );
or ( n3980 , n3977 , n3979 );
and ( n3981 , n3980 , n3493 );
or ( n3982 , n3975 , n3981 );
not ( n3983 , n3982 );
and ( n3984 , n2083 , n3983 );
buf ( n3985 , n676 );
and ( n3986 , n3985 , n3583 );
not ( n3987 , n3777 );
and ( n3988 , n3987 , n3675 );
xor ( n3989 , n3851 , n3868 );
and ( n3990 , n3989 , n3777 );
or ( n3991 , n3988 , n3990 );
and ( n3992 , n3991 , n3493 );
or ( n3993 , n3986 , n3992 );
not ( n3994 , n3993 );
and ( n3995 , n2059 , n3994 );
buf ( n3996 , n677 );
and ( n3997 , n3996 , n3583 );
not ( n3998 , n3777 );
and ( n3999 , n3998 , n3665 );
xor ( n4000 , n3852 , n3867 );
and ( n4001 , n4000 , n3777 );
or ( n4002 , n3999 , n4001 );
and ( n4003 , n4002 , n3493 );
or ( n4004 , n3997 , n4003 );
not ( n4005 , n4004 );
and ( n4006 , n2035 , n4005 );
buf ( n4007 , n678 );
and ( n4008 , n4007 , n3583 );
not ( n4009 , n3777 );
and ( n4010 , n4009 , n3655 );
xor ( n4011 , n3853 , n3866 );
and ( n4012 , n4011 , n3777 );
or ( n4013 , n4010 , n4012 );
and ( n4014 , n4013 , n3493 );
or ( n4015 , n4008 , n4014 );
not ( n4016 , n4015 );
and ( n4017 , n2011 , n4016 );
buf ( n4018 , n679 );
and ( n4019 , n4018 , n3583 );
not ( n4020 , n3777 );
and ( n4021 , n4020 , n3645 );
xor ( n4022 , n3854 , n3865 );
and ( n4023 , n4022 , n3777 );
or ( n4024 , n4021 , n4023 );
and ( n4025 , n4024 , n3493 );
or ( n4026 , n4019 , n4025 );
not ( n4027 , n4026 );
and ( n4028 , n1987 , n4027 );
buf ( n4029 , n680 );
and ( n4030 , n4029 , n3583 );
not ( n4031 , n3777 );
and ( n4032 , n4031 , n3635 );
xor ( n4033 , n3855 , n3864 );
and ( n4034 , n4033 , n3777 );
or ( n4035 , n4032 , n4034 );
and ( n4036 , n4035 , n3493 );
or ( n4037 , n4030 , n4036 );
not ( n4038 , n4037 );
and ( n4039 , n1963 , n4038 );
buf ( n4040 , n681 );
and ( n4041 , n4040 , n3583 );
not ( n4042 , n3777 );
and ( n4043 , n4042 , n3625 );
xor ( n4044 , n3856 , n3863 );
and ( n4045 , n4044 , n3777 );
or ( n4046 , n4043 , n4045 );
and ( n4047 , n4046 , n3493 );
or ( n4048 , n4041 , n4047 );
not ( n4049 , n4048 );
and ( n4050 , n1939 , n4049 );
buf ( n4051 , n682 );
and ( n4052 , n4051 , n3583 );
not ( n4053 , n3777 );
and ( n4054 , n4053 , n3615 );
xor ( n4055 , n3857 , n3862 );
and ( n4056 , n4055 , n3777 );
or ( n4057 , n4054 , n4056 );
and ( n4058 , n4057 , n3493 );
or ( n4059 , n4052 , n4058 );
not ( n4060 , n4059 );
and ( n4061 , n1915 , n4060 );
buf ( n4062 , n683 );
and ( n4063 , n4062 , n3583 );
not ( n4064 , n3777 );
and ( n4065 , n4064 , n3605 );
xor ( n4066 , n3858 , n3861 );
and ( n4067 , n4066 , n3777 );
or ( n4068 , n4065 , n4067 );
and ( n4069 , n4068 , n3493 );
or ( n4070 , n4063 , n4069 );
not ( n4071 , n4070 );
and ( n4072 , n1891 , n4071 );
buf ( n4073 , n684 );
and ( n4074 , n4073 , n3583 );
not ( n4075 , n3777 );
and ( n4076 , n4075 , n3595 );
xor ( n4077 , n3859 , n3860 );
and ( n4078 , n4077 , n3777 );
or ( n4079 , n4076 , n4078 );
and ( n4080 , n4079 , n3493 );
or ( n4081 , n4074 , n4080 );
not ( n4082 , n4081 );
and ( n4083 , n1868 , n4082 );
not ( n4084 , n3785 );
or ( n4085 , n1850 , n4084 );
and ( n4086 , n4082 , n4085 );
and ( n4087 , n1868 , n4085 );
or ( n4088 , n4083 , n4086 , n4087 );
and ( n4089 , n4071 , n4088 );
and ( n4090 , n1891 , n4088 );
or ( n4091 , n4072 , n4089 , n4090 );
and ( n4092 , n4060 , n4091 );
and ( n4093 , n1915 , n4091 );
or ( n4094 , n4061 , n4092 , n4093 );
and ( n4095 , n4049 , n4094 );
and ( n4096 , n1939 , n4094 );
or ( n4097 , n4050 , n4095 , n4096 );
and ( n4098 , n4038 , n4097 );
and ( n4099 , n1963 , n4097 );
or ( n4100 , n4039 , n4098 , n4099 );
and ( n4101 , n4027 , n4100 );
and ( n4102 , n1987 , n4100 );
or ( n4103 , n4028 , n4101 , n4102 );
and ( n4104 , n4016 , n4103 );
and ( n4105 , n2011 , n4103 );
or ( n4106 , n4017 , n4104 , n4105 );
and ( n4107 , n4005 , n4106 );
and ( n4108 , n2035 , n4106 );
or ( n4109 , n4006 , n4107 , n4108 );
and ( n4110 , n3994 , n4109 );
and ( n4111 , n2059 , n4109 );
or ( n4112 , n3995 , n4110 , n4111 );
and ( n4113 , n3983 , n4112 );
and ( n4114 , n2083 , n4112 );
or ( n4115 , n3984 , n4113 , n4114 );
and ( n4116 , n3972 , n4115 );
and ( n4117 , n2107 , n4115 );
or ( n4118 , n3973 , n4116 , n4117 );
and ( n4119 , n3961 , n4118 );
and ( n4120 , n2131 , n4118 );
or ( n4121 , n3962 , n4119 , n4120 );
and ( n4122 , n3950 , n4121 );
and ( n4123 , n2155 , n4121 );
or ( n4124 , n3951 , n4122 , n4123 );
and ( n4125 , n3939 , n4124 );
and ( n4126 , n2179 , n4124 );
or ( n4127 , n3940 , n4125 , n4126 );
and ( n4128 , n3928 , n4127 );
and ( n4129 , n2203 , n4127 );
or ( n4130 , n3929 , n4128 , n4129 );
and ( n4131 , n3917 , n4130 );
and ( n4132 , n2227 , n4130 );
or ( n4133 , n3918 , n4131 , n4132 );
and ( n4134 , n3906 , n4133 );
and ( n4135 , n2251 , n4133 );
or ( n4136 , n3907 , n4134 , n4135 );
and ( n4137 , n3895 , n4136 );
and ( n4138 , n2275 , n4136 );
or ( n4139 , n3896 , n4137 , n4138 );
and ( n4140 , n3884 , n4139 );
and ( n4141 , n2299 , n4139 );
or ( n4142 , n3885 , n4140 , n4141 );
and ( n4143 , n3835 , n4142 );
and ( n4144 , n2323 , n4142 );
or ( n4145 , n3836 , n4143 , n4144 );
and ( n4146 , n3831 , n4145 );
and ( n4147 , n2347 , n4145 );
or ( n4148 , n3832 , n4146 , n4147 );
and ( n4149 , n3827 , n4148 );
and ( n4150 , n2371 , n4148 );
or ( n4151 , n3828 , n4149 , n4150 );
and ( n4152 , n3823 , n4151 );
and ( n4153 , n2395 , n4151 );
or ( n4154 , n3824 , n4152 , n4153 );
and ( n4155 , n3819 , n4154 );
and ( n4156 , n2419 , n4154 );
or ( n4157 , n3820 , n4155 , n4156 );
and ( n4158 , n3815 , n4157 );
and ( n4159 , n2443 , n4157 );
or ( n4160 , n3816 , n4158 , n4159 );
and ( n4161 , n3811 , n4160 );
and ( n4162 , n2467 , n4160 );
or ( n4163 , n3812 , n4161 , n4162 );
and ( n4164 , n3807 , n4163 );
and ( n4165 , n2491 , n4163 );
or ( n4166 , n3808 , n4164 , n4165 );
and ( n4167 , n3803 , n4166 );
and ( n4168 , n2515 , n4166 );
or ( n4169 , n3804 , n4167 , n4168 );
and ( n4170 , n3799 , n4169 );
and ( n4171 , n2728 , n4169 );
or ( n4172 , n3800 , n4170 , n4171 );
and ( n4173 , n3795 , n4172 );
and ( n4174 , n2717 , n4172 );
or ( n4175 , n3796 , n4173 , n4174 );
xor ( n4176 , n3792 , n4175 );
not ( n4177 , n4176 );
xor ( n4178 , n1868 , n4082 );
xor ( n4179 , n4178 , n4085 );
and ( n4180 , n4177 , n4179 );
not ( n4181 , n4179 );
not ( n4182 , n3786 );
xor ( n4183 , n4181 , n4182 );
and ( n4184 , n4183 , n4176 );
or ( n4185 , n4180 , n4184 );
not ( n4186 , n4185 );
not ( n4187 , n4186 );
or ( n4188 , n3788 , n4187 );
not ( n4189 , n4176 );
xor ( n4190 , n1891 , n4071 );
xor ( n4191 , n4190 , n4088 );
and ( n4192 , n4189 , n4191 );
not ( n4193 , n4191 );
and ( n4194 , n4181 , n4182 );
xor ( n4195 , n4193 , n4194 );
and ( n4196 , n4195 , n4176 );
or ( n4197 , n4192 , n4196 );
not ( n4198 , n4197 );
not ( n4199 , n4198 );
or ( n4200 , n4188 , n4199 );
not ( n4201 , n4176 );
xor ( n4202 , n1915 , n4060 );
xor ( n4203 , n4202 , n4091 );
and ( n4204 , n4201 , n4203 );
not ( n4205 , n4203 );
and ( n4206 , n4193 , n4194 );
xor ( n4207 , n4205 , n4206 );
and ( n4208 , n4207 , n4176 );
or ( n4209 , n4204 , n4208 );
not ( n4210 , n4209 );
not ( n4211 , n4210 );
or ( n4212 , n4200 , n4211 );
not ( n4213 , n4176 );
xor ( n4214 , n1939 , n4049 );
xor ( n4215 , n4214 , n4094 );
and ( n4216 , n4213 , n4215 );
not ( n4217 , n4215 );
and ( n4218 , n4205 , n4206 );
xor ( n4219 , n4217 , n4218 );
and ( n4220 , n4219 , n4176 );
or ( n4221 , n4216 , n4220 );
not ( n4222 , n4221 );
not ( n4223 , n4222 );
or ( n4224 , n4212 , n4223 );
not ( n4225 , n4176 );
xor ( n4226 , n1963 , n4038 );
xor ( n4227 , n4226 , n4097 );
and ( n4228 , n4225 , n4227 );
not ( n4229 , n4227 );
and ( n4230 , n4217 , n4218 );
xor ( n4231 , n4229 , n4230 );
and ( n4232 , n4231 , n4176 );
or ( n4233 , n4228 , n4232 );
not ( n4234 , n4233 );
not ( n4235 , n4234 );
or ( n4236 , n4224 , n4235 );
not ( n4237 , n4176 );
xor ( n4238 , n1987 , n4027 );
xor ( n4239 , n4238 , n4100 );
and ( n4240 , n4237 , n4239 );
not ( n4241 , n4239 );
and ( n4242 , n4229 , n4230 );
xor ( n4243 , n4241 , n4242 );
and ( n4244 , n4243 , n4176 );
or ( n4245 , n4240 , n4244 );
not ( n4246 , n4245 );
not ( n4247 , n4246 );
or ( n4248 , n4236 , n4247 );
not ( n4249 , n4176 );
xor ( n4250 , n2011 , n4016 );
xor ( n4251 , n4250 , n4103 );
and ( n4252 , n4249 , n4251 );
not ( n4253 , n4251 );
and ( n4254 , n4241 , n4242 );
xor ( n4255 , n4253 , n4254 );
and ( n4256 , n4255 , n4176 );
or ( n4257 , n4252 , n4256 );
not ( n4258 , n4257 );
not ( n4259 , n4258 );
or ( n4260 , n4248 , n4259 );
not ( n4261 , n4176 );
xor ( n4262 , n2035 , n4005 );
xor ( n4263 , n4262 , n4106 );
and ( n4264 , n4261 , n4263 );
not ( n4265 , n4263 );
and ( n4266 , n4253 , n4254 );
xor ( n4267 , n4265 , n4266 );
and ( n4268 , n4267 , n4176 );
or ( n4269 , n4264 , n4268 );
not ( n4270 , n4269 );
not ( n4271 , n4270 );
or ( n4272 , n4260 , n4271 );
not ( n4273 , n4176 );
xor ( n4274 , n2059 , n3994 );
xor ( n4275 , n4274 , n4109 );
and ( n4276 , n4273 , n4275 );
not ( n4277 , n4275 );
and ( n4278 , n4265 , n4266 );
xor ( n4279 , n4277 , n4278 );
and ( n4280 , n4279 , n4176 );
or ( n4281 , n4276 , n4280 );
not ( n4282 , n4281 );
not ( n4283 , n4282 );
or ( n4284 , n4272 , n4283 );
not ( n4285 , n4176 );
xor ( n4286 , n2083 , n3983 );
xor ( n4287 , n4286 , n4112 );
and ( n4288 , n4285 , n4287 );
not ( n4289 , n4287 );
and ( n4290 , n4277 , n4278 );
xor ( n4291 , n4289 , n4290 );
and ( n4292 , n4291 , n4176 );
or ( n4293 , n4288 , n4292 );
not ( n4294 , n4293 );
not ( n4295 , n4294 );
or ( n4296 , n4284 , n4295 );
not ( n4297 , n4176 );
xor ( n4298 , n2107 , n3972 );
xor ( n4299 , n4298 , n4115 );
and ( n4300 , n4297 , n4299 );
not ( n4301 , n4299 );
and ( n4302 , n4289 , n4290 );
xor ( n4303 , n4301 , n4302 );
and ( n4304 , n4303 , n4176 );
or ( n4305 , n4300 , n4304 );
not ( n4306 , n4305 );
not ( n4307 , n4306 );
or ( n4308 , n4296 , n4307 );
not ( n4309 , n4176 );
xor ( n4310 , n2131 , n3961 );
xor ( n4311 , n4310 , n4118 );
and ( n4312 , n4309 , n4311 );
not ( n4313 , n4311 );
and ( n4314 , n4301 , n4302 );
xor ( n4315 , n4313 , n4314 );
and ( n4316 , n4315 , n4176 );
or ( n4317 , n4312 , n4316 );
not ( n4318 , n4317 );
not ( n4319 , n4318 );
or ( n4320 , n4308 , n4319 );
not ( n4321 , n4176 );
xor ( n4322 , n2155 , n3950 );
xor ( n4323 , n4322 , n4121 );
and ( n4324 , n4321 , n4323 );
not ( n4325 , n4323 );
and ( n4326 , n4313 , n4314 );
xor ( n4327 , n4325 , n4326 );
and ( n4328 , n4327 , n4176 );
or ( n4329 , n4324 , n4328 );
not ( n4330 , n4329 );
not ( n4331 , n4330 );
or ( n4332 , n4320 , n4331 );
not ( n4333 , n4176 );
xor ( n4334 , n2179 , n3939 );
xor ( n4335 , n4334 , n4124 );
and ( n4336 , n4333 , n4335 );
not ( n4337 , n4335 );
and ( n4338 , n4325 , n4326 );
xor ( n4339 , n4337 , n4338 );
and ( n4340 , n4339 , n4176 );
or ( n4341 , n4336 , n4340 );
not ( n4342 , n4341 );
not ( n4343 , n4342 );
or ( n4344 , n4332 , n4343 );
not ( n4345 , n4176 );
xor ( n4346 , n2203 , n3928 );
xor ( n4347 , n4346 , n4127 );
and ( n4348 , n4345 , n4347 );
not ( n4349 , n4347 );
and ( n4350 , n4337 , n4338 );
xor ( n4351 , n4349 , n4350 );
and ( n4352 , n4351 , n4176 );
or ( n4353 , n4348 , n4352 );
not ( n4354 , n4353 );
not ( n4355 , n4354 );
or ( n4356 , n4344 , n4355 );
not ( n4357 , n4176 );
xor ( n4358 , n2227 , n3917 );
xor ( n4359 , n4358 , n4130 );
and ( n4360 , n4357 , n4359 );
not ( n4361 , n4359 );
and ( n4362 , n4349 , n4350 );
xor ( n4363 , n4361 , n4362 );
and ( n4364 , n4363 , n4176 );
or ( n4365 , n4360 , n4364 );
not ( n4366 , n4365 );
not ( n4367 , n4366 );
or ( n4368 , n4356 , n4367 );
not ( n4369 , n4176 );
xor ( n4370 , n2251 , n3906 );
xor ( n4371 , n4370 , n4133 );
and ( n4372 , n4369 , n4371 );
not ( n4373 , n4371 );
and ( n4374 , n4361 , n4362 );
xor ( n4375 , n4373 , n4374 );
and ( n4376 , n4375 , n4176 );
or ( n4377 , n4372 , n4376 );
not ( n4378 , n4377 );
not ( n4379 , n4378 );
or ( n4380 , n4368 , n4379 );
not ( n4381 , n4176 );
xor ( n4382 , n2275 , n3895 );
xor ( n4383 , n4382 , n4136 );
and ( n4384 , n4381 , n4383 );
not ( n4385 , n4383 );
and ( n4386 , n4373 , n4374 );
xor ( n4387 , n4385 , n4386 );
and ( n4388 , n4387 , n4176 );
or ( n4389 , n4384 , n4388 );
not ( n4390 , n4389 );
not ( n4391 , n4390 );
or ( n4392 , n4380 , n4391 );
not ( n4393 , n4176 );
xor ( n4394 , n2299 , n3884 );
xor ( n4395 , n4394 , n4139 );
and ( n4396 , n4393 , n4395 );
not ( n4397 , n4395 );
and ( n4398 , n4385 , n4386 );
xor ( n4399 , n4397 , n4398 );
and ( n4400 , n4399 , n4176 );
or ( n4401 , n4396 , n4400 );
not ( n4402 , n4401 );
not ( n4403 , n4402 );
or ( n4404 , n4392 , n4403 );
not ( n4405 , n4176 );
xor ( n4406 , n2323 , n3835 );
xor ( n4407 , n4406 , n4142 );
and ( n4408 , n4405 , n4407 );
not ( n4409 , n4407 );
and ( n4410 , n4397 , n4398 );
xor ( n4411 , n4409 , n4410 );
and ( n4412 , n4411 , n4176 );
or ( n4413 , n4408 , n4412 );
not ( n4414 , n4413 );
not ( n4415 , n4414 );
or ( n4416 , n4404 , n4415 );
not ( n4417 , n4176 );
xor ( n4418 , n2347 , n3831 );
xor ( n4419 , n4418 , n4145 );
and ( n4420 , n4417 , n4419 );
not ( n4421 , n4419 );
and ( n4422 , n4409 , n4410 );
xor ( n4423 , n4421 , n4422 );
and ( n4424 , n4423 , n4176 );
or ( n4425 , n4420 , n4424 );
not ( n4426 , n4425 );
not ( n4427 , n4426 );
or ( n4428 , n4416 , n4427 );
not ( n4429 , n4176 );
xor ( n4430 , n2371 , n3827 );
xor ( n4431 , n4430 , n4148 );
and ( n4432 , n4429 , n4431 );
not ( n4433 , n4431 );
and ( n4434 , n4421 , n4422 );
xor ( n4435 , n4433 , n4434 );
and ( n4436 , n4435 , n4176 );
or ( n4437 , n4432 , n4436 );
not ( n4438 , n4437 );
not ( n4439 , n4438 );
or ( n4440 , n4428 , n4439 );
not ( n4441 , n4176 );
xor ( n4442 , n2395 , n3823 );
xor ( n4443 , n4442 , n4151 );
and ( n4444 , n4441 , n4443 );
not ( n4445 , n4443 );
and ( n4446 , n4433 , n4434 );
xor ( n4447 , n4445 , n4446 );
and ( n4448 , n4447 , n4176 );
or ( n4449 , n4444 , n4448 );
not ( n4450 , n4449 );
not ( n4451 , n4450 );
or ( n4452 , n4440 , n4451 );
not ( n4453 , n4176 );
xor ( n4454 , n2419 , n3819 );
xor ( n4455 , n4454 , n4154 );
and ( n4456 , n4453 , n4455 );
not ( n4457 , n4455 );
and ( n4458 , n4445 , n4446 );
xor ( n4459 , n4457 , n4458 );
and ( n4460 , n4459 , n4176 );
or ( n4461 , n4456 , n4460 );
not ( n4462 , n4461 );
not ( n4463 , n4462 );
or ( n4464 , n4452 , n4463 );
not ( n4465 , n4176 );
xor ( n4466 , n2443 , n3815 );
xor ( n4467 , n4466 , n4157 );
and ( n4468 , n4465 , n4467 );
not ( n4469 , n4467 );
and ( n4470 , n4457 , n4458 );
xor ( n4471 , n4469 , n4470 );
and ( n4472 , n4471 , n4176 );
or ( n4473 , n4468 , n4472 );
not ( n4474 , n4473 );
not ( n4475 , n4474 );
or ( n4476 , n4464 , n4475 );
not ( n4477 , n4176 );
xor ( n4478 , n2467 , n3811 );
xor ( n4479 , n4478 , n4160 );
and ( n4480 , n4477 , n4479 );
not ( n4481 , n4479 );
and ( n4482 , n4469 , n4470 );
xor ( n4483 , n4481 , n4482 );
and ( n4484 , n4483 , n4176 );
or ( n4485 , n4480 , n4484 );
not ( n4486 , n4485 );
not ( n4487 , n4486 );
or ( n4488 , n4476 , n4487 );
not ( n4489 , n4176 );
xor ( n4490 , n2491 , n3807 );
xor ( n4491 , n4490 , n4163 );
and ( n4492 , n4489 , n4491 );
not ( n4493 , n4491 );
and ( n4494 , n4481 , n4482 );
xor ( n4495 , n4493 , n4494 );
and ( n4496 , n4495 , n4176 );
or ( n4497 , n4492 , n4496 );
not ( n4498 , n4497 );
not ( n4499 , n4498 );
or ( n4500 , n4488 , n4499 );
not ( n4501 , n4176 );
xor ( n4502 , n2515 , n3803 );
xor ( n4503 , n4502 , n4166 );
and ( n4504 , n4501 , n4503 );
not ( n4505 , n4503 );
and ( n4506 , n4493 , n4494 );
xor ( n4507 , n4505 , n4506 );
and ( n4508 , n4507 , n4176 );
or ( n4509 , n4504 , n4508 );
not ( n4510 , n4509 );
not ( n4511 , n4510 );
or ( n4512 , n4500 , n4511 );
not ( n4513 , n4176 );
xor ( n4514 , n2728 , n3799 );
xor ( n4515 , n4514 , n4169 );
and ( n4516 , n4513 , n4515 );
not ( n4517 , n4515 );
and ( n4518 , n4505 , n4506 );
xor ( n4519 , n4517 , n4518 );
and ( n4520 , n4519 , n4176 );
or ( n4521 , n4516 , n4520 );
not ( n4522 , n4521 );
not ( n4523 , n4522 );
or ( n4524 , n4512 , n4523 );
and ( n4525 , n4524 , n4176 );
not ( n4526 , n4525 );
and ( n4527 , n4526 , n4187 );
xor ( n4528 , n4187 , n4176 );
xor ( n4529 , n3788 , n4176 );
and ( n4530 , n4529 , n4176 );
xor ( n4531 , n4528 , n4530 );
and ( n4532 , n4531 , n4525 );
or ( n4533 , n4527 , n4532 );
and ( n4534 , n4533 , n3569 );
and ( n4535 , n1447 , n3576 );
or ( n4536 , n4534 , n4535 );
not ( n4537 , n1705 );
and ( n4538 , n1707 , n1690 , n1698 , n4537 );
and ( n4539 , n1683 , n1690 , n1698 , n4537 );
or ( n4540 , n4538 , n4539 );
nor ( n4541 , n1707 , n1690 , n1698 , n4537 );
or ( n4542 , n4540 , n4541 );
nor ( n4543 , n1707 , n1691 , n1698 , n4537 );
or ( n4544 , n4542 , n4543 );
and ( n4545 , n4536 , n4544 );
xor ( n4546 , n1850 , n3785 );
not ( n4547 , n4546 );
not ( n4548 , n4547 );
xor ( n4549 , n1859 , n3790 );
and ( n4550 , n2717 , n3794 );
and ( n4551 , n2728 , n3798 );
and ( n4552 , n2515 , n3802 );
and ( n4553 , n2491 , n3806 );
and ( n4554 , n2467 , n3810 );
and ( n4555 , n2443 , n3814 );
and ( n4556 , n2419 , n3818 );
and ( n4557 , n2395 , n3822 );
and ( n4558 , n2371 , n3826 );
and ( n4559 , n2347 , n3830 );
and ( n4560 , n2323 , n3834 );
and ( n4561 , n2299 , n3883 );
and ( n4562 , n2275 , n3894 );
and ( n4563 , n2251 , n3905 );
and ( n4564 , n2227 , n3916 );
and ( n4565 , n2203 , n3927 );
and ( n4566 , n2179 , n3938 );
and ( n4567 , n2155 , n3949 );
and ( n4568 , n2131 , n3960 );
and ( n4569 , n2107 , n3971 );
and ( n4570 , n2083 , n3982 );
and ( n4571 , n2059 , n3993 );
and ( n4572 , n2035 , n4004 );
and ( n4573 , n2011 , n4015 );
and ( n4574 , n1987 , n4026 );
and ( n4575 , n1963 , n4037 );
and ( n4576 , n1939 , n4048 );
and ( n4577 , n1915 , n4059 );
and ( n4578 , n1891 , n4070 );
and ( n4579 , n1868 , n4081 );
and ( n4580 , n1850 , n3785 );
and ( n4581 , n4081 , n4580 );
and ( n4582 , n1868 , n4580 );
or ( n4583 , n4579 , n4581 , n4582 );
and ( n4584 , n4070 , n4583 );
and ( n4585 , n1891 , n4583 );
or ( n4586 , n4578 , n4584 , n4585 );
and ( n4587 , n4059 , n4586 );
and ( n4588 , n1915 , n4586 );
or ( n4589 , n4577 , n4587 , n4588 );
and ( n4590 , n4048 , n4589 );
and ( n4591 , n1939 , n4589 );
or ( n4592 , n4576 , n4590 , n4591 );
and ( n4593 , n4037 , n4592 );
and ( n4594 , n1963 , n4592 );
or ( n4595 , n4575 , n4593 , n4594 );
and ( n4596 , n4026 , n4595 );
and ( n4597 , n1987 , n4595 );
or ( n4598 , n4574 , n4596 , n4597 );
and ( n4599 , n4015 , n4598 );
and ( n4600 , n2011 , n4598 );
or ( n4601 , n4573 , n4599 , n4600 );
and ( n4602 , n4004 , n4601 );
and ( n4603 , n2035 , n4601 );
or ( n4604 , n4572 , n4602 , n4603 );
and ( n4605 , n3993 , n4604 );
and ( n4606 , n2059 , n4604 );
or ( n4607 , n4571 , n4605 , n4606 );
and ( n4608 , n3982 , n4607 );
and ( n4609 , n2083 , n4607 );
or ( n4610 , n4570 , n4608 , n4609 );
and ( n4611 , n3971 , n4610 );
and ( n4612 , n2107 , n4610 );
or ( n4613 , n4569 , n4611 , n4612 );
and ( n4614 , n3960 , n4613 );
and ( n4615 , n2131 , n4613 );
or ( n4616 , n4568 , n4614 , n4615 );
and ( n4617 , n3949 , n4616 );
and ( n4618 , n2155 , n4616 );
or ( n4619 , n4567 , n4617 , n4618 );
and ( n4620 , n3938 , n4619 );
and ( n4621 , n2179 , n4619 );
or ( n4622 , n4566 , n4620 , n4621 );
and ( n4623 , n3927 , n4622 );
and ( n4624 , n2203 , n4622 );
or ( n4625 , n4565 , n4623 , n4624 );
and ( n4626 , n3916 , n4625 );
and ( n4627 , n2227 , n4625 );
or ( n4628 , n4564 , n4626 , n4627 );
and ( n4629 , n3905 , n4628 );
and ( n4630 , n2251 , n4628 );
or ( n4631 , n4563 , n4629 , n4630 );
and ( n4632 , n3894 , n4631 );
and ( n4633 , n2275 , n4631 );
or ( n4634 , n4562 , n4632 , n4633 );
and ( n4635 , n3883 , n4634 );
and ( n4636 , n2299 , n4634 );
or ( n4637 , n4561 , n4635 , n4636 );
and ( n4638 , n3834 , n4637 );
and ( n4639 , n2323 , n4637 );
or ( n4640 , n4560 , n4638 , n4639 );
and ( n4641 , n3830 , n4640 );
and ( n4642 , n2347 , n4640 );
or ( n4643 , n4559 , n4641 , n4642 );
and ( n4644 , n3826 , n4643 );
and ( n4645 , n2371 , n4643 );
or ( n4646 , n4558 , n4644 , n4645 );
and ( n4647 , n3822 , n4646 );
and ( n4648 , n2395 , n4646 );
or ( n4649 , n4557 , n4647 , n4648 );
and ( n4650 , n3818 , n4649 );
and ( n4651 , n2419 , n4649 );
or ( n4652 , n4556 , n4650 , n4651 );
and ( n4653 , n3814 , n4652 );
and ( n4654 , n2443 , n4652 );
or ( n4655 , n4555 , n4653 , n4654 );
and ( n4656 , n3810 , n4655 );
and ( n4657 , n2467 , n4655 );
or ( n4658 , n4554 , n4656 , n4657 );
and ( n4659 , n3806 , n4658 );
and ( n4660 , n2491 , n4658 );
or ( n4661 , n4553 , n4659 , n4660 );
and ( n4662 , n3802 , n4661 );
and ( n4663 , n2515 , n4661 );
or ( n4664 , n4552 , n4662 , n4663 );
and ( n4665 , n3798 , n4664 );
and ( n4666 , n2728 , n4664 );
or ( n4667 , n4551 , n4665 , n4666 );
and ( n4668 , n3794 , n4667 );
and ( n4669 , n2717 , n4667 );
or ( n4670 , n4550 , n4668 , n4669 );
xor ( n4671 , n4549 , n4670 );
not ( n4672 , n4671 );
xor ( n4673 , n1868 , n4081 );
xor ( n4674 , n4673 , n4580 );
and ( n4675 , n4672 , n4674 );
not ( n4676 , n4674 );
not ( n4677 , n4546 );
xor ( n4678 , n4676 , n4677 );
and ( n4679 , n4678 , n4671 );
or ( n4680 , n4675 , n4679 );
not ( n4681 , n4680 );
not ( n4682 , n4681 );
or ( n4683 , n4548 , n4682 );
not ( n4684 , n4671 );
xor ( n4685 , n1891 , n4070 );
xor ( n4686 , n4685 , n4583 );
and ( n4687 , n4684 , n4686 );
not ( n4688 , n4686 );
and ( n4689 , n4676 , n4677 );
xor ( n4690 , n4688 , n4689 );
and ( n4691 , n4690 , n4671 );
or ( n4692 , n4687 , n4691 );
not ( n4693 , n4692 );
not ( n4694 , n4693 );
or ( n4695 , n4683 , n4694 );
not ( n4696 , n4671 );
xor ( n4697 , n1915 , n4059 );
xor ( n4698 , n4697 , n4586 );
and ( n4699 , n4696 , n4698 );
not ( n4700 , n4698 );
and ( n4701 , n4688 , n4689 );
xor ( n4702 , n4700 , n4701 );
and ( n4703 , n4702 , n4671 );
or ( n4704 , n4699 , n4703 );
not ( n4705 , n4704 );
not ( n4706 , n4705 );
or ( n4707 , n4695 , n4706 );
not ( n4708 , n4671 );
xor ( n4709 , n1939 , n4048 );
xor ( n4710 , n4709 , n4589 );
and ( n4711 , n4708 , n4710 );
not ( n4712 , n4710 );
and ( n4713 , n4700 , n4701 );
xor ( n4714 , n4712 , n4713 );
and ( n4715 , n4714 , n4671 );
or ( n4716 , n4711 , n4715 );
not ( n4717 , n4716 );
not ( n4718 , n4717 );
or ( n4719 , n4707 , n4718 );
not ( n4720 , n4671 );
xor ( n4721 , n1963 , n4037 );
xor ( n4722 , n4721 , n4592 );
and ( n4723 , n4720 , n4722 );
not ( n4724 , n4722 );
and ( n4725 , n4712 , n4713 );
xor ( n4726 , n4724 , n4725 );
and ( n4727 , n4726 , n4671 );
or ( n4728 , n4723 , n4727 );
not ( n4729 , n4728 );
not ( n4730 , n4729 );
or ( n4731 , n4719 , n4730 );
not ( n4732 , n4671 );
xor ( n4733 , n1987 , n4026 );
xor ( n4734 , n4733 , n4595 );
and ( n4735 , n4732 , n4734 );
not ( n4736 , n4734 );
and ( n4737 , n4724 , n4725 );
xor ( n4738 , n4736 , n4737 );
and ( n4739 , n4738 , n4671 );
or ( n4740 , n4735 , n4739 );
not ( n4741 , n4740 );
not ( n4742 , n4741 );
or ( n4743 , n4731 , n4742 );
not ( n4744 , n4671 );
xor ( n4745 , n2011 , n4015 );
xor ( n4746 , n4745 , n4598 );
and ( n4747 , n4744 , n4746 );
not ( n4748 , n4746 );
and ( n4749 , n4736 , n4737 );
xor ( n4750 , n4748 , n4749 );
and ( n4751 , n4750 , n4671 );
or ( n4752 , n4747 , n4751 );
not ( n4753 , n4752 );
not ( n4754 , n4753 );
or ( n4755 , n4743 , n4754 );
not ( n4756 , n4671 );
xor ( n4757 , n2035 , n4004 );
xor ( n4758 , n4757 , n4601 );
and ( n4759 , n4756 , n4758 );
not ( n4760 , n4758 );
and ( n4761 , n4748 , n4749 );
xor ( n4762 , n4760 , n4761 );
and ( n4763 , n4762 , n4671 );
or ( n4764 , n4759 , n4763 );
not ( n4765 , n4764 );
not ( n4766 , n4765 );
or ( n4767 , n4755 , n4766 );
not ( n4768 , n4671 );
xor ( n4769 , n2059 , n3993 );
xor ( n4770 , n4769 , n4604 );
and ( n4771 , n4768 , n4770 );
not ( n4772 , n4770 );
and ( n4773 , n4760 , n4761 );
xor ( n4774 , n4772 , n4773 );
and ( n4775 , n4774 , n4671 );
or ( n4776 , n4771 , n4775 );
not ( n4777 , n4776 );
not ( n4778 , n4777 );
or ( n4779 , n4767 , n4778 );
not ( n4780 , n4671 );
xor ( n4781 , n2083 , n3982 );
xor ( n4782 , n4781 , n4607 );
and ( n4783 , n4780 , n4782 );
not ( n4784 , n4782 );
and ( n4785 , n4772 , n4773 );
xor ( n4786 , n4784 , n4785 );
and ( n4787 , n4786 , n4671 );
or ( n4788 , n4783 , n4787 );
not ( n4789 , n4788 );
not ( n4790 , n4789 );
or ( n4791 , n4779 , n4790 );
not ( n4792 , n4671 );
xor ( n4793 , n2107 , n3971 );
xor ( n4794 , n4793 , n4610 );
and ( n4795 , n4792 , n4794 );
not ( n4796 , n4794 );
and ( n4797 , n4784 , n4785 );
xor ( n4798 , n4796 , n4797 );
and ( n4799 , n4798 , n4671 );
or ( n4800 , n4795 , n4799 );
not ( n4801 , n4800 );
not ( n4802 , n4801 );
or ( n4803 , n4791 , n4802 );
not ( n4804 , n4671 );
xor ( n4805 , n2131 , n3960 );
xor ( n4806 , n4805 , n4613 );
and ( n4807 , n4804 , n4806 );
not ( n4808 , n4806 );
and ( n4809 , n4796 , n4797 );
xor ( n4810 , n4808 , n4809 );
and ( n4811 , n4810 , n4671 );
or ( n4812 , n4807 , n4811 );
not ( n4813 , n4812 );
not ( n4814 , n4813 );
or ( n4815 , n4803 , n4814 );
not ( n4816 , n4671 );
xor ( n4817 , n2155 , n3949 );
xor ( n4818 , n4817 , n4616 );
and ( n4819 , n4816 , n4818 );
not ( n4820 , n4818 );
and ( n4821 , n4808 , n4809 );
xor ( n4822 , n4820 , n4821 );
and ( n4823 , n4822 , n4671 );
or ( n4824 , n4819 , n4823 );
not ( n4825 , n4824 );
not ( n4826 , n4825 );
or ( n4827 , n4815 , n4826 );
not ( n4828 , n4671 );
xor ( n4829 , n2179 , n3938 );
xor ( n4830 , n4829 , n4619 );
and ( n4831 , n4828 , n4830 );
not ( n4832 , n4830 );
and ( n4833 , n4820 , n4821 );
xor ( n4834 , n4832 , n4833 );
and ( n4835 , n4834 , n4671 );
or ( n4836 , n4831 , n4835 );
not ( n4837 , n4836 );
not ( n4838 , n4837 );
or ( n4839 , n4827 , n4838 );
not ( n4840 , n4671 );
xor ( n4841 , n2203 , n3927 );
xor ( n4842 , n4841 , n4622 );
and ( n4843 , n4840 , n4842 );
not ( n4844 , n4842 );
and ( n4845 , n4832 , n4833 );
xor ( n4846 , n4844 , n4845 );
and ( n4847 , n4846 , n4671 );
or ( n4848 , n4843 , n4847 );
not ( n4849 , n4848 );
not ( n4850 , n4849 );
or ( n4851 , n4839 , n4850 );
not ( n4852 , n4671 );
xor ( n4853 , n2227 , n3916 );
xor ( n4854 , n4853 , n4625 );
and ( n4855 , n4852 , n4854 );
not ( n4856 , n4854 );
and ( n4857 , n4844 , n4845 );
xor ( n4858 , n4856 , n4857 );
and ( n4859 , n4858 , n4671 );
or ( n4860 , n4855 , n4859 );
not ( n4861 , n4860 );
not ( n4862 , n4861 );
or ( n4863 , n4851 , n4862 );
not ( n4864 , n4671 );
xor ( n4865 , n2251 , n3905 );
xor ( n4866 , n4865 , n4628 );
and ( n4867 , n4864 , n4866 );
not ( n4868 , n4866 );
and ( n4869 , n4856 , n4857 );
xor ( n4870 , n4868 , n4869 );
and ( n4871 , n4870 , n4671 );
or ( n4872 , n4867 , n4871 );
not ( n4873 , n4872 );
not ( n4874 , n4873 );
or ( n4875 , n4863 , n4874 );
not ( n4876 , n4671 );
xor ( n4877 , n2275 , n3894 );
xor ( n4878 , n4877 , n4631 );
and ( n4879 , n4876 , n4878 );
not ( n4880 , n4878 );
and ( n4881 , n4868 , n4869 );
xor ( n4882 , n4880 , n4881 );
and ( n4883 , n4882 , n4671 );
or ( n4884 , n4879 , n4883 );
not ( n4885 , n4884 );
not ( n4886 , n4885 );
or ( n4887 , n4875 , n4886 );
not ( n4888 , n4671 );
xor ( n4889 , n2299 , n3883 );
xor ( n4890 , n4889 , n4634 );
and ( n4891 , n4888 , n4890 );
not ( n4892 , n4890 );
and ( n4893 , n4880 , n4881 );
xor ( n4894 , n4892 , n4893 );
and ( n4895 , n4894 , n4671 );
or ( n4896 , n4891 , n4895 );
not ( n4897 , n4896 );
not ( n4898 , n4897 );
or ( n4899 , n4887 , n4898 );
not ( n4900 , n4671 );
xor ( n4901 , n2323 , n3834 );
xor ( n4902 , n4901 , n4637 );
and ( n4903 , n4900 , n4902 );
not ( n4904 , n4902 );
and ( n4905 , n4892 , n4893 );
xor ( n4906 , n4904 , n4905 );
and ( n4907 , n4906 , n4671 );
or ( n4908 , n4903 , n4907 );
not ( n4909 , n4908 );
not ( n4910 , n4909 );
or ( n4911 , n4899 , n4910 );
not ( n4912 , n4671 );
xor ( n4913 , n2347 , n3830 );
xor ( n4914 , n4913 , n4640 );
and ( n4915 , n4912 , n4914 );
not ( n4916 , n4914 );
and ( n4917 , n4904 , n4905 );
xor ( n4918 , n4916 , n4917 );
and ( n4919 , n4918 , n4671 );
or ( n4920 , n4915 , n4919 );
not ( n4921 , n4920 );
not ( n4922 , n4921 );
or ( n4923 , n4911 , n4922 );
not ( n4924 , n4671 );
xor ( n4925 , n2371 , n3826 );
xor ( n4926 , n4925 , n4643 );
and ( n4927 , n4924 , n4926 );
not ( n4928 , n4926 );
and ( n4929 , n4916 , n4917 );
xor ( n4930 , n4928 , n4929 );
and ( n4931 , n4930 , n4671 );
or ( n4932 , n4927 , n4931 );
not ( n4933 , n4932 );
not ( n4934 , n4933 );
or ( n4935 , n4923 , n4934 );
not ( n4936 , n4671 );
xor ( n4937 , n2395 , n3822 );
xor ( n4938 , n4937 , n4646 );
and ( n4939 , n4936 , n4938 );
not ( n4940 , n4938 );
and ( n4941 , n4928 , n4929 );
xor ( n4942 , n4940 , n4941 );
and ( n4943 , n4942 , n4671 );
or ( n4944 , n4939 , n4943 );
not ( n4945 , n4944 );
not ( n4946 , n4945 );
or ( n4947 , n4935 , n4946 );
not ( n4948 , n4671 );
xor ( n4949 , n2419 , n3818 );
xor ( n4950 , n4949 , n4649 );
and ( n4951 , n4948 , n4950 );
not ( n4952 , n4950 );
and ( n4953 , n4940 , n4941 );
xor ( n4954 , n4952 , n4953 );
and ( n4955 , n4954 , n4671 );
or ( n4956 , n4951 , n4955 );
not ( n4957 , n4956 );
not ( n4958 , n4957 );
or ( n4959 , n4947 , n4958 );
not ( n4960 , n4671 );
xor ( n4961 , n2443 , n3814 );
xor ( n4962 , n4961 , n4652 );
and ( n4963 , n4960 , n4962 );
not ( n4964 , n4962 );
and ( n4965 , n4952 , n4953 );
xor ( n4966 , n4964 , n4965 );
and ( n4967 , n4966 , n4671 );
or ( n4968 , n4963 , n4967 );
not ( n4969 , n4968 );
not ( n4970 , n4969 );
or ( n4971 , n4959 , n4970 );
not ( n4972 , n4671 );
xor ( n4973 , n2467 , n3810 );
xor ( n4974 , n4973 , n4655 );
and ( n4975 , n4972 , n4974 );
not ( n4976 , n4974 );
and ( n4977 , n4964 , n4965 );
xor ( n4978 , n4976 , n4977 );
and ( n4979 , n4978 , n4671 );
or ( n4980 , n4975 , n4979 );
not ( n4981 , n4980 );
not ( n4982 , n4981 );
or ( n4983 , n4971 , n4982 );
not ( n4984 , n4671 );
xor ( n4985 , n2491 , n3806 );
xor ( n4986 , n4985 , n4658 );
and ( n4987 , n4984 , n4986 );
not ( n4988 , n4986 );
and ( n4989 , n4976 , n4977 );
xor ( n4990 , n4988 , n4989 );
and ( n4991 , n4990 , n4671 );
or ( n4992 , n4987 , n4991 );
not ( n4993 , n4992 );
not ( n4994 , n4993 );
or ( n4995 , n4983 , n4994 );
not ( n4996 , n4671 );
xor ( n4997 , n2515 , n3802 );
xor ( n4998 , n4997 , n4661 );
and ( n4999 , n4996 , n4998 );
not ( n5000 , n4998 );
and ( n5001 , n4988 , n4989 );
xor ( n5002 , n5000 , n5001 );
and ( n5003 , n5002 , n4671 );
or ( n5004 , n4999 , n5003 );
not ( n5005 , n5004 );
not ( n5006 , n5005 );
or ( n5007 , n4995 , n5006 );
not ( n5008 , n4671 );
xor ( n5009 , n2728 , n3798 );
xor ( n5010 , n5009 , n4664 );
and ( n5011 , n5008 , n5010 );
not ( n5012 , n5010 );
and ( n5013 , n5000 , n5001 );
xor ( n5014 , n5012 , n5013 );
and ( n5015 , n5014 , n4671 );
or ( n5016 , n5011 , n5015 );
not ( n5017 , n5016 );
not ( n5018 , n5017 );
or ( n5019 , n5007 , n5018 );
and ( n5020 , n5019 , n4671 );
not ( n5021 , n5020 );
and ( n5022 , n5021 , n4682 );
xor ( n5023 , n4682 , n4671 );
xor ( n5024 , n4548 , n4671 );
and ( n5025 , n5024 , n4671 );
xor ( n5026 , n5023 , n5025 );
and ( n5027 , n5026 , n5020 );
or ( n5028 , n5022 , n5027 );
and ( n5029 , n5028 , n3569 );
and ( n5030 , n1447 , n3576 );
or ( n5031 , n5029 , n5030 );
and ( n5032 , n1707 , n1691 , n1698 , n4537 );
and ( n5033 , n1683 , n1691 , n1698 , n4537 );
or ( n5034 , n5032 , n5033 );
nor ( n5035 , n1683 , n1690 , n1698 , n4537 );
or ( n5036 , n5034 , n5035 );
nor ( n5037 , n1683 , n1691 , n1698 , n4537 );
or ( n5038 , n5036 , n5037 );
and ( n5039 , n5031 , n5038 );
and ( n5040 , n4081 , n3569 );
and ( n5041 , n1447 , n3576 );
or ( n5042 , n5040 , n5041 );
nor ( n5043 , n1683 , n1691 , n1698 , n1705 );
nor ( n5044 , n1707 , n1691 , n1698 , n1705 );
or ( n5045 , n5043 , n5044 );
and ( n5046 , n5042 , n5045 );
nor ( n5047 , n1707 , n1690 , n1698 , n1705 );
and ( n5048 , n4081 , n5047 );
not ( n5049 , n4081 );
not ( n5050 , n3785 );
xor ( n5051 , n5049 , n5050 );
and ( n5052 , n5051 , n3569 );
and ( n5053 , n1447 , n3576 );
or ( n5054 , n5052 , n5053 );
nor ( n5055 , n1683 , n1690 , n1698 , n1705 );
and ( n5056 , n5054 , n5055 );
or ( n5057 , n1712 , n3580 , n4545 , n5039 , n5046 , n5048 , n5056 );
and ( n5058 , n1442 , n5057 );
and ( n5059 , n1447 , n1441 );
or ( n5060 , n5058 , n5059 );
buf ( n5061 , n686 );
and ( n5062 , n5060 , n5061 );
not ( n5063 , n5061 );
and ( n5064 , n1443 , n5063 );
or ( n5065 , n5062 , n5064 );
buf ( n5066 , n5065 );
buf ( n5067 , n5066 );
buf ( n5068 , n653 );
buf ( n5069 , n5068 );
buf ( n5070 , n847 );
not ( n5071 , n1441 );
and ( n5072 , n1883 , n1711 );
not ( n5073 , n2525 );
and ( n5074 , n5073 , n1876 );
xor ( n5075 , n1876 , n1859 );
and ( n5076 , n2528 , n1859 );
xor ( n5077 , n5075 , n5076 );
and ( n5078 , n5077 , n2525 );
or ( n5079 , n5074 , n5078 );
and ( n5080 , n5079 , n2671 );
and ( n5081 , n5079 , n2674 );
not ( n5082 , n2676 );
and ( n5083 , n5082 , n3080 );
not ( n5084 , n3480 );
and ( n5085 , n5084 , n3088 );
xor ( n5086 , n3088 , n3064 );
and ( n5087 , n3483 , n3485 );
xor ( n5088 , n5086 , n5087 );
and ( n5089 , n5088 , n3480 );
or ( n5090 , n5085 , n5089 );
and ( n5091 , n5090 , n2676 );
or ( n5092 , n5083 , n5091 );
and ( n5093 , n5092 , n3491 );
and ( n5094 , n3080 , n3493 );
or ( n5095 , n5080 , n5081 , n5093 , n5094 );
and ( n5096 , n5095 , n3569 );
and ( n5097 , n1883 , n3576 );
or ( n5098 , n5096 , n5097 );
and ( n5099 , n5098 , n3579 );
not ( n5100 , n4525 );
and ( n5101 , n5100 , n4199 );
xor ( n5102 , n4199 , n4176 );
and ( n5103 , n4528 , n4530 );
xor ( n5104 , n5102 , n5103 );
and ( n5105 , n5104 , n4525 );
or ( n5106 , n5101 , n5105 );
and ( n5107 , n5106 , n3569 );
and ( n5108 , n1883 , n3576 );
or ( n5109 , n5107 , n5108 );
and ( n5110 , n5109 , n4544 );
not ( n5111 , n5020 );
and ( n5112 , n5111 , n4694 );
xor ( n5113 , n4694 , n4671 );
and ( n5114 , n5023 , n5025 );
xor ( n5115 , n5113 , n5114 );
and ( n5116 , n5115 , n5020 );
or ( n5117 , n5112 , n5116 );
and ( n5118 , n5117 , n3569 );
and ( n5119 , n1883 , n3576 );
or ( n5120 , n5118 , n5119 );
and ( n5121 , n5120 , n5038 );
and ( n5122 , n4070 , n3569 );
and ( n5123 , n1883 , n3576 );
or ( n5124 , n5122 , n5123 );
and ( n5125 , n5124 , n5045 );
and ( n5126 , n4070 , n5047 );
not ( n5127 , n4070 );
and ( n5128 , n5049 , n5050 );
xor ( n5129 , n5127 , n5128 );
and ( n5130 , n5129 , n3569 );
and ( n5131 , n1883 , n3576 );
or ( n5132 , n5130 , n5131 );
and ( n5133 , n5132 , n5055 );
or ( n5134 , n5072 , n5099 , n5110 , n5121 , n5125 , n5126 , n5133 );
and ( n5135 , n5071 , n5134 );
and ( n5136 , n1883 , n1441 );
or ( n5137 , n5135 , n5136 );
and ( n5138 , n5137 , n5061 );
and ( n5139 , n1879 , n5063 );
or ( n5140 , n5138 , n5139 );
buf ( n5141 , n5140 );
buf ( n5142 , n5141 );
buf ( n5143 , n5068 );
buf ( n5144 , n847 );
not ( n5145 , n1441 );
and ( n5146 , n1907 , n1711 );
not ( n5147 , n2525 );
and ( n5148 , n5147 , n1899 );
xor ( n5149 , n1899 , n1859 );
and ( n5150 , n5075 , n5076 );
xor ( n5151 , n5149 , n5150 );
and ( n5152 , n5151 , n2525 );
or ( n5153 , n5148 , n5152 );
and ( n5154 , n5153 , n2671 );
and ( n5155 , n5153 , n2674 );
not ( n5156 , n2676 );
and ( n5157 , n5156 , n3095 );
not ( n5158 , n3480 );
and ( n5159 , n5158 , n3103 );
xor ( n5160 , n3103 , n3064 );
and ( n5161 , n5086 , n5087 );
xor ( n5162 , n5160 , n5161 );
and ( n5163 , n5162 , n3480 );
or ( n5164 , n5159 , n5163 );
and ( n5165 , n5164 , n2676 );
or ( n5166 , n5157 , n5165 );
and ( n5167 , n5166 , n3491 );
and ( n5168 , n3095 , n3493 );
or ( n5169 , n5154 , n5155 , n5167 , n5168 );
and ( n5170 , n5169 , n3569 );
and ( n5171 , n1907 , n3576 );
or ( n5172 , n5170 , n5171 );
and ( n5173 , n5172 , n3579 );
not ( n5174 , n4525 );
and ( n5175 , n5174 , n4211 );
xor ( n5176 , n4211 , n4176 );
and ( n5177 , n5102 , n5103 );
xor ( n5178 , n5176 , n5177 );
and ( n5179 , n5178 , n4525 );
or ( n5180 , n5175 , n5179 );
and ( n5181 , n5180 , n3569 );
and ( n5182 , n1907 , n3576 );
or ( n5183 , n5181 , n5182 );
and ( n5184 , n5183 , n4544 );
not ( n5185 , n5020 );
and ( n5186 , n5185 , n4706 );
xor ( n5187 , n4706 , n4671 );
and ( n5188 , n5113 , n5114 );
xor ( n5189 , n5187 , n5188 );
and ( n5190 , n5189 , n5020 );
or ( n5191 , n5186 , n5190 );
and ( n5192 , n5191 , n3569 );
and ( n5193 , n1907 , n3576 );
or ( n5194 , n5192 , n5193 );
and ( n5195 , n5194 , n5038 );
and ( n5196 , n4059 , n3569 );
and ( n5197 , n1907 , n3576 );
or ( n5198 , n5196 , n5197 );
and ( n5199 , n5198 , n5045 );
and ( n5200 , n4059 , n5047 );
not ( n5201 , n4059 );
and ( n5202 , n5127 , n5128 );
xor ( n5203 , n5201 , n5202 );
and ( n5204 , n5203 , n3569 );
and ( n5205 , n1907 , n3576 );
or ( n5206 , n5204 , n5205 );
and ( n5207 , n5206 , n5055 );
or ( n5208 , n5146 , n5173 , n5184 , n5195 , n5199 , n5200 , n5207 );
and ( n5209 , n5145 , n5208 );
and ( n5210 , n1907 , n1441 );
or ( n5211 , n5209 , n5210 );
and ( n5212 , n5211 , n5061 );
and ( n5213 , n1902 , n5063 );
or ( n5214 , n5212 , n5213 );
buf ( n5215 , n5214 );
buf ( n5216 , n5215 );
buf ( n5217 , n5068 );
buf ( n5218 , n847 );
not ( n5219 , n1441 );
and ( n5220 , n1931 , n1711 );
not ( n5221 , n2525 );
and ( n5222 , n5221 , n1923 );
xor ( n5223 , n1923 , n1859 );
and ( n5224 , n5149 , n5150 );
xor ( n5225 , n5223 , n5224 );
and ( n5226 , n5225 , n2525 );
or ( n5227 , n5222 , n5226 );
and ( n5228 , n5227 , n2671 );
and ( n5229 , n5227 , n2674 );
not ( n5230 , n2676 );
and ( n5231 , n5230 , n3110 );
not ( n5232 , n3480 );
and ( n5233 , n5232 , n3118 );
xor ( n5234 , n3118 , n3064 );
and ( n5235 , n5160 , n5161 );
xor ( n5236 , n5234 , n5235 );
and ( n5237 , n5236 , n3480 );
or ( n5238 , n5233 , n5237 );
and ( n5239 , n5238 , n2676 );
or ( n5240 , n5231 , n5239 );
and ( n5241 , n5240 , n3491 );
and ( n5242 , n3110 , n3493 );
or ( n5243 , n5228 , n5229 , n5241 , n5242 );
and ( n5244 , n5243 , n3569 );
and ( n5245 , n1931 , n3576 );
or ( n5246 , n5244 , n5245 );
and ( n5247 , n5246 , n3579 );
not ( n5248 , n4525 );
and ( n5249 , n5248 , n4223 );
xor ( n5250 , n4223 , n4176 );
and ( n5251 , n5176 , n5177 );
xor ( n5252 , n5250 , n5251 );
and ( n5253 , n5252 , n4525 );
or ( n5254 , n5249 , n5253 );
and ( n5255 , n5254 , n3569 );
and ( n5256 , n1931 , n3576 );
or ( n5257 , n5255 , n5256 );
and ( n5258 , n5257 , n4544 );
not ( n5259 , n5020 );
and ( n5260 , n5259 , n4718 );
xor ( n5261 , n4718 , n4671 );
and ( n5262 , n5187 , n5188 );
xor ( n5263 , n5261 , n5262 );
and ( n5264 , n5263 , n5020 );
or ( n5265 , n5260 , n5264 );
and ( n5266 , n5265 , n3569 );
and ( n5267 , n1931 , n3576 );
or ( n5268 , n5266 , n5267 );
and ( n5269 , n5268 , n5038 );
and ( n5270 , n4048 , n3569 );
and ( n5271 , n1931 , n3576 );
or ( n5272 , n5270 , n5271 );
and ( n5273 , n5272 , n5045 );
and ( n5274 , n4048 , n5047 );
not ( n5275 , n4048 );
and ( n5276 , n5201 , n5202 );
xor ( n5277 , n5275 , n5276 );
and ( n5278 , n5277 , n3569 );
and ( n5279 , n1931 , n3576 );
or ( n5280 , n5278 , n5279 );
and ( n5281 , n5280 , n5055 );
or ( n5282 , n5220 , n5247 , n5258 , n5269 , n5273 , n5274 , n5281 );
and ( n5283 , n5219 , n5282 );
and ( n5284 , n1931 , n1441 );
or ( n5285 , n5283 , n5284 );
and ( n5286 , n5285 , n5061 );
and ( n5287 , n1926 , n5063 );
or ( n5288 , n5286 , n5287 );
buf ( n5289 , n5288 );
buf ( n5290 , n5289 );
endmodule
