//
// Conformal-LEC Version 16.10-d005 ( 21-Apr-2016 ) ( 64 bit executable )
//
module top ( n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 );
input n0 , n1 , n2 , n3 , n4 , n5 , n6 , n7 , n8 , n9 , n10 , n11 , n12 , n13 , n14 , n15 , n16 , n17 , n18 , n19 , n20 , n21 , n22 , n23 , n24 , n25 , n26 , n27 , n28 , n29 , n30 , n31 , n32 , n33 , n34 , n35 , n36 , n37 , n38 , n39 , n40 , n41 , n42 , n43 , n44 , n45 , n46 , n47 , n48 , n49 , n50 , n51 , n52 , n53 , n54 , n55 , n56 , n57 , n58 , n59 , n60 , n61 , n62 , n63 , n64 , n65 , n66 , n67 , n68 , n69 , n70 , n71 , n72 , n73 , n74 , n75 , n76 , n77 , n78 , n79 , n80 , n81 , n82 , n83 , n84 , n85 , n86 , n87 , n88 , n89 , n90 , n91 , n92 , n93 , n94 , n95 , n96 , n97 , n98 , n99 , n100 , n101 , n102 , n103 , n104 , n105 , n106 , n107 , n108 , n109 , n110 , n111 , n112 , n113 , n114 , n115 , n116 , n117 , n118 , n119 , n120 , n121 , n122 , n123 , n124 , n125 , n126 , n127 , n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n136 , n137 , n138 , n139 , n140 , n141 , n142 , n143 , n144 , n145 , n146 , n147 , n148 , n149 , n150 , n151 , n152 , n153 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 , n163 , n164 , n165 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 , n174 , n175 , n176 , n177 , n178 , n179 , n180 , n181 , n182 , n183 , n184 , n185 , n186 , n187 , n188 , n189 , n190 , n191 ;
output n192 , n193 , n194 , n195 , n196 , n197 , n198 , n199 , n200 , n201 ;

wire n404 , n405 , n406 , n407 , n408 , n409 , n410 , n411 , n412 ,
     n413 , n414 , n415 , n416 , n417 , n418 , n419 , n420 , n421 , n422 ,
     n423 , n424 , n425 , n426 , n427 , n428 , n429 , n430 , n431 , n432 ,
     n433 , n434 , n435 , n436 , n437 , n438 , n439 , n440 , n441 , n442 ,
     n443 , n444 , n445 , n446 , n447 , n448 , n449 , n450 , n451 , n452 ,
     n453 , n454 , n455 , n456 , n457 , n458 , n459 , n460 , n461 , n462 ,
     n463 , n464 , n465 , n466 , n467 , n468 , n469 , n470 , n471 , n472 ,
     n473 , n474 , n475 , n476 , n477 , n478 , n479 , n480 , n481 , n482 ,
     n483 , n484 , n485 , n486 , n487 , n488 , n489 , n490 , n491 , n492 ,
     n493 , n494 , n495 , n496 , n497 , n498 , n499 , n500 , n501 , n502 ,
     n503 , n504 , n505 , n506 , n507 , n508 , n509 , n510 , n511 , n512 ,
     n513 , n514 , n515 , n516 , n517 , n518 , n519 , n520 , n521 , n522 ,
     n523 , n524 , n525 , n526 , n527 , n528 , n529 , n530 , n531 , n532 ,
     n533 , n534 , n535 , n536 , n537 , n538 , n539 , n540 , n541 , n542 ,
     n543 , n544 , n545 , n546 , n547 , n548 , n549 , n550 , n551 , n552 ,
     n553 , n554 , n555 , n556 , n557 , n558 , n559 , n560 , n561 , n562 ,
     n563 , n564 , n565 , n566 , n567 , n568 , n569 , n570 , n571 , n572 ,
     n573 , n574 , n575 , n576 , n577 , n578 , n579 , n580 , n581 , n582 ,
     n583 , n584 , n585 , n586 , n587 , n588 , n589 , n590 , n591 , n592 ,
     n593 , n594 , n595 , n596 , n597 , n598 , n599 , n600 , n601 , n602 ,
     n603 , n604 , n605 , n606 , n607 , n608 , n609 , n610 , n611 , n612 ,
     n613 , n614 , n615 , n616 , n617 , n618 , n619 , n620 , n621 , n622 ,
     n623 , n624 , n625 , n626 , n627 , n628 , n629 , n630 , n631 , n632 ,
     n633 , n634 , n635 , n636 , n637 , n638 , n639 , n640 , n641 , n642 ,
     n643 , n644 , n645 , n646 , n647 , n648 , n649 , n650 , n651 , n652 ,
     n653 , n654 , n655 , n656 , n657 , n658 , n659 , n660 , n661 , n662 ,
     n663 , n664 , n665 , n666 , n667 , n668 , n669 , n670 , n671 , n672 ,
     n673 , n674 , n675 , n676 , n677 , n678 , n679 , n680 , n681 , n682 ,
     n683 , n684 , n685 , n686 , n687 , n688 , n689 , n690 , n691 , n692 ,
     n693 , n694 , n695 , n696 , n697 , n698 , n699 , n700 , n701 , n702 ,
     n703 , n704 , n705 , n706 , n707 , n708 , n709 , n710 , n711 , n712 ,
     n713 , n714 , n715 , n716 , n717 , n718 , n719 , n720 , n721 , n722 ,
     n723 , n724 , n725 , n726 , n727 , n728 , n729 , n730 , n731 , n732 ,
     n733 , n734 , n735 , n736 , n737 , n738 , n739 , n740 , n741 , n742 ,
     n743 , n744 , n745 , n746 , n747 , n748 , n749 , n750 , n751 , n752 ,
     n753 , n754 , n755 , n756 , n757 , n758 , n759 , n760 , n761 , n762 ,
     n763 , n764 , n765 , n766 , n767 , n768 , n769 , n770 , n771 , n772 ,
     n773 , n774 , n775 , n776 , n777 , n778 , n779 , n780 , n781 , n782 ,
     n783 , n784 , n785 , n786 , n787 , n788 , n789 , n790 , n791 , n792 ,
     n793 , n794 , n795 , n796 , n797 , n798 , n799 , n800 , n801 , n802 ,
     n803 , n804 , n805 , n806 , n807 , n808 , n809 , n810 , n811 , n812 ,
     n813 , n814 , n815 , n816 , n817 , n818 , n819 , n820 , n821 , n822 ,
     n823 , n824 , n825 , n826 , n827 , n828 , n829 , n830 , n831 , n832 ,
     n833 , n834 , n835 , n836 , n837 , n838 , n839 , n840 , n841 , n842 ,
     n843 , n844 , n845 , n846 , n847 , n848 , n849 , n850 , n851 , n852 ,
     n853 , n854 , n855 , n856 , n857 , n858 , n859 , n860 , n861 , n862 ,
     n863 , n864 , n865 , n866 , n867 , n868 , n869 , n870 , n871 , n872 ,
     n873 , n874 , n875 , n876 , n877 , n878 , n879 , n880 , n881 , n882 ,
     n883 , n884 , n885 , n886 , n887 , n888 , n889 , n890 , n891 , n892 ,
     n893 , n894 , n895 , n896 , n897 , n898 , n899 , n900 , n901 , n902 ,
     n903 , n904 , n905 , n906 , n907 , n908 , n909 , n910 , n911 , n912 ,
     n913 , n914 , n915 , n916 , n917 , n918 , n919 , n920 , n921 , n922 ,
     n923 , n924 , n925 , n926 , n927 , n928 , n929 , n930 , n931 , n932 ,
     n933 , n934 , n935 , n936 , n937 , n938 , n939 , n940 , n941 , n942 ,
     n943 , n944 , n945 , n946 , n947 , n948 , n949 , n950 , n951 , n952 ,
     n953 , n954 , n955 , n956 , n957 , n958 , n959 , n960 , n961 , n962 ,
     n963 , n964 , n965 , n966 , n967 , n968 , n969 , n970 , n971 , n972 ,
     n973 , n974 , n975 , n976 , n977 , n978 , n979 , n980 , n981 , n982 ,
     n983 , n984 , n985 , n986 , n987 , n988 , n989 , n990 , n991 , n992 ,
     n993 , n994 , n995 , n996 , n997 , n998 , n999 , n1000 , n1001 , n1002 ,
     n1003 , n1004 , n1005 , n1006 , n1007 , n1008 , n1009 , n1010 , n1011 , n1012 ,
     n1013 , n1014 , n1015 , n1016 , n1017 , n1018 , n1019 , n1020 , n1021 , n1022 ,
     n1023 , n1024 , n1025 , n1026 , n1027 , n1028 , n1029 , n1030 , n1031 , n1032 ,
     n1033 , n1034 , n1035 , n1036 , n1037 , n1038 , n1039 , n1040 , n1041 , n1042 ,
     n1043 , n1044 , n1045 , n1046 , n1047 , n1048 , n1049 , n1050 , n1051 , n1052 ,
     n1053 , n1054 , n1055 , n1056 , n1057 , n1058 , n1059 , n1060 , n1061 , n1062 ,
     n1063 , n1064 , n1065 , n1066 , n1067 , n1068 , n1069 , n1070 , n1071 , n1072 ,
     n1073 , n1074 , n1075 , n1076 , n1077 , n1078 , n1079 , n1080 , n1081 , n1082 ,
     n1083 , n1084 , n1085 , n1086 , n1087 , n1088 , n1089 , n1090 , n1091 , n1092 ,
     n1093 , n1094 , n1095 , n1096 , n1097 , n1098 , n1099 , n1100 , n1101 , n1102 ,
     n1103 , n1104 , n1105 , n1106 , n1107 , n1108 , n1109 , n1110 , n1111 , n1112 ,
     n1113 , n1114 , n1115 , n1116 , n1117 , n1118 , n1119 , n1120 , n1121 , n1122 ,
     n1123 , n1124 , n1125 , n1126 , n1127 , n1128 , n1129 , n1130 , n1131 , n1132 ,
     n1133 , n1134 , n1135 , n1136 , n1137 , n1138 , n1139 , n1140 , n1141 , n1142 ,
     n1143 , n1144 , n1145 , n1146 , n1147 , n1148 , n1149 , n1150 , n1151 , n1152 ,
     n1153 , n1154 , n1155 , n1156 , n1157 , n1158 , n1159 , n1160 , n1161 , n1162 ,
     n1163 , n1164 , n1165 , n1166 , n1167 , n1168 , n1169 , n1170 , n1171 , n1172 ,
     n1173 , n1174 , n1175 , n1176 , n1177 , n1178 , n1179 , n1180 , n1181 , n1182 ,
     n1183 , n1184 , n1185 , n1186 , n1187 , n1188 , n1189 , n1190 , n1191 , n1192 ,
     n1193 , n1194 , n1195 , n1196 , n1197 , n1198 , n1199 , n1200 , n1201 , n1202 ,
     n1203 , n1204 , n1205 , n1206 , n1207 , n1208 , n1209 , n1210 , n1211 , n1212 ,
     n1213 , n1214 , n1215 , n1216 , n1217 , n1218 , n1219 , n1220 , n1221 , n1222 ,
     n1223 , n1224 , n1225 , n1226 , n1227 , n1228 , n1229 , n1230 , n1231 , n1232 ,
     n1233 , n1234 , n1235 , n1236 , n1237 , n1238 , n1239 , n1240 , n1241 , n1242 ,
     n1243 , n1244 , n1245 , n1246 , n1247 , n1248 , n1249 , n1250 , n1251 , n1252 ,
     n1253 , n1254 , n1255 , n1256 , n1257 , n1258 , n1259 , n1260 , n1261 , n1262 ,
     n1263 , n1264 , n1265 , n1266 , n1267 , n1268 , n1269 , n1270 , n1271 , n1272 ,
     n1273 , n1274 , n1275 , n1276 , n1277 , n1278 , n1279 , n1280 , n1281 , n1282 ,
     n1283 , n1284 , n1285 , n1286 , n1287 , n1288 , n1289 , n1290 , n1291 , n1292 ,
     n1293 , n1294 , n1295 , n1296 , n1297 , n1298 , n1299 , n1300 , n1301 , n1302 ,
     n1303 , n1304 , n1305 , n1306 , n1307 , n1308 , n1309 , n1310 , n1311 , n1312 ,
     n1313 , n1314 , n1315 , n1316 , n1317 , n1318 , n1319 , n1320 , n1321 , n1322 ,
     n1323 , n1324 , n1325 , n1326 , n1327 , n1328 , n1329 , n1330 , n1331 , n1332 ,
     n1333 , n1334 , n1335 , n1336 , n1337 , n1338 , n1339 , n1340 , n1341 , n1342 ,
     n1343 , n1344 , n1345 , n1346 , n1347 , n1348 , n1349 , n1350 , n1351 , n1352 ,
     n1353 , n1354 , n1355 , n1356 , n1357 , n1358 , n1359 , n1360 , n1361 , n1362 ,
     n1363 , n1364 , n1365 , n1366 , n1367 , n1368 , n1369 , n1370 , n1371 , n1372 ,
     n1373 , n1374 , n1375 , n1376 , n1377 , n1378 , n1379 , n1380 , n1381 , n1382 ,
     n1383 , n1384 , n1385 , n1386 , n1387 , n1388 , n1389 , n1390 , n1391 , n1392 ,
     n1393 , n1394 , n1395 , n1396 , n1397 , n1398 , n1399 , n1400 , n1401 , n1402 ,
     n1403 , n1404 , n1405 , n1406 , n1407 , n1408 , n1409 , n1410 , n1411 , n1412 ,
     n1413 , n1414 , n1415 , n1416 , n1417 , n1418 , n1419 , n1420 , n1421 , n1422 ,
     n1423 , n1424 , n1425 , n1426 , n1427 , n1428 , n1429 , n1430 , n1431 , n1432 ,
     n1433 , n1434 , n1435 , n1436 , n1437 , n1438 , n1439 , n1440 , n1441 , n1442 ,
     n1443 , n1444 , n1445 , n1446 , n1447 , n1448 , n1449 , n1450 , n1451 , n1452 ,
     n1453 , n1454 , n1455 , n1456 , n1457 , n1458 , n1459 , n1460 , n1461 , n1462 ,
     n1463 , n1464 , n1465 , n1466 , n1467 , n1468 , n1469 , n1470 , n1471 , n1472 ,
     n1473 , n1474 , n1475 , n1476 , n1477 , n1478 , n1479 , n1480 , n1481 , n1482 ,
     n1483 , n1484 , n1485 , n1486 , n1487 , n1488 , n1489 , n1490 , n1491 , n1492 ,
     n1493 , n1494 , n1495 , n1496 , n1497 , n1498 , n1499 , n1500 , n1501 , n1502 ,
     n1503 , n1504 , n1505 , n1506 , n1507 , n1508 , n1509 , n1510 , n1511 , n1512 ,
     n1513 , n1514 , n1515 , n1516 , n1517 , n1518 , n1519 , n1520 , n1521 , n1522 ,
     n1523 , n1524 , n1525 , n1526 , n1527 , n1528 , n1529 , n1530 , n1531 , n1532 ,
     n1533 , n1534 , n1535 , n1536 , n1537 , n1538 , n1539 , n1540 , n1541 , n1542 ,
     n1543 , n1544 , n1545 , n1546 , n1547 , n1548 , n1549 , n1550 , n1551 , n1552 ,
     n1553 , n1554 , n1555 , n1556 , n1557 , n1558 , n1559 , n1560 , n1561 , n1562 ,
     n1563 , n1564 , n1565 , n1566 , n1567 , n1568 , n1569 , n1570 , n1571 , n1572 ,
     n1573 , n1574 , n1575 , n1576 , n1577 , n1578 , n1579 , n1580 , n1581 , n1582 ,
     n1583 , n1584 , n1585 , n1586 , n1587 , n1588 , n1589 , n1590 , n1591 , n1592 ,
     n1593 , n1594 , n1595 , n1596 , n1597 , n1598 , n1599 , n1600 , n1601 , n1602 ,
     n1603 , n1604 , n1605 , n1606 , n1607 , n1608 , n1609 , n1610 , n1611 , n1612 ,
     n1613 , n1614 , n1615 , n1616 , n1617 , n1618 , n1619 , n1620 , n1621 , n1622 ,
     n1623 , n1624 , n1625 , n1626 , n1627 , n1628 , n1629 , n1630 , n1631 , n1632 ,
     n1633 , n1634 , n1635 , n1636 , n1637 , n1638 , n1639 , n1640 , n1641 , n1642 ,
     n1643 , n1644 , n1645 , n1646 , n1647 , n1648 , n1649 , n1650 , n1651 , n1652 ,
     n1653 , n1654 , n1655 , n1656 , n1657 , n1658 , n1659 , n1660 , n1661 , n1662 ,
     n1663 , n1664 , n1665 , n1666 , n1667 , n1668 , n1669 , n1670 , n1671 , n1672 ,
     n1673 , n1674 , n1675 , n1676 , n1677 , n1678 , n1679 , n1680 , n1681 , n1682 ,
     n1683 , n1684 , n1685 , n1686 , n1687 , n1688 , n1689 , n1690 , n1691 , n1692 ,
     n1693 , n1694 , n1695 , n1696 , n1697 , n1698 , n1699 , n1700 , n1701 , n1702 ,
     n1703 , n1704 , n1705 , n1706 , n1707 , n1708 , n1709 , n1710 , n1711 , n1712 ,
     n1713 , n1714 , n1715 , n1716 , n1717 , n1718 , n1719 , n1720 , n1721 , n1722 ,
     n1723 , n1724 , n1725 , n1726 , n1727 , n1728 , n1729 , n1730 , n1731 , n1732 ,
     n1733 , n1734 , n1735 , n1736 , n1737 , n1738 , n1739 , n1740 , n1741 , n1742 ,
     n1743 , n1744 , n1745 , n1746 , n1747 , n1748 , n1749 , n1750 , n1751 , n1752 ,
     n1753 , n1754 , n1755 , n1756 , n1757 , n1758 , n1759 , n1760 , n1761 , n1762 ,
     n1763 , n1764 , n1765 , n1766 , n1767 , n1768 , n1769 , n1770 , n1771 , n1772 ,
     n1773 , n1774 , n1775 , n1776 , n1777 , n1778 , n1779 , n1780 , n1781 , n1782 ,
     n1783 , n1784 , n1785 , n1786 , n1787 , n1788 , n1789 , n1790 , n1791 , n1792 ,
     n1793 , n1794 , n1795 , n1796 , n1797 , n1798 , n1799 , n1800 , n1801 , n1802 ,
     n1803 , n1804 , n1805 , n1806 , n1807 , n1808 , n1809 , n1810 , n1811 , n1812 ,
     n1813 , n1814 , n1815 , n1816 , n1817 , n1818 , n1819 , n1820 , n1821 , n1822 ,
     n1823 , n1824 , n1825 , n1826 , n1827 , n1828 , n1829 , n1830 , n1831 , n1832 ,
     n1833 , n1834 , n1835 , n1836 , n1837 , n1838 , n1839 , n1840 , n1841 , n1842 ,
     n1843 , n1844 , n1845 , n1846 , n1847 , n1848 , n1849 , n1850 , n1851 , n1852 ,
     n1853 , n1854 , n1855 , n1856 , n1857 , n1858 , n1859 , n1860 , n1861 , n1862 ,
     n1863 , n1864 , n1865 , n1866 , n1867 , n1868 , n1869 , n1870 , n1871 , n1872 ,
     n1873 , n1874 , n1875 , n1876 , n1877 , n1878 , n1879 , n1880 , n1881 , n1882 ,
     n1883 , n1884 , n1885 , n1886 , n1887 , n1888 , n1889 , n1890 , n1891 , n1892 ,
     n1893 , n1894 , n1895 , n1896 , n1897 , n1898 , n1899 , n1900 , n1901 , n1902 ,
     n1903 , n1904 , n1905 , n1906 , n1907 , n1908 , n1909 , n1910 , n1911 , n1912 ,
     n1913 , n1914 , n1915 , n1916 , n1917 , n1918 , n1919 , n1920 , n1921 , n1922 ,
     n1923 , n1924 , n1925 , n1926 , n1927 , n1928 , n1929 , n1930 , n1931 , n1932 ,
     n1933 , n1934 , n1935 , n1936 , n1937 , n1938 , n1939 , n1940 , n1941 , n1942 ,
     n1943 , n1944 , n1945 , n1946 , n1947 , n1948 , n1949 , n1950 , n1951 , n1952 ,
     n1953 , n1954 , n1955 , n1956 , n1957 , n1958 , n1959 , n1960 , n1961 , n1962 ,
     n1963 , n1964 , n1965 , n1966 , n1967 , n1968 , n1969 , n1970 , n1971 , n1972 ,
     n1973 , n1974 , n1975 , n1976 , n1977 , n1978 , n1979 , n1980 , n1981 , n1982 ,
     n1983 , n1984 , n1985 , n1986 , n1987 , n1988 , n1989 , n1990 , n1991 , n1992 ,
     n1993 , n1994 , n1995 , n1996 , n1997 , n1998 , n1999 , n2000 , n2001 , n2002 ,
     n2003 , n2004 , n2005 , n2006 , n2007 , n2008 , n2009 , n2010 , n2011 , n2012 ,
     n2013 , n2014 , n2015 , n2016 , n2017 , n2018 , n2019 , n2020 , n2021 , n2022 ,
     n2023 , n2024 , n2025 , n2026 , n2027 , n2028 , n2029 , n2030 , n2031 , n2032 ,
     n2033 , n2034 , n2035 , n2036 , n2037 , n2038 , n2039 , n2040 , n2041 , n2042 ,
     n2043 , n2044 , n2045 , n2046 , n2047 , n2048 , n2049 , n2050 , n2051 , n2052 ,
     n2053 , n2054 , n2055 , n2056 , n2057 , n2058 , n2059 , n2060 , n2061 , n2062 ,
     n2063 , n2064 , n2065 , n2066 , n2067 , n2068 , n2069 , n2070 , n2071 , n2072 ,
     n2073 , n2074 , n2075 , n2076 , n2077 , n2078 , n2079 , n2080 , n2081 , n2082 ,
     n2083 , n2084 , n2085 , n2086 , n2087 , n2088 , n2089 , n2090 , n2091 , n2092 ,
     n2093 , n2094 , n2095 , n2096 , n2097 , n2098 , n2099 , n2100 , n2101 , n2102 ,
     n2103 , n2104 , n2105 , n2106 , n2107 , n2108 , n2109 , n2110 , n2111 , n2112 ,
     n2113 , n2114 , n2115 , n2116 , n2117 , n2118 , n2119 , n2120 , n2121 , n2122 ,
     n2123 , n2124 , n2125 , n2126 , n2127 , n2128 , n2129 , n2130 , n2131 , n2132 ,
     n2133 , n2134 , n2135 , n2136 , n2137 , n2138 , n2139 , n2140 , n2141 , n2142 ,
     n2143 , n2144 , n2145 , n2146 , n2147 , n2148 , n2149 , n2150 , n2151 , n2152 ,
     n2153 , n2154 , n2155 , n2156 , n2157 , n2158 , n2159 , n2160 , n2161 , n2162 ,
     n2163 , n2164 , n2165 , n2166 , n2167 , n2168 , n2169 , n2170 , n2171 , n2172 ,
     n2173 , n2174 , n2175 , n2176 , n2177 , n2178 , n2179 , n2180 , n2181 , n2182 ,
     n2183 , n2184 , n2185 , n2186 , n2187 , n2188 , n2189 , n2190 , n2191 , n2192 ,
     n2193 , n2194 , n2195 , n2196 , n2197 , n2198 , n2199 , n2200 , n2201 , n2202 ,
     n2203 , n2204 , n2205 , n2206 , n2207 , n2208 , n2209 , n2210 , n2211 , n2212 ,
     n2213 , n2214 , n2215 , n2216 , n2217 , n2218 , n2219 , n2220 , n2221 , n2222 ,
     n2223 , n2224 , n2225 , n2226 , n2227 , n2228 , n2229 , n2230 , n2231 , n2232 ,
     n2233 , n2234 , n2235 , n2236 , n2237 , n2238 , n2239 , n2240 , n2241 , n2242 ,
     n2243 , n2244 , n2245 , n2246 , n2247 , n2248 , n2249 , n2250 , n2251 , n2252 ,
     n2253 , n2254 , n2255 , n2256 , n2257 , n2258 , n2259 , n2260 , n2261 , n2262 ,
     n2263 , n2264 , n2265 , n2266 , n2267 , n2268 , n2269 , n2270 , n2271 , n2272 ,
     n2273 , n2274 , n2275 , n2276 , n2277 , n2278 , n2279 , n2280 , n2281 , n2282 ,
     n2283 , n2284 , n2285 , n2286 , n2287 , n2288 , n2289 , n2290 , n2291 , n2292 ,
     n2293 , n2294 , n2295 , n2296 , n2297 , n2298 , n2299 , n2300 , n2301 , n2302 ,
     n2303 , n2304 , n2305 , n2306 , n2307 , n2308 , n2309 , n2310 , n2311 , n2312 ,
     n2313 , n2314 , n2315 , n2316 , n2317 , n2318 , n2319 , n2320 , n2321 , n2322 ,
     n2323 , n2324 , n2325 , n2326 , n2327 , n2328 , n2329 , n2330 , n2331 , n2332 ,
     n2333 , n2334 , n2335 , n2336 , n2337 , n2338 , n2339 , n2340 , n2341 , n2342 ,
     n2343 , n2344 , n2345 , n2346 , n2347 , n2348 , n2349 , n2350 , n2351 , n2352 ,
     n2353 , n2354 , n2355 , n2356 , n2357 , n2358 , n2359 , n2360 , n2361 , n2362 ,
     n2363 , n2364 , n2365 , n2366 , n2367 , n2368 , n2369 , n2370 , n2371 , n2372 ,
     n2373 , n2374 , n2375 , n2376 , n2377 , n2378 , n2379 , n2380 , n2381 , n2382 ,
     n2383 , n2384 , n2385 , n2386 , n2387 , n2388 , n2389 , n2390 , n2391 , n2392 ,
     n2393 , n2394 , n2395 , n2396 , n2397 , n2398 , n2399 , n2400 , n2401 , n2402 ,
     n2403 , n2404 , n2405 , n2406 , n2407 , n2408 , n2409 , n2410 , n2411 , n2412 ,
     n2413 , n2414 , n2415 , n2416 , n2417 , n2418 , n2419 , n2420 , n2421 , n2422 ,
     n2423 , n2424 , n2425 , n2426 , n2427 , n2428 , n2429 , n2430 , n2431 , n2432 ,
     n2433 , n2434 , n2435 , n2436 , n2437 , n2438 , n2439 , n2440 , n2441 , n2442 ,
     n2443 , n2444 , n2445 , n2446 , n2447 , n2448 , n2449 , n2450 , n2451 , n2452 ,
     n2453 , n2454 , n2455 , n2456 , n2457 , n2458 , n2459 , n2460 , n2461 , n2462 ,
     n2463 , n2464 , n2465 , n2466 , n2467 , n2468 , n2469 , n2470 , n2471 , n2472 ,
     n2473 , n2474 , n2475 , n2476 , n2477 , n2478 , n2479 , n2480 , n2481 , n2482 ,
     n2483 , n2484 , n2485 , n2486 , n2487 , n2488 , n2489 , n2490 , n2491 , n2492 ,
     n2493 , n2494 , n2495 , n2496 , n2497 , n2498 , n2499 , n2500 , n2501 , n2502 ,
     n2503 , n2504 , n2505 , n2506 , n2507 , n2508 , n2509 , n2510 , n2511 , n2512 ,
     n2513 , n2514 , n2515 , n2516 , n2517 , n2518 , n2519 , n2520 , n2521 , n2522 ,
     n2523 , n2524 , n2525 , n2526 , n2527 , n2528 , n2529 , n2530 , n2531 , n2532 ,
     n2533 , n2534 , n2535 , n2536 , n2537 , n2538 , n2539 , n2540 , n2541 , n2542 ,
     n2543 , n2544 , n2545 , n2546 , n2547 , n2548 , n2549 , n2550 , n2551 , n2552 ,
     n2553 , n2554 , n2555 , n2556 , n2557 , n2558 , n2559 , n2560 , n2561 , n2562 ,
     n2563 , n2564 , n2565 , n2566 , n2567 , n2568 , n2569 , n2570 , n2571 , n2572 ,
     n2573 , n2574 , n2575 , n2576 , n2577 , n2578 , n2579 , n2580 , n2581 , n2582 ,
     n2583 , n2584 , n2585 , n2586 , n2587 , n2588 , n2589 , n2590 , n2591 , n2592 ,
     n2593 , n2594 , n2595 , n2596 , n2597 , n2598 , n2599 , n2600 , n2601 , n2602 ,
     n2603 , n2604 , n2605 , n2606 , n2607 , n2608 , n2609 , n2610 , n2611 , n2612 ,
     n2613 , n2614 , n2615 , n2616 , n2617 , n2618 , n2619 , n2620 , n2621 , n2622 ,
     n2623 , n2624 , n2625 , n2626 , n2627 , n2628 , n2629 , n2630 , n2631 , n2632 ,
     n2633 , n2634 , n2635 , n2636 , n2637 , n2638 , n2639 , n2640 , n2641 , n2642 ,
     n2643 , n2644 , n2645 , n2646 , n2647 , n2648 , n2649 , n2650 , n2651 , n2652 ,
     n2653 , n2654 , n2655 , n2656 , n2657 , n2658 , n2659 , n2660 , n2661 , n2662 ,
     n2663 , n2664 , n2665 , n2666 , n2667 , n2668 , n2669 , n2670 , n2671 , n2672 ,
     n2673 , n2674 , n2675 , n2676 , n2677 , n2678 , n2679 , n2680 , n2681 , n2682 ,
     n2683 , n2684 , n2685 , n2686 , n2687 , n2688 , n2689 , n2690 , n2691 , n2692 ,
     n2693 , n2694 , n2695 , n2696 , n2697 , n2698 , n2699 , n2700 , n2701 , n2702 ,
     n2703 , n2704 , n2705 , n2706 , n2707 , n2708 , n2709 , n2710 , n2711 , n2712 ,
     n2713 , n2714 , n2715 , n2716 , n2717 , n2718 , n2719 , n2720 , n2721 , n2722 ,
     n2723 , n2724 , n2725 , n2726 , n2727 , n2728 , n2729 , n2730 , n2731 , n2732 ,
     n2733 , n2734 , n2735 , n2736 , n2737 , n2738 , n2739 , n2740 , n2741 , n2742 ,
     n2743 , n2744 , n2745 , n2746 , n2747 , n2748 , n2749 , n2750 , n2751 , n2752 ,
     n2753 , n2754 , n2755 , n2756 , n2757 , n2758 , n2759 , n2760 , n2761 , n2762 ,
     n2763 , n2764 , n2765 , n2766 , n2767 , n2768 , n2769 , n2770 , n2771 , n2772 ,
     n2773 , n2774 , n2775 , n2776 , n2777 , n2778 , n2779 , n2780 , n2781 , n2782 ,
     n2783 , n2784 , n2785 , n2786 , n2787 , n2788 , n2789 , n2790 , n2791 , n2792 ,
     n2793 , n2794 , n2795 , n2796 , n2797 , n2798 , n2799 , n2800 , n2801 , n2802 ,
     n2803 , n2804 , n2805 , n2806 , n2807 , n2808 , n2809 , n2810 , n2811 , n2812 ,
     n2813 , n2814 , n2815 , n2816 , n2817 , n2818 , n2819 , n2820 , n2821 , n2822 ,
     n2823 , n2824 , n2825 , n2826 , n2827 , n2828 , n2829 , n2830 , n2831 , n2832 ,
     n2833 , n2834 , n2835 , n2836 , n2837 , n2838 , n2839 , n2840 , n2841 , n2842 ,
     n2843 , n2844 , n2845 , n2846 , n2847 , n2848 , n2849 , n2850 , n2851 , n2852 ,
     n2853 , n2854 , n2855 , n2856 , n2857 , n2858 , n2859 , n2860 , n2861 , n2862 ,
     n2863 , n2864 , n2865 , n2866 , n2867 , n2868 , n2869 , n2870 , n2871 , n2872 ,
     n2873 , n2874 , n2875 , n2876 , n2877 , n2878 , n2879 , n2880 , n2881 , n2882 ,
     n2883 , n2884 , n2885 , n2886 , n2887 , n2888 , n2889 , n2890 , n2891 , n2892 ,
     n2893 , n2894 , n2895 , n2896 , n2897 , n2898 , n2899 , n2900 , n2901 , n2902 ,
     n2903 , n2904 , n2905 , n2906 , n2907 , n2908 , n2909 , n2910 , n2911 , n2912 ,
     n2913 , n2914 , n2915 , n2916 , n2917 , n2918 , n2919 , n2920 , n2921 , n2922 ,
     n2923 , n2924 , n2925 , n2926 , n2927 , n2928 , n2929 , n2930 , n2931 , n2932 ,
     n2933 , n2934 , n2935 , n2936 , n2937 , n2938 , n2939 , n2940 , n2941 , n2942 ,
     n2943 , n2944 , n2945 , n2946 , n2947 , n2948 , n2949 , n2950 , n2951 , n2952 ,
     n2953 , n2954 , n2955 , n2956 , n2957 , n2958 , n2959 , n2960 , n2961 , n2962 ,
     n2963 , n2964 , n2965 , n2966 , n2967 , n2968 , n2969 , n2970 , n2971 , n2972 ,
     n2973 , n2974 , n2975 , n2976 , n2977 , n2978 , n2979 , n2980 , n2981 , n2982 ,
     n2983 , n2984 , n2985 , n2986 , n2987 , n2988 , n2989 , n2990 , n2991 , n2992 ,
     n2993 , n2994 , n2995 , n2996 , n2997 , n2998 , n2999 , n3000 , n3001 , n3002 ,
     n3003 , n3004 , n3005 , n3006 , n3007 , n3008 , n3009 , n3010 , n3011 , n3012 ,
     n3013 , n3014 , n3015 , n3016 , n3017 , n3018 , n3019 , n3020 , n3021 , n3022 ,
     n3023 , n3024 , n3025 , n3026 , n3027 , n3028 , n3029 , n3030 , n3031 , n3032 ,
     n3033 , n3034 , n3035 , n3036 , n3037 , n3038 , n3039 , n3040 , n3041 , n3042 ,
     n3043 , n3044 , n3045 , n3046 , n3047 , n3048 , n3049 , n3050 , n3051 , n3052 ,
     n3053 , n3054 , n3055 , n3056 , n3057 , n3058 , n3059 , n3060 , n3061 , n3062 ,
     n3063 , n3064 , n3065 , n3066 , n3067 , n3068 , n3069 , n3070 , n3071 , n3072 ,
     n3073 , n3074 , n3075 , n3076 , n3077 , n3078 , n3079 , n3080 , n3081 , n3082 ,
     n3083 , n3084 , n3085 , n3086 , n3087 , n3088 , n3089 , n3090 , n3091 , n3092 ,
     n3093 , n3094 , n3095 , n3096 , n3097 , n3098 , n3099 , n3100 , n3101 , n3102 ,
     n3103 , n3104 , n3105 , n3106 , n3107 , n3108 , n3109 , n3110 , n3111 , n3112 ,
     n3113 , n3114 , n3115 , n3116 , n3117 , n3118 , n3119 , n3120 , n3121 , n3122 ,
     n3123 , n3124 , n3125 , n3126 , n3127 , n3128 , n3129 , n3130 , n3131 , n3132 ,
     n3133 , n3134 , n3135 , n3136 , n3137 , n3138 , n3139 , n3140 , n3141 , n3142 ,
     n3143 , n3144 , n3145 , n3146 , n3147 , n3148 , n3149 , n3150 , n3151 , n3152 ,
     n3153 , n3154 , n3155 , n3156 , n3157 , n3158 , n3159 , n3160 , n3161 , n3162 ,
     n3163 , n3164 , n3165 , n3166 , n3167 , n3168 , n3169 , n3170 , n3171 , n3172 ,
     n3173 , n3174 , n3175 , n3176 , n3177 , n3178 , n3179 , n3180 , n3181 , n3182 ,
     n3183 , n3184 , n3185 , n3186 , n3187 , n3188 , n3189 , n3190 , n3191 , n3192 ,
     n3193 , n3194 , n3195 , n3196 , n3197 , n3198 , n3199 , n3200 , n3201 , n3202 ,
     n3203 , n3204 , n3205 , n3206 , n3207 , n3208 , n3209 , n3210 , n3211 , n3212 ,
     n3213 , n3214 , n3215 , n3216 , n3217 , n3218 , n3219 , n3220 , n3221 , n3222 ,
     n3223 , n3224 , n3225 , n3226 , n3227 , n3228 , n3229 , n3230 , n3231 , n3232 ,
     n3233 , n3234 , n3235 , n3236 , n3237 , n3238 , n3239 , n3240 , n3241 , n3242 ,
     n3243 , n3244 , n3245 , n3246 , n3247 , n3248 , n3249 , n3250 , n3251 , n3252 ,
     n3253 , n3254 , n3255 , n3256 , n3257 , n3258 , n3259 , n3260 , n3261 , n3262 ,
     n3263 , n3264 , n3265 , n3266 , n3267 , n3268 , n3269 , n3270 , n3271 , n3272 ,
     n3273 , n3274 , n3275 , n3276 , n3277 , n3278 , n3279 , n3280 , n3281 , n3282 ,
     n3283 , n3284 , n3285 , n3286 , n3287 , n3288 , n3289 , n3290 , n3291 , n3292 ,
     n3293 , n3294 , n3295 , n3296 , n3297 , n3298 , n3299 , n3300 , n3301 , n3302 ,
     n3303 , n3304 , n3305 , n3306 , n3307 , n3308 , n3309 , n3310 , n3311 , n3312 ,
     n3313 , n3314 , n3315 , n3316 , n3317 , n3318 , n3319 , n3320 , n3321 , n3322 ,
     n3323 , n3324 , n3325 , n3326 , n3327 , n3328 , n3329 , n3330 , n3331 , n3332 ,
     n3333 , n3334 , n3335 , n3336 , n3337 , n3338 , n3339 , n3340 , n3341 , n3342 ,
     n3343 , n3344 , n3345 , n3346 , n3347 , n3348 , n3349 , n3350 , n3351 , n3352 ,
     n3353 , n3354 , n3355 , n3356 , n3357 , n3358 , n3359 , n3360 , n3361 , n3362 ,
     n3363 , n3364 , n3365 , n3366 , n3367 , n3368 , n3369 , n3370 , n3371 , n3372 ,
     n3373 , n3374 , n3375 , n3376 , n3377 , n3378 , n3379 , n3380 , n3381 , n3382 ,
     n3383 , n3384 , n3385 , n3386 , n3387 , n3388 , n3389 , n3390 , n3391 , n3392 ,
     n3393 , n3394 , n3395 , n3396 , n3397 , n3398 , n3399 , n3400 , n3401 , n3402 ,
     n3403 , n3404 , n3405 , n3406 , n3407 , n3408 , n3409 , n3410 , n3411 , n3412 ,
     n3413 , n3414 , n3415 , n3416 , n3417 , n3418 , n3419 , n3420 , n3421 , n3422 ,
     n3423 , n3424 , n3425 , n3426 , n3427 , n3428 , n3429 , n3430 , n3431 , n3432 ,
     n3433 , n3434 , n3435 , n3436 , n3437 , n3438 , n3439 , n3440 , n3441 , n3442 ,
     n3443 , n3444 , n3445 , n3446 , n3447 , n3448 , n3449 , n3450 , n3451 , n3452 ,
     n3453 , n3454 , n3455 , n3456 , n3457 , n3458 , n3459 , n3460 , n3461 , n3462 ,
     n3463 , n3464 , n3465 , n3466 , n3467 , n3468 , n3469 , n3470 , n3471 , n3472 ,
     n3473 , n3474 , n3475 , n3476 , n3477 , n3478 , n3479 , n3480 , n3481 , n3482 ,
     n3483 , n3484 , n3485 , n3486 , n3487 , n3488 , n3489 , n3490 , n3491 , n3492 ,
     n3493 , n3494 , n3495 , n3496 , n3497 , n3498 , n3499 , n3500 , n3501 , n3502 ,
     n3503 , n3504 , n3505 , n3506 , n3507 , n3508 , n3509 , n3510 , n3511 , n3512 ,
     n3513 , n3514 , n3515 , n3516 , n3517 , n3518 , n3519 , n3520 , n3521 , n3522 ,
     n3523 , n3524 , n3525 , n3526 , n3527 , n3528 , n3529 , n3530 , n3531 , n3532 ,
     n3533 , n3534 , n3535 , n3536 , n3537 , n3538 , n3539 , n3540 , n3541 , n3542 ,
     n3543 , n3544 , n3545 , n3546 , n3547 , n3548 , n3549 , n3550 , n3551 , n3552 ,
     n3553 , n3554 , n3555 , n3556 , n3557 , n3558 , n3559 , n3560 , n3561 , n3562 ,
     n3563 , n3564 , n3565 , n3566 , n3567 , n3568 , n3569 , n3570 , n3571 , n3572 ,
     n3573 , n3574 , n3575 , n3576 , n3577 , n3578 , n3579 , n3580 , n3581 , n3582 ,
     n3583 , n3584 , n3585 , n3586 , n3587 , n3588 , n3589 , n3590 , n3591 , n3592 ,
     n3593 , n3594 , n3595 , n3596 , n3597 , n3598 , n3599 , n3600 , n3601 , n3602 ,
     n3603 , n3604 , n3605 , n3606 , n3607 , n3608 , n3609 , n3610 , n3611 , n3612 ,
     n3613 , n3614 , n3615 , n3616 , n3617 , n3618 , n3619 , n3620 , n3621 , n3622 ,
     n3623 , n3624 , n3625 , n3626 , n3627 , n3628 , n3629 , n3630 , n3631 , n3632 ,
     n3633 , n3634 , n3635 , n3636 , n3637 , n3638 , n3639 , n3640 , n3641 , n3642 ,
     n3643 , n3644 , n3645 , n3646 , n3647 , n3648 , n3649 , n3650 , n3651 , n3652 ,
     n3653 , n3654 , n3655 , n3656 , n3657 , n3658 , n3659 , n3660 , n3661 , n3662 ,
     n3663 , n3664 , n3665 , n3666 , n3667 , n3668 , n3669 , n3670 , n3671 , n3672 ,
     n3673 , n3674 , n3675 , n3676 , n3677 , n3678 , n3679 , n3680 , n3681 , n3682 ,
     n3683 , n3684 , n3685 , n3686 , n3687 , n3688 , n3689 , n3690 , n3691 , n3692 ,
     n3693 , n3694 , n3695 , n3696 , n3697 , n3698 , n3699 , n3700 , n3701 , n3702 ,
     n3703 , n3704 , n3705 , n3706 , n3707 , n3708 , n3709 , n3710 , n3711 , n3712 ,
     n3713 , n3714 , n3715 , n3716 , n3717 , n3718 , n3719 , n3720 , n3721 , n3722 ,
     n3723 , n3724 , n3725 , n3726 , n3727 , n3728 , n3729 , n3730 , n3731 , n3732 ,
     n3733 , n3734 , n3735 , n3736 , n3737 , n3738 , n3739 , n3740 , n3741 , n3742 ,
     n3743 , n3744 , n3745 , n3746 , n3747 , n3748 , n3749 , n3750 , n3751 , n3752 ,
     n3753 , n3754 , n3755 , n3756 , n3757 , n3758 , n3759 , n3760 , n3761 , n3762 ,
     n3763 , n3764 , n3765 , n3766 , n3767 , n3768 , n3769 , n3770 , n3771 , n3772 ,
     n3773 , n3774 , n3775 , n3776 , n3777 , n3778 , n3779 , n3780 , n3781 , n3782 ,
     n3783 , n3784 , n3785 , n3786 , n3787 , n3788 , n3789 , n3790 , n3791 , n3792 ,
     n3793 , n3794 , n3795 , n3796 , n3797 , n3798 , n3799 , n3800 , n3801 , n3802 ,
     n3803 , n3804 , n3805 , n3806 , n3807 , n3808 , n3809 , n3810 , n3811 , n3812 ,
     n3813 , n3814 , n3815 , n3816 , n3817 , n3818 , n3819 , n3820 , n3821 , n3822 ,
     n3823 , n3824 , n3825 , n3826 , n3827 , n3828 , n3829 , n3830 , n3831 , n3832 ,
     n3833 , n3834 , n3835 , n3836 , n3837 , n3838 , n3839 , n3840 , n3841 , n3842 ,
     n3843 , n3844 , n3845 , n3846 , n3847 , n3848 , n3849 , n3850 , n3851 , n3852 ,
     n3853 , n3854 , n3855 , n3856 , n3857 , n3858 , n3859 , n3860 , n3861 , n3862 ,
     n3863 , n3864 , n3865 , n3866 , n3867 , n3868 , n3869 , n3870 , n3871 , n3872 ,
     n3873 , n3874 , n3875 , n3876 , n3877 , n3878 , n3879 , n3880 , n3881 , n3882 ,
     n3883 , n3884 , n3885 , n3886 , n3887 , n3888 , n3889 , n3890 , n3891 , n3892 ,
     n3893 , n3894 , n3895 , n3896 , n3897 , n3898 , n3899 , n3900 , n3901 , n3902 ,
     n3903 , n3904 , n3905 , n3906 , n3907 , n3908 , n3909 , n3910 , n3911 , n3912 ,
     n3913 , n3914 , n3915 , n3916 , n3917 , n3918 , n3919 , n3920 , n3921 , n3922 ,
     n3923 , n3924 , n3925 , n3926 , n3927 , n3928 , n3929 , n3930 , n3931 , n3932 ,
     n3933 , n3934 , n3935 , n3936 , n3937 , n3938 , n3939 , n3940 , n3941 , n3942 ,
     n3943 , n3944 , n3945 , n3946 , n3947 , n3948 , n3949 , n3950 , n3951 , n3952 ,
     n3953 , n3954 , n3955 , n3956 , n3957 , n3958 , n3959 , n3960 , n3961 , n3962 ,
     n3963 , n3964 , n3965 , n3966 , n3967 , n3968 , n3969 , n3970 , n3971 , n3972 ,
     n3973 , n3974 , n3975 , n3976 , n3977 , n3978 , n3979 , n3980 , n3981 , n3982 ,
     n3983 , n3984 , n3985 , n3986 , n3987 , n3988 , n3989 , n3990 , n3991 , n3992 ,
     n3993 , n3994 , n3995 , n3996 , n3997 , n3998 , n3999 , n4000 , n4001 , n4002 ,
     n4003 , n4004 , n4005 , n4006 , n4007 , n4008 , n4009 , n4010 , n4011 , n4012 ,
     n4013 , n4014 , n4015 , n4016 , n4017 , n4018 , n4019 , n4020 , n4021 , n4022 ,
     n4023 , n4024 , n4025 , n4026 , n4027 , n4028 , n4029 , n4030 , n4031 , n4032 ,
     n4033 , n4034 , n4035 , n4036 , n4037 , n4038 , n4039 , n4040 , n4041 , n4042 ,
     n4043 , n4044 , n4045 , n4046 , n4047 , n4048 , n4049 , n4050 , n4051 , n4052 ,
     n4053 , n4054 , n4055 , n4056 , n4057 , n4058 , n4059 , n4060 , n4061 , n4062 ,
     n4063 , n4064 , n4065 , n4066 , n4067 , n4068 , n4069 , n4070 , n4071 , n4072 ,
     n4073 , n4074 , n4075 , n4076 , n4077 , n4078 , n4079 , n4080 , n4081 , n4082 ,
     n4083 , n4084 , n4085 , n4086 , n4087 , n4088 , n4089 , n4090 , n4091 , n4092 ,
     n4093 , n4094 , n4095 , n4096 , n4097 , n4098 , n4099 , n4100 , n4101 , n4102 ,
     n4103 , n4104 , n4105 , n4106 , n4107 , n4108 , n4109 , n4110 , n4111 , n4112 ,
     n4113 , n4114 , n4115 , n4116 , n4117 , n4118 , n4119 , n4120 , n4121 , n4122 ,
     n4123 , n4124 , n4125 , n4126 , n4127 , n4128 , n4129 , n4130 , n4131 , n4132 ,
     n4133 , n4134 , n4135 , n4136 , n4137 , n4138 , n4139 , n4140 , n4141 , n4142 ,
     n4143 , n4144 , n4145 , n4146 , n4147 , n4148 , n4149 , n4150 , n4151 , n4152 ,
     n4153 , n4154 , n4155 , n4156 , n4157 , n4158 , n4159 , n4160 , n4161 , n4162 ,
     n4163 , n4164 , n4165 , n4166 , n4167 , n4168 , n4169 , n4170 , n4171 , n4172 ,
     n4173 , n4174 , n4175 , n4176 , n4177 , n4178 , n4179 , n4180 , n4181 , n4182 ,
     n4183 , n4184 , n4185 , n4186 , n4187 , n4188 , n4189 , n4190 , n4191 , n4192 ,
     n4193 , n4194 , n4195 , n4196 , n4197 , n4198 , n4199 , n4200 , n4201 , n4202 ,
     n4203 , n4204 , n4205 , n4206 , n4207 , n4208 , n4209 , n4210 , n4211 , n4212 ,
     n4213 , n4214 , n4215 , n4216 , n4217 , n4218 , n4219 , n4220 , n4221 , n4222 ,
     n4223 , n4224 , n4225 , n4226 , n4227 , n4228 , n4229 , n4230 , n4231 , n4232 ,
     n4233 , n4234 , n4235 , n4236 , n4237 , n4238 , n4239 , n4240 , n4241 , n4242 ,
     n4243 , n4244 , n4245 , n4246 , n4247 , n4248 , n4249 , n4250 , n4251 , n4252 ,
     n4253 , n4254 , n4255 , n4256 , n4257 , n4258 , n4259 , n4260 , n4261 , n4262 ,
     n4263 , n4264 , n4265 , n4266 , n4267 , n4268 , n4269 , n4270 , n4271 , n4272 ,
     n4273 , n4274 , n4275 , n4276 , n4277 , n4278 , n4279 , n4280 , n4281 , n4282 ,
     n4283 , n4284 , n4285 , n4286 , n4287 , n4288 , n4289 , n4290 , n4291 , n4292 ,
     n4293 , n4294 , n4295 , n4296 , n4297 , n4298 , n4299 , n4300 , n4301 , n4302 ,
     n4303 , n4304 , n4305 , n4306 , n4307 , n4308 , n4309 , n4310 , n4311 , n4312 ,
     n4313 , n4314 , n4315 , n4316 , n4317 , n4318 , n4319 , n4320 , n4321 , n4322 ,
     n4323 , n4324 , n4325 , n4326 , n4327 , n4328 , n4329 , n4330 , n4331 , n4332 ,
     n4333 , n4334 , n4335 , n4336 , n4337 , n4338 , n4339 , n4340 , n4341 , n4342 ,
     n4343 , n4344 , n4345 , n4346 , n4347 , n4348 , n4349 , n4350 , n4351 , n4352 ,
     n4353 , n4354 , n4355 , n4356 , n4357 , n4358 , n4359 , n4360 , n4361 , n4362 ,
     n4363 , n4364 , n4365 , n4366 , n4367 , n4368 , n4369 , n4370 , n4371 , n4372 ,
     n4373 , n4374 , n4375 , n4376 , n4377 , n4378 , n4379 , n4380 , n4381 , n4382 ,
     n4383 , n4384 , n4385 , n4386 , n4387 , n4388 , n4389 , n4390 , n4391 , n4392 ,
     n4393 , n4394 , n4395 , n4396 , n4397 , n4398 , n4399 , n4400 , n4401 , n4402 ,
     n4403 , n4404 , n4405 , n4406 , n4407 , n4408 , n4409 , n4410 , n4411 , n4412 ,
     n4413 , n4414 , n4415 , n4416 , n4417 , n4418 , n4419 , n4420 , n4421 , n4422 ,
     n4423 , n4424 , n4425 , n4426 , n4427 , n4428 , n4429 , n4430 , n4431 , n4432 ,
     n4433 , n4434 , n4435 , n4436 , n4437 , n4438 , n4439 , n4440 , n4441 , n4442 ,
     n4443 , n4444 , n4445 , n4446 , n4447 , n4448 , n4449 , n4450 , n4451 , n4452 ,
     n4453 , n4454 , n4455 , n4456 , n4457 , n4458 , n4459 , n4460 , n4461 , n4462 ,
     n4463 , n4464 , n4465 , n4466 , n4467 , n4468 , n4469 , n4470 , n4471 , n4472 ,
     n4473 , n4474 , n4475 , n4476 , n4477 , n4478 , n4479 , n4480 , n4481 , n4482 ,
     n4483 , n4484 , n4485 , n4486 , n4487 , n4488 , n4489 , n4490 , n4491 , n4492 ,
     n4493 , n4494 , n4495 , n4496 , n4497 , n4498 , n4499 , n4500 , n4501 , n4502 ,
     n4503 , n4504 , n4505 , n4506 , n4507 , n4508 , n4509 , n4510 , n4511 , n4512 ,
     n4513 , n4514 , n4515 , n4516 , n4517 , n4518 , n4519 , n4520 , n4521 , n4522 ,
     n4523 , n4524 , n4525 , n4526 , n4527 , n4528 , n4529 , n4530 , n4531 , n4532 ,
     n4533 , n4534 , n4535 , n4536 , n4537 , n4538 , n4539 , n4540 , n4541 , n4542 ,
     n4543 , n4544 , n4545 , n4546 , n4547 , n4548 , n4549 , n4550 , n4551 , n4552 ,
     n4553 , n4554 , n4555 , n4556 , n4557 , n4558 , n4559 , n4560 , n4561 , n4562 ,
     n4563 , n4564 , n4565 , n4566 , n4567 , n4568 , n4569 , n4570 , n4571 , n4572 ,
     n4573 , n4574 , n4575 , n4576 , n4577 , n4578 , n4579 , n4580 , n4581 , n4582 ,
     n4583 , n4584 , n4585 , n4586 , n4587 , n4588 , n4589 , n4590 , n4591 , n4592 ,
     n4593 , n4594 , n4595 , n4596 , n4597 , n4598 , n4599 , n4600 , n4601 , n4602 ,
     n4603 , n4604 , n4605 , n4606 , n4607 , n4608 , n4609 , n4610 , n4611 , n4612 ,
     n4613 , n4614 , n4615 , n4616 , n4617 , n4618 , n4619 , n4620 , n4621 , n4622 ,
     n4623 , n4624 , n4625 , n4626 , n4627 , n4628 , n4629 , n4630 , n4631 , n4632 ,
     n4633 , n4634 , n4635 , n4636 , n4637 , n4638 , n4639 , n4640 , n4641 , n4642 ,
     n4643 , n4644 , n4645 , n4646 , n4647 , n4648 , n4649 , n4650 , n4651 , n4652 ,
     n4653 , n4654 , n4655 , n4656 , n4657 , n4658 , n4659 , n4660 , n4661 , n4662 ,
     n4663 , n4664 , n4665 , n4666 , n4667 , n4668 , n4669 , n4670 , n4671 , n4672 ,
     n4673 , n4674 , n4675 , n4676 , n4677 , n4678 , n4679 , n4680 , n4681 , n4682 ,
     n4683 , n4684 , n4685 , n4686 , n4687 , n4688 , n4689 , n4690 , n4691 , n4692 ,
     n4693 , n4694 , n4695 , n4696 , n4697 , n4698 , n4699 , n4700 , n4701 , n4702 ,
     n4703 , n4704 , n4705 , n4706 , n4707 , n4708 , n4709 , n4710 , n4711 , n4712 ,
     n4713 , n4714 , n4715 , n4716 , n4717 , n4718 , n4719 , n4720 , n4721 , n4722 ,
     n4723 , n4724 , n4725 , n4726 , n4727 , n4728 , n4729 , n4730 , n4731 , n4732 ,
     n4733 , n4734 , n4735 , n4736 , n4737 , n4738 , n4739 , n4740 , n4741 , n4742 ,
     n4743 , n4744 , n4745 , n4746 , n4747 , n4748 , n4749 , n4750 , n4751 , n4752 ,
     n4753 , n4754 , n4755 , n4756 , n4757 , n4758 , n4759 , n4760 , n4761 , n4762 ,
     n4763 , n4764 , n4765 , n4766 , n4767 , n4768 , n4769 , n4770 , n4771 , n4772 ,
     n4773 , n4774 , n4775 , n4776 , n4777 , n4778 , n4779 , n4780 , n4781 , n4782 ,
     n4783 , n4784 , n4785 , n4786 , n4787 , n4788 , n4789 , n4790 , n4791 , n4792 ,
     n4793 , n4794 , n4795 , n4796 , n4797 , n4798 , n4799 , n4800 , n4801 , n4802 ,
     n4803 , n4804 , n4805 , n4806 , n4807 , n4808 , n4809 , n4810 , n4811 , n4812 ,
     n4813 , n4814 , n4815 , n4816 , n4817 , n4818 , n4819 , n4820 , n4821 , n4822 ,
     n4823 , n4824 , n4825 , n4826 , n4827 , n4828 , n4829 , n4830 , n4831 , n4832 ,
     n4833 , n4834 , n4835 , n4836 , n4837 , n4838 , n4839 , n4840 , n4841 , n4842 ,
     n4843 , n4844 , n4845 , n4846 , n4847 , n4848 , n4849 , n4850 , n4851 , n4852 ,
     n4853 , n4854 , n4855 , n4856 , n4857 , n4858 , n4859 , n4860 , n4861 , n4862 ,
     n4863 , n4864 , n4865 , n4866 , n4867 , n4868 , n4869 , n4870 , n4871 , n4872 ,
     n4873 , n4874 , n4875 , n4876 , n4877 , n4878 , n4879 , n4880 , n4881 , n4882 ,
     n4883 , n4884 , n4885 , n4886 , n4887 , n4888 , n4889 , n4890 , n4891 , n4892 ,
     n4893 , n4894 , n4895 , n4896 , n4897 , n4898 , n4899 , n4900 , n4901 , n4902 ,
     n4903 , n4904 , n4905 , n4906 , n4907 , n4908 , n4909 , n4910 , n4911 , n4912 ,
     n4913 , n4914 , n4915 , n4916 , n4917 , n4918 , n4919 , n4920 , n4921 , n4922 ,
     n4923 , n4924 , n4925 , n4926 , n4927 , n4928 , n4929 , n4930 , n4931 , n4932 ,
     n4933 , n4934 , n4935 , n4936 , n4937 , n4938 , n4939 , n4940 , n4941 , n4942 ,
     n4943 , n4944 , n4945 , n4946 , n4947 , n4948 , n4949 , n4950 , n4951 , n4952 ,
     n4953 , n4954 , n4955 , n4956 , n4957 , n4958 , n4959 , n4960 , n4961 , n4962 ,
     n4963 , n4964 , n4965 , n4966 , n4967 , n4968 , n4969 , n4970 , n4971 , n4972 ,
     n4973 , n4974 , n4975 , n4976 , n4977 , n4978 , n4979 , n4980 , n4981 , n4982 ,
     n4983 , n4984 , n4985 , n4986 , n4987 , n4988 , n4989 , n4990 , n4991 , n4992 ,
     n4993 , n4994 , n4995 , n4996 , n4997 , n4998 , n4999 , n5000 , n5001 , n5002 ,
     n5003 , n5004 , n5005 , n5006 , n5007 , n5008 , n5009 , n5010 , n5011 , n5012 ,
     n5013 , n5014 , n5015 , n5016 , n5017 , n5018 , n5019 , n5020 , n5021 , n5022 ,
     n5023 , n5024 , n5025 , n5026 , n5027 , n5028 , n5029 , n5030 , n5031 , n5032 ,
     n5033 , n5034 , n5035 , n5036 , n5037 , n5038 , n5039 , n5040 , n5041 , n5042 ,
     n5043 , n5044 , n5045 , n5046 , n5047 , n5048 , n5049 , n5050 , n5051 , n5052 ,
     n5053 , n5054 , n5055 , n5056 , n5057 , n5058 , n5059 , n5060 , n5061 , n5062 ,
     n5063 , n5064 , n5065 , n5066 , n5067 , n5068 , n5069 , n5070 , n5071 , n5072 ,
     n5073 , n5074 , n5075 , n5076 , n5077 , n5078 , n5079 , n5080 , n5081 , n5082 ,
     n5083 , n5084 , n5085 , n5086 , n5087 , n5088 , n5089 , n5090 , n5091 , n5092 ,
     n5093 , n5094 , n5095 , n5096 , n5097 , n5098 , n5099 , n5100 , n5101 , n5102 ,
     n5103 , n5104 , n5105 , n5106 , n5107 , n5108 , n5109 , n5110 , n5111 , n5112 ,
     n5113 , n5114 , n5115 , n5116 , n5117 , n5118 , n5119 , n5120 , n5121 , n5122 ,
     n5123 , n5124 , n5125 , n5126 , n5127 , n5128 , n5129 , n5130 , n5131 , n5132 ,
     n5133 , n5134 , n5135 , n5136 , n5137 , n5138 , n5139 , n5140 , n5141 , n5142 ,
     n5143 , n5144 , n5145 , n5146 , n5147 , n5148 , n5149 , n5150 , n5151 , n5152 ,
     n5153 , n5154 , n5155 , n5156 , n5157 , n5158 , n5159 , n5160 , n5161 , n5162 ,
     n5163 , n5164 , n5165 , n5166 , n5167 , n5168 , n5169 , n5170 , n5171 , n5172 ,
     n5173 , n5174 , n5175 , n5176 , n5177 , n5178 , n5179 , n5180 , n5181 , n5182 ,
     n5183 , n5184 , n5185 , n5186 , n5187 , n5188 , n5189 , n5190 , n5191 , n5192 ,
     n5193 , n5194 , n5195 , n5196 , n5197 , n5198 , n5199 , n5200 , n5201 , n5202 ,
     n5203 , n5204 , n5205 , n5206 , n5207 , n5208 , n5209 , n5210 , n5211 , n5212 ,
     n5213 , n5214 , n5215 , n5216 , n5217 , n5218 , n5219 , n5220 , n5221 , n5222 ,
     n5223 , n5224 , n5225 , n5226 , n5227 , n5228 , n5229 , n5230 , n5231 , n5232 ,
     n5233 , n5234 , n5235 , n5236 , n5237 , n5238 , n5239 , n5240 , n5241 , n5242 ,
     n5243 , n5244 , n5245 , n5246 , n5247 , n5248 , n5249 , n5250 , n5251 , n5252 ,
     n5253 , n5254 , n5255 , n5256 , n5257 , n5258 , n5259 , n5260 , n5261 , n5262 ,
     n5263 , n5264 , n5265 , n5266 , n5267 , n5268 , n5269 , n5270 , n5271 , n5272 ,
     n5273 , n5274 , n5275 , n5276 , n5277 , n5278 , n5279 , n5280 , n5281 , n5282 ,
     n5283 , n5284 , n5285 , n5286 , n5287 , n5288 , n5289 , n5290 , n5291 , n5292 ,
     n5293 , n5294 , n5295 , n5296 , n5297 , n5298 , n5299 , n5300 , n5301 , n5302 ,
     n5303 , n5304 , n5305 , n5306 , n5307 , n5308 , n5309 , n5310 , n5311 , n5312 ,
     n5313 , n5314 , n5315 , n5316 , n5317 , n5318 , n5319 , n5320 , n5321 , n5322 ,
     n5323 , n5324 , n5325 , n5326 , n5327 , n5328 , n5329 , n5330 , n5331 , n5332 ,
     n5333 , n5334 , n5335 , n5336 , n5337 , n5338 , n5339 , n5340 , n5341 , n5342 ,
     n5343 , n5344 , n5345 , n5346 , n5347 , n5348 , n5349 , n5350 , n5351 , n5352 ,
     n5353 , n5354 , n5355 , n5356 , n5357 , n5358 , n5359 , n5360 , n5361 , n5362 ,
     n5363 , n5364 , n5365 , n5366 , n5367 , n5368 , n5369 , n5370 , n5371 , n5372 ,
     n5373 , n5374 , n5375 , n5376 , n5377 , n5378 , n5379 , n5380 , n5381 , n5382 ,
     n5383 , n5384 , n5385 , n5386 , n5387 , n5388 , n5389 , n5390 , n5391 , n5392 ,
     n5393 , n5394 , n5395 , n5396 , n5397 , n5398 , n5399 , n5400 , n5401 , n5402 ,
     n5403 , n5404 , n5405 , n5406 , n5407 , n5408 , n5409 , n5410 , n5411 , n5412 ,
     n5413 , n5414 , n5415 , n5416 , n5417 , n5418 , n5419 , n5420 , n5421 , n5422 ,
     n5423 , n5424 , n5425 , n5426 , n5427 , n5428 , n5429 , n5430 , n5431 , n5432 ,
     n5433 , n5434 , n5435 , n5436 , n5437 , n5438 , n5439 , n5440 , n5441 , n5442 ,
     n5443 , n5444 , n5445 , n5446 , n5447 , n5448 , n5449 , n5450 , n5451 , n5452 ,
     n5453 , n5454 , n5455 , n5456 , n5457 , n5458 , n5459 , n5460 , n5461 , n5462 ,
     n5463 , n5464 , n5465 , n5466 , n5467 , n5468 , n5469 , n5470 , n5471 , n5472 ,
     n5473 , n5474 , n5475 , n5476 , n5477 , n5478 , n5479 , n5480 , n5481 , n5482 ,
     n5483 , n5484 , n5485 , n5486 , n5487 , n5488 , n5489 , n5490 , n5491 , n5492 ,
     n5493 , n5494 , n5495 , n5496 , n5497 , n5498 , n5499 , n5500 , n5501 , n5502 ,
     n5503 , n5504 , n5505 , n5506 , n5507 , n5508 , n5509 , n5510 , n5511 , n5512 ,
     n5513 , n5514 , n5515 , n5516 , n5517 , n5518 , n5519 , n5520 , n5521 , n5522 ,
     n5523 , n5524 , n5525 , n5526 , n5527 , n5528 , n5529 , n5530 , n5531 , n5532 ,
     n5533 , n5534 , n5535 , n5536 , n5537 , n5538 , n5539 , n5540 , n5541 , n5542 ,
     n5543 , n5544 , n5545 , n5546 , n5547 , n5548 , n5549 , n5550 , n5551 , n5552 ,
     n5553 , n5554 , n5555 , n5556 , n5557 , n5558 , n5559 , n5560 , n5561 , n5562 ,
     n5563 , n5564 , n5565 , n5566 , n5567 , n5568 , n5569 , n5570 , n5571 , n5572 ,
     n5573 , n5574 , n5575 , n5576 , n5577 , n5578 , n5579 , n5580 , n5581 , n5582 ,
     n5583 , n5584 , n5585 , n5586 , n5587 , n5588 , n5589 , n5590 , n5591 , n5592 ,
     n5593 , n5594 , n5595 , n5596 , n5597 , n5598 , n5599 , n5600 , n5601 , n5602 ,
     n5603 , n5604 , n5605 , n5606 , n5607 , n5608 , n5609 , n5610 , n5611 , n5612 ,
     n5613 , n5614 , n5615 , n5616 , n5617 , n5618 , n5619 , n5620 , n5621 , n5622 ,
     n5623 , n5624 , n5625 , n5626 , n5627 , n5628 , n5629 , n5630 , n5631 , n5632 ,
     n5633 , n5634 , n5635 , n5636 , n5637 , n5638 , n5639 , n5640 , n5641 , n5642 ,
     n5643 , n5644 , n5645 , n5646 , n5647 , n5648 , n5649 , n5650 , n5651 , n5652 ,
     n5653 , n5654 , n5655 , n5656 , n5657 , n5658 , n5659 , n5660 , n5661 , n5662 ,
     n5663 , n5664 , n5665 , n5666 , n5667 , n5668 , n5669 , n5670 , n5671 , n5672 ,
     n5673 , n5674 , n5675 , n5676 , n5677 , n5678 , n5679 , n5680 , n5681 , n5682 ,
     n5683 , n5684 , n5685 , n5686 , n5687 , n5688 , n5689 , n5690 , n5691 , n5692 ,
     n5693 , n5694 , n5695 , n5696 , n5697 , n5698 , n5699 , n5700 , n5701 , n5702 ,
     n5703 , n5704 , n5705 , n5706 , n5707 , n5708 , n5709 , n5710 , n5711 , n5712 ,
     n5713 , n5714 , n5715 , n5716 , n5717 , n5718 , n5719 , n5720 , n5721 , n5722 ,
     n5723 , n5724 , n5725 , n5726 , n5727 , n5728 , n5729 , n5730 , n5731 , n5732 ,
     n5733 , n5734 , n5735 , n5736 , n5737 , n5738 , n5739 , n5740 , n5741 , n5742 ,
     n5743 , n5744 , n5745 , n5746 , n5747 , n5748 , n5749 , n5750 , n5751 , n5752 ,
     n5753 , n5754 , n5755 , n5756 , n5757 , n5758 , n5759 , n5760 , n5761 , n5762 ,
     n5763 , n5764 , n5765 , n5766 , n5767 , n5768 , n5769 , n5770 , n5771 , n5772 ,
     n5773 , n5774 , n5775 , n5776 , n5777 , n5778 , n5779 , n5780 , n5781 , n5782 ,
     n5783 , n5784 , n5785 , n5786 , n5787 , n5788 , n5789 , n5790 , n5791 , n5792 ,
     n5793 , n5794 , n5795 , n5796 , n5797 , n5798 , n5799 , n5800 , n5801 , n5802 ,
     n5803 , n5804 , n5805 , n5806 , n5807 , n5808 , n5809 , n5810 , n5811 , n5812 ,
     n5813 , n5814 , n5815 , n5816 , n5817 , n5818 , n5819 , n5820 , n5821 , n5822 ,
     n5823 , n5824 , n5825 , n5826 , n5827 , n5828 , n5829 , n5830 , n5831 , n5832 ,
     n5833 , n5834 , n5835 , n5836 , n5837 , n5838 , n5839 , n5840 , n5841 , n5842 ,
     n5843 , n5844 , n5845 , n5846 , n5847 , n5848 , n5849 , n5850 , n5851 , n5852 ,
     n5853 , n5854 , n5855 , n5856 , n5857 , n5858 , n5859 , n5860 , n5861 , n5862 ,
     n5863 , n5864 , n5865 , n5866 , n5867 , n5868 , n5869 , n5870 , n5871 , n5872 ,
     n5873 , n5874 , n5875 , n5876 , n5877 , n5878 , n5879 , n5880 , n5881 , n5882 ,
     n5883 , n5884 , n5885 , n5886 , n5887 , n5888 , n5889 , n5890 , n5891 , n5892 ,
     n5893 , n5894 , n5895 , n5896 , n5897 , n5898 , n5899 , n5900 , n5901 , n5902 ,
     n5903 , n5904 , n5905 , n5906 , n5907 , n5908 , n5909 , n5910 , n5911 , n5912 ,
     n5913 , n5914 , n5915 , n5916 , n5917 , n5918 , n5919 , n5920 , n5921 , n5922 ,
     n5923 , n5924 , n5925 , n5926 , n5927 , n5928 , n5929 , n5930 , n5931 , n5932 ,
     n5933 , n5934 , n5935 , n5936 , n5937 , n5938 , n5939 , n5940 , n5941 , n5942 ,
     n5943 , n5944 , n5945 , n5946 , n5947 , n5948 , n5949 , n5950 , n5951 , n5952 ,
     n5953 , n5954 , n5955 , n5956 , n5957 , n5958 , n5959 , n5960 , n5961 , n5962 ,
     n5963 , n5964 , n5965 , n5966 , n5967 , n5968 , n5969 , n5970 , n5971 , n5972 ,
     n5973 , n5974 , n5975 , n5976 , n5977 , n5978 , n5979 , n5980 , n5981 , n5982 ,
     n5983 , n5984 , n5985 , n5986 , n5987 , n5988 , n5989 , n5990 , n5991 , n5992 ,
     n5993 , n5994 , n5995 , n5996 , n5997 , n5998 , n5999 , n6000 , n6001 , n6002 ,
     n6003 , n6004 , n6005 , n6006 , n6007 , n6008 , n6009 , n6010 , n6011 , n6012 ,
     n6013 , n6014 , n6015 , n6016 , n6017 , n6018 , n6019 , n6020 , n6021 , n6022 ,
     n6023 , n6024 , n6025 , n6026 , n6027 , n6028 , n6029 , n6030 , n6031 , n6032 ,
     n6033 , n6034 , n6035 , n6036 , n6037 , n6038 , n6039 , n6040 , n6041 , n6042 ,
     n6043 , n6044 , n6045 , n6046 , n6047 , n6048 , n6049 , n6050 , n6051 , n6052 ,
     n6053 , n6054 , n6055 , n6056 , n6057 , n6058 , n6059 , n6060 , n6061 , n6062 ,
     n6063 , n6064 , n6065 , n6066 , n6067 , n6068 , n6069 , n6070 , n6071 , n6072 ,
     n6073 , n6074 , n6075 , n6076 , n6077 , n6078 , n6079 , n6080 , n6081 , n6082 ,
     n6083 , n6084 , n6085 , n6086 , n6087 , n6088 , n6089 , n6090 , n6091 , n6092 ,
     n6093 , n6094 , n6095 , n6096 , n6097 , n6098 , n6099 , n6100 , n6101 , n6102 ,
     n6103 , n6104 , n6105 , n6106 , n6107 , n6108 , n6109 , n6110 , n6111 , n6112 ,
     n6113 , n6114 , n6115 , n6116 , n6117 , n6118 , n6119 , n6120 , n6121 , n6122 ,
     n6123 , n6124 , n6125 , n6126 , n6127 , n6128 , n6129 , n6130 , n6131 , n6132 ,
     n6133 , n6134 , n6135 , n6136 , n6137 , n6138 , n6139 , n6140 , n6141 , n6142 ,
     n6143 , n6144 , n6145 , n6146 , n6147 , n6148 , n6149 , n6150 , n6151 , n6152 ,
     n6153 , n6154 , n6155 , n6156 , n6157 , n6158 , n6159 , n6160 , n6161 , n6162 ,
     n6163 , n6164 , n6165 , n6166 , n6167 , n6168 , n6169 , n6170 , n6171 , n6172 ,
     n6173 , n6174 , n6175 , n6176 , n6177 , n6178 , n6179 , n6180 , n6181 , n6182 ,
     n6183 , n6184 , n6185 , n6186 , n6187 , n6188 , n6189 , n6190 , n6191 , n6192 ,
     n6193 , n6194 , n6195 , n6196 , n6197 , n6198 , n6199 , n6200 , n6201 , n6202 ,
     n6203 , n6204 , n6205 , n6206 , n6207 , n6208 , n6209 , n6210 , n6211 , n6212 ,
     n6213 , n6214 , n6215 , n6216 , n6217 , n6218 , n6219 , n6220 , n6221 , n6222 ,
     n6223 , n6224 , n6225 , n6226 , n6227 , n6228 , n6229 , n6230 , n6231 , n6232 ,
     n6233 , n6234 , n6235 , n6236 , n6237 , n6238 , n6239 , n6240 , n6241 , n6242 ,
     n6243 , n6244 , n6245 , n6246 , n6247 , n6248 , n6249 , n6250 , n6251 , n6252 ,
     n6253 , n6254 , n6255 , n6256 , n6257 , n6258 , n6259 , n6260 , n6261 , n6262 ,
     n6263 , n6264 , n6265 , n6266 , n6267 , n6268 , n6269 , n6270 , n6271 , n6272 ,
     n6273 , n6274 , n6275 , n6276 , n6277 , n6278 , n6279 , n6280 , n6281 , n6282 ,
     n6283 , n6284 , n6285 , n6286 , n6287 , n6288 , n6289 , n6290 , n6291 , n6292 ,
     n6293 , n6294 , n6295 , n6296 , n6297 , n6298 , n6299 , n6300 , n6301 , n6302 ,
     n6303 , n6304 , n6305 , n6306 , n6307 , n6308 , n6309 , n6310 , n6311 , n6312 ,
     n6313 , n6314 , n6315 , n6316 , n6317 , n6318 , n6319 , n6320 , n6321 , n6322 ,
     n6323 , n6324 , n6325 , n6326 , n6327 , n6328 , n6329 , n6330 , n6331 , n6332 ,
     n6333 , n6334 , n6335 , n6336 , n6337 , n6338 , n6339 , n6340 , n6341 , n6342 ,
     n6343 , n6344 , n6345 , n6346 , n6347 , n6348 , n6349 , n6350 , n6351 , n6352 ,
     n6353 , n6354 , n6355 , n6356 , n6357 , n6358 , n6359 , n6360 , n6361 , n6362 ,
     n6363 , n6364 , n6365 , n6366 , n6367 , n6368 , n6369 , n6370 , n6371 , n6372 ,
     n6373 , n6374 , n6375 , n6376 , n6377 , n6378 , n6379 , n6380 , n6381 , n6382 ,
     n6383 , n6384 , n6385 , n6386 , n6387 , n6388 , n6389 , n6390 , n6391 , n6392 ,
     n6393 , n6394 , n6395 , n6396 , n6397 , n6398 , n6399 , n6400 , n6401 , n6402 ,
     n6403 , n6404 , n6405 , n6406 , n6407 , n6408 , n6409 , n6410 , n6411 , n6412 ,
     n6413 , n6414 , n6415 , n6416 , n6417 , n6418 , n6419 , n6420 , n6421 , n6422 ,
     n6423 , n6424 , n6425 , n6426 , n6427 , n6428 , n6429 , n6430 , n6431 , n6432 ,
     n6433 , n6434 , n6435 , n6436 , n6437 , n6438 , n6439 , n6440 , n6441 , n6442 ,
     n6443 , n6444 , n6445 , n6446 , n6447 , n6448 , n6449 , n6450 , n6451 , n6452 ,
     n6453 , n6454 , n6455 , n6456 , n6457 , n6458 , n6459 , n6460 , n6461 , n6462 ,
     n6463 , n6464 , n6465 , n6466 , n6467 , n6468 , n6469 , n6470 , n6471 , n6472 ,
     n6473 , n6474 , n6475 , n6476 , n6477 , n6478 , n6479 , n6480 , n6481 , n6482 ,
     n6483 , n6484 , n6485 , n6486 , n6487 , n6488 , n6489 , n6490 , n6491 , n6492 ,
     n6493 , n6494 , n6495 , n6496 , n6497 , n6498 , n6499 , n6500 , n6501 , n6502 ,
     n6503 , n6504 , n6505 , n6506 , n6507 , n6508 , n6509 , n6510 , n6511 , n6512 ,
     n6513 , n6514 , n6515 , n6516 , n6517 , n6518 , n6519 , n6520 , n6521 , n6522 ,
     n6523 , n6524 , n6525 , n6526 , n6527 , n6528 , n6529 , n6530 , n6531 , n6532 ,
     n6533 , n6534 , n6535 , n6536 , n6537 , n6538 , n6539 , n6540 , n6541 , n6542 ,
     n6543 , n6544 , n6545 , n6546 , n6547 , n6548 , n6549 , n6550 , n6551 , n6552 ,
     n6553 , n6554 , n6555 , n6556 , n6557 , n6558 , n6559 , n6560 , n6561 , n6562 ,
     n6563 , n6564 , n6565 , n6566 , n6567 , n6568 , n6569 , n6570 , n6571 , n6572 ,
     n6573 , n6574 , n6575 , n6576 , n6577 , n6578 , n6579 , n6580 , n6581 , n6582 ,
     n6583 , n6584 , n6585 , n6586 , n6587 , n6588 , n6589 , n6590 , n6591 , n6592 ,
     n6593 , n6594 , n6595 , n6596 , n6597 , n6598 , n6599 , n6600 , n6601 , n6602 ,
     n6603 , n6604 , n6605 , n6606 , n6607 , n6608 , n6609 , n6610 , n6611 , n6612 ,
     n6613 , n6614 , n6615 , n6616 , n6617 , n6618 , n6619 , n6620 , n6621 , n6622 ,
     n6623 , n6624 , n6625 , n6626 , n6627 , n6628 , n6629 , n6630 , n6631 , n6632 ,
     n6633 , n6634 , n6635 , n6636 , n6637 , n6638 , n6639 , n6640 , n6641 , n6642 ,
     n6643 , n6644 , n6645 , n6646 , n6647 , n6648 , n6649 , n6650 , n6651 , n6652 ,
     n6653 , n6654 , n6655 , n6656 , n6657 , n6658 , n6659 , n6660 , n6661 , n6662 ,
     n6663 , n6664 , n6665 , n6666 , n6667 , n6668 , n6669 , n6670 , n6671 , n6672 ,
     n6673 , n6674 , n6675 , n6676 , n6677 , n6678 , n6679 , n6680 , n6681 , n6682 ,
     n6683 , n6684 , n6685 , n6686 , n6687 , n6688 , n6689 , n6690 , n6691 , n6692 ,
     n6693 , n6694 , n6695 , n6696 , n6697 , n6698 , n6699 , n6700 , n6701 , n6702 ,
     n6703 , n6704 , n6705 , n6706 , n6707 , n6708 , n6709 , n6710 , n6711 , n6712 ,
     n6713 , n6714 , n6715 , n6716 , n6717 , n6718 , n6719 , n6720 , n6721 , n6722 ,
     n6723 , n6724 , n6725 , n6726 , n6727 , n6728 , n6729 , n6730 , n6731 , n6732 ,
     n6733 , n6734 , n6735 , n6736 , n6737 , n6738 , n6739 , n6740 , n6741 , n6742 ,
     n6743 , n6744 , n6745 , n6746 , n6747 , n6748 , n6749 , n6750 , n6751 , n6752 ,
     n6753 , n6754 , n6755 , n6756 , n6757 , n6758 , n6759 , n6760 , n6761 , n6762 ,
     n6763 , n6764 , n6765 , n6766 , n6767 , n6768 , n6769 , n6770 , n6771 , n6772 ,
     n6773 , n6774 , n6775 , n6776 , n6777 , n6778 , n6779 , n6780 , n6781 , n6782 ,
     n6783 , n6784 , n6785 , n6786 , n6787 , n6788 , n6789 , n6790 , n6791 , n6792 ,
     n6793 , n6794 , n6795 , n6796 , n6797 , n6798 , n6799 , n6800 , n6801 , n6802 ,
     n6803 , n6804 , n6805 , n6806 , n6807 , n6808 , n6809 , n6810 , n6811 , n6812 ,
     n6813 , n6814 , n6815 , n6816 , n6817 , n6818 , n6819 , n6820 , n6821 , n6822 ,
     n6823 , n6824 , n6825 , n6826 , n6827 , n6828 , n6829 , n6830 , n6831 , n6832 ,
     n6833 , n6834 , n6835 , n6836 , n6837 , n6838 , n6839 , n6840 , n6841 , n6842 ,
     n6843 , n6844 , n6845 , n6846 , n6847 , n6848 , n6849 , n6850 , n6851 , n6852 ,
     n6853 , n6854 , n6855 , n6856 , n6857 , n6858 , n6859 , n6860 , n6861 , n6862 ,
     n6863 , n6864 , n6865 , n6866 , n6867 , n6868 , n6869 , n6870 , n6871 , n6872 ,
     n6873 , n6874 , n6875 , n6876 , n6877 , n6878 , n6879 , n6880 , n6881 , n6882 ,
     n6883 , n6884 , n6885 , n6886 , n6887 , n6888 , n6889 , n6890 , n6891 , n6892 ,
     n6893 , n6894 , n6895 , n6896 , n6897 , n6898 , n6899 , n6900 , n6901 , n6902 ,
     n6903 , n6904 , n6905 , n6906 , n6907 , n6908 , n6909 , n6910 , n6911 , n6912 ,
     n6913 , n6914 , n6915 , n6916 , n6917 , n6918 , n6919 , n6920 , n6921 , n6922 ,
     n6923 , n6924 , n6925 , n6926 , n6927 , n6928 , n6929 , n6930 , n6931 , n6932 ,
     n6933 , n6934 , n6935 , n6936 , n6937 , n6938 , n6939 , n6940 , n6941 , n6942 ,
     n6943 , n6944 , n6945 , n6946 , n6947 , n6948 , n6949 , n6950 , n6951 , n6952 ,
     n6953 , n6954 , n6955 , n6956 , n6957 , n6958 , n6959 , n6960 , n6961 , n6962 ,
     n6963 , n6964 , n6965 , n6966 , n6967 , n6968 , n6969 , n6970 , n6971 , n6972 ,
     n6973 , n6974 , n6975 , n6976 , n6977 , n6978 , n6979 , n6980 , n6981 , n6982 ,
     n6983 , n6984 , n6985 , n6986 , n6987 , n6988 , n6989 , n6990 , n6991 , n6992 ,
     n6993 , n6994 , n6995 , n6996 , n6997 , n6998 , n6999 , n7000 , n7001 , n7002 ,
     n7003 , n7004 , n7005 , n7006 , n7007 , n7008 , n7009 , n7010 , n7011 , n7012 ,
     n7013 , n7014 , n7015 , n7016 , n7017 , n7018 , n7019 , n7020 , n7021 , n7022 ,
     n7023 , n7024 , n7025 , n7026 , n7027 , n7028 , n7029 , n7030 , n7031 , n7032 ,
     n7033 , n7034 , n7035 , n7036 , n7037 , n7038 , n7039 , n7040 , n7041 , n7042 ,
     n7043 , n7044 , n7045 , n7046 , n7047 , n7048 , n7049 , n7050 , n7051 , n7052 ,
     n7053 , n7054 , n7055 , n7056 , n7057 , n7058 , n7059 , n7060 , n7061 , n7062 ,
     n7063 , n7064 , n7065 , n7066 , n7067 , n7068 , n7069 , n7070 , n7071 , n7072 ,
     n7073 , n7074 , n7075 , n7076 , n7077 , n7078 , n7079 , n7080 , n7081 , n7082 ,
     n7083 , n7084 , n7085 , n7086 , n7087 , n7088 , n7089 , n7090 , n7091 , n7092 ,
     n7093 , n7094 , n7095 , n7096 , n7097 , n7098 , n7099 , n7100 , n7101 , n7102 ,
     n7103 , n7104 , n7105 , n7106 , n7107 , n7108 , n7109 , n7110 , n7111 , n7112 ,
     n7113 , n7114 , n7115 , n7116 , n7117 , n7118 , n7119 , n7120 , n7121 , n7122 ,
     n7123 , n7124 , n7125 , n7126 , n7127 , n7128 , n7129 , n7130 , n7131 , n7132 ,
     n7133 , n7134 , n7135 , n7136 , n7137 , n7138 , n7139 , n7140 , n7141 , n7142 ,
     n7143 , n7144 , n7145 , n7146 , n7147 , n7148 , n7149 , n7150 , n7151 , n7152 ,
     n7153 , n7154 , n7155 , n7156 , n7157 , n7158 , n7159 , n7160 , n7161 , n7162 ,
     n7163 , n7164 , n7165 , n7166 , n7167 , n7168 , n7169 , n7170 , n7171 , n7172 ,
     n7173 , n7174 , n7175 , n7176 , n7177 , n7178 , n7179 , n7180 , n7181 , n7182 ,
     n7183 , n7184 , n7185 , n7186 , n7187 , n7188 , n7189 , n7190 , n7191 , n7192 ,
     n7193 , n7194 , n7195 , n7196 , n7197 , n7198 , n7199 , n7200 , n7201 , n7202 ,
     n7203 , n7204 , n7205 , n7206 , n7207 , n7208 , n7209 , n7210 , n7211 , n7212 ,
     n7213 , n7214 , n7215 , n7216 , n7217 , n7218 , n7219 , n7220 , n7221 , n7222 ,
     n7223 , n7224 , n7225 , n7226 , n7227 , n7228 , n7229 , n7230 , n7231 , n7232 ,
     n7233 , n7234 , n7235 , n7236 , n7237 , n7238 , n7239 , n7240 , n7241 , n7242 ,
     n7243 , n7244 , n7245 , n7246 , n7247 , n7248 , n7249 , n7250 , n7251 , n7252 ,
     n7253 , n7254 , n7255 , n7256 , n7257 , n7258 , n7259 , n7260 , n7261 , n7262 ,
     n7263 , n7264 , n7265 , n7266 , n7267 , n7268 , n7269 , n7270 , n7271 , n7272 ,
     n7273 , n7274 , n7275 , n7276 , n7277 , n7278 , n7279 , n7280 , n7281 , n7282 ,
     n7283 , n7284 , n7285 , n7286 , n7287 , n7288 , n7289 , n7290 , n7291 , n7292 ,
     n7293 , n7294 , n7295 , n7296 , n7297 , n7298 , n7299 , n7300 , n7301 , n7302 ,
     n7303 , n7304 , n7305 , n7306 , n7307 , n7308 , n7309 , n7310 , n7311 , n7312 ,
     n7313 , n7314 , n7315 , n7316 , n7317 , n7318 , n7319 , n7320 , n7321 , n7322 ,
     n7323 , n7324 , n7325 , n7326 , n7327 , n7328 , n7329 , n7330 , n7331 , n7332 ,
     n7333 , n7334 , n7335 , n7336 , n7337 , n7338 , n7339 , n7340 , n7341 , n7342 ,
     n7343 , n7344 , n7345 , n7346 , n7347 , n7348 , n7349 , n7350 , n7351 , n7352 ,
     n7353 , n7354 , n7355 , n7356 , n7357 , n7358 , n7359 , n7360 , n7361 , n7362 ,
     n7363 , n7364 , n7365 , n7366 , n7367 , n7368 , n7369 , n7370 , n7371 , n7372 ,
     n7373 , n7374 , n7375 , n7376 , n7377 , n7378 , n7379 , n7380 , n7381 , n7382 ,
     n7383 , n7384 , n7385 , n7386 , n7387 , n7388 , n7389 , n7390 , n7391 , n7392 ,
     n7393 , n7394 , n7395 , n7396 , n7397 , n7398 , n7399 , n7400 , n7401 , n7402 ,
     n7403 , n7404 , n7405 , n7406 , n7407 , n7408 , n7409 , n7410 , n7411 , n7412 ,
     n7413 , n7414 , n7415 , n7416 , n7417 , n7418 , n7419 , n7420 , n7421 , n7422 ,
     n7423 , n7424 , n7425 , n7426 , n7427 , n7428 , n7429 , n7430 , n7431 , n7432 ,
     n7433 , n7434 , n7435 , n7436 , n7437 , n7438 , n7439 , n7440 , n7441 , n7442 ,
     n7443 , n7444 , n7445 , n7446 , n7447 , n7448 , n7449 , n7450 , n7451 , n7452 ,
     n7453 , n7454 , n7455 , n7456 , n7457 , n7458 , n7459 , n7460 , n7461 , n7462 ,
     n7463 , n7464 , n7465 , n7466 , n7467 , n7468 , n7469 , n7470 , n7471 , n7472 ,
     n7473 , n7474 , n7475 , n7476 , n7477 , n7478 , n7479 , n7480 , n7481 , n7482 ,
     n7483 , n7484 , n7485 , n7486 , n7487 , n7488 , n7489 , n7490 , n7491 , n7492 ,
     n7493 , n7494 , n7495 , n7496 , n7497 , n7498 , n7499 , n7500 , n7501 , n7502 ,
     n7503 , n7504 , n7505 , n7506 , n7507 , n7508 , n7509 , n7510 , n7511 , n7512 ,
     n7513 , n7514 , n7515 , n7516 , n7517 , n7518 , n7519 , n7520 , n7521 , n7522 ,
     n7523 , n7524 , n7525 , n7526 , n7527 , n7528 , n7529 , n7530 , n7531 , n7532 ,
     n7533 , n7534 , n7535 , n7536 , n7537 , n7538 , n7539 , n7540 , n7541 , n7542 ,
     n7543 , n7544 , n7545 , n7546 , n7547 , n7548 , n7549 , n7550 , n7551 , n7552 ,
     n7553 , n7554 , n7555 , n7556 , n7557 , n7558 , n7559 , n7560 , n7561 , n7562 ,
     n7563 , n7564 , n7565 , n7566 , n7567 , n7568 , n7569 , n7570 , n7571 , n7572 ,
     n7573 , n7574 , n7575 , n7576 , n7577 , n7578 , n7579 , n7580 , n7581 , n7582 ,
     n7583 , n7584 , n7585 , n7586 , n7587 , n7588 , n7589 , n7590 , n7591 , n7592 ,
     n7593 , n7594 , n7595 , n7596 , n7597 , n7598 , n7599 , n7600 , n7601 , n7602 ,
     n7603 , n7604 , n7605 , n7606 , n7607 , n7608 , n7609 , n7610 , n7611 , n7612 ,
     n7613 , n7614 , n7615 , n7616 , n7617 , n7618 , n7619 , n7620 , n7621 , n7622 ,
     n7623 , n7624 , n7625 , n7626 , n7627 , n7628 , n7629 , n7630 , n7631 , n7632 ,
     n7633 , n7634 , n7635 , n7636 , n7637 , n7638 , n7639 , n7640 , n7641 , n7642 ,
     n7643 , n7644 , n7645 , n7646 , n7647 , n7648 , n7649 , n7650 , n7651 , n7652 ,
     n7653 , n7654 , n7655 , n7656 , n7657 , n7658 , n7659 , n7660 , n7661 , n7662 ,
     n7663 , n7664 , n7665 , n7666 , n7667 , n7668 , n7669 , n7670 , n7671 , n7672 ,
     n7673 , n7674 , n7675 , n7676 , n7677 , n7678 , n7679 , n7680 , n7681 , n7682 ,
     n7683 , n7684 , n7685 , n7686 , n7687 , n7688 , n7689 , n7690 , n7691 , n7692 ,
     n7693 , n7694 , n7695 , n7696 , n7697 , n7698 , n7699 , n7700 , n7701 , n7702 ,
     n7703 , n7704 , n7705 , n7706 , n7707 , n7708 , n7709 , n7710 , n7711 , n7712 ,
     n7713 , n7714 , n7715 , n7716 , n7717 , n7718 , n7719 , n7720 , n7721 , n7722 ,
     n7723 , n7724 , n7725 , n7726 , n7727 , n7728 , n7729 , n7730 , n7731 , n7732 ,
     n7733 , n7734 , n7735 , n7736 , n7737 , n7738 , n7739 , n7740 , n7741 , n7742 ,
     n7743 , n7744 , n7745 , n7746 , n7747 , n7748 , n7749 , n7750 , n7751 , n7752 ,
     n7753 , n7754 , n7755 , n7756 , n7757 , n7758 , n7759 , n7760 , n7761 , n7762 ,
     n7763 , n7764 , n7765 , n7766 , n7767 , n7768 , n7769 , n7770 , n7771 , n7772 ,
     n7773 , n7774 , n7775 , n7776 , n7777 , n7778 , n7779 , n7780 , n7781 , n7782 ,
     n7783 , n7784 , n7785 , n7786 , n7787 , n7788 , n7789 , n7790 , n7791 , n7792 ,
     n7793 , n7794 , n7795 , n7796 , n7797 , n7798 , n7799 , n7800 , n7801 , n7802 ,
     n7803 , n7804 , n7805 , n7806 , n7807 , n7808 , n7809 , n7810 , n7811 , n7812 ,
     n7813 , n7814 , n7815 , n7816 , n7817 , n7818 , n7819 , n7820 , n7821 , n7822 ,
     n7823 , n7824 , n7825 , n7826 , n7827 , n7828 , n7829 , n7830 , n7831 , n7832 ,
     n7833 , n7834 , n7835 , n7836 , n7837 , n7838 , n7839 , n7840 , n7841 , n7842 ,
     n7843 , n7844 , n7845 , n7846 , n7847 , n7848 , n7849 , n7850 , n7851 , n7852 ,
     n7853 , n7854 , n7855 , n7856 , n7857 , n7858 , n7859 , n7860 , n7861 , n7862 ,
     n7863 , n7864 , n7865 , n7866 , n7867 , n7868 , n7869 , n7870 , n7871 , n7872 ,
     n7873 , n7874 , n7875 , n7876 , n7877 , n7878 , n7879 , n7880 , n7881 , n7882 ,
     n7883 , n7884 , n7885 , n7886 , n7887 , n7888 , n7889 , n7890 , n7891 , n7892 ,
     n7893 , n7894 , n7895 , n7896 , n7897 , n7898 , n7899 , n7900 , n7901 , n7902 ,
     n7903 , n7904 , n7905 , n7906 , n7907 , n7908 , n7909 , n7910 , n7911 , n7912 ,
     n7913 , n7914 , n7915 , n7916 , n7917 , n7918 , n7919 , n7920 , n7921 , n7922 ,
     n7923 , n7924 , n7925 , n7926 , n7927 , n7928 , n7929 , n7930 , n7931 , n7932 ,
     n7933 , n7934 , n7935 , n7936 , n7937 , n7938 , n7939 , n7940 , n7941 , n7942 ,
     n7943 , n7944 , n7945 , n7946 , n7947 , n7948 , n7949 , n7950 , n7951 , n7952 ,
     n7953 , n7954 , n7955 , n7956 , n7957 , n7958 , n7959 , n7960 , n7961 , n7962 ,
     n7963 , n7964 , n7965 , n7966 , n7967 , n7968 , n7969 , n7970 , n7971 , n7972 ,
     n7973 , n7974 , n7975 , n7976 , n7977 , n7978 , n7979 , n7980 , n7981 , n7982 ,
     n7983 , n7984 , n7985 , n7986 , n7987 , n7988 , n7989 , n7990 , n7991 , n7992 ,
     n7993 , n7994 , n7995 , n7996 , n7997 , n7998 , n7999 , n8000 , n8001 , n8002 ,
     n8003 , n8004 , n8005 , n8006 , n8007 , n8008 , n8009 , n8010 , n8011 , n8012 ,
     n8013 , n8014 , n8015 , n8016 , n8017 , n8018 , n8019 , n8020 , n8021 , n8022 ,
     n8023 , n8024 , n8025 , n8026 , n8027 , n8028 , n8029 , n8030 , n8031 , n8032 ,
     n8033 , n8034 , n8035 , n8036 , n8037 , n8038 , n8039 , n8040 , n8041 , n8042 ,
     n8043 , n8044 , n8045 , n8046 , n8047 , n8048 , n8049 , n8050 , n8051 , n8052 ,
     n8053 , n8054 , n8055 , n8056 , n8057 , n8058 , n8059 , n8060 , n8061 , n8062 ,
     n8063 , n8064 , n8065 , n8066 , n8067 , n8068 , n8069 , n8070 , n8071 , n8072 ,
     n8073 , n8074 , n8075 , n8076 , n8077 , n8078 , n8079 , n8080 , n8081 , n8082 ,
     n8083 , n8084 , n8085 , n8086 , n8087 , n8088 , n8089 , n8090 , n8091 , n8092 ,
     n8093 , n8094 , n8095 , n8096 , n8097 , n8098 , n8099 , n8100 , n8101 , n8102 ,
     n8103 , n8104 , n8105 , n8106 , n8107 , n8108 , n8109 , n8110 , n8111 , n8112 ,
     n8113 , n8114 , n8115 , n8116 , n8117 , n8118 , n8119 , n8120 , n8121 , n8122 ,
     n8123 , n8124 , n8125 , n8126 , n8127 , n8128 , n8129 , n8130 , n8131 , n8132 ,
     n8133 , n8134 , n8135 , n8136 , n8137 , n8138 , n8139 , n8140 , n8141 , n8142 ,
     n8143 , n8144 , n8145 , n8146 , n8147 , n8148 , n8149 , n8150 , n8151 , n8152 ,
     n8153 , n8154 , n8155 , n8156 , n8157 , n8158 , n8159 , n8160 , n8161 , n8162 ,
     n8163 , n8164 , n8165 , n8166 , n8167 , n8168 , n8169 , n8170 , n8171 , n8172 ,
     n8173 , n8174 , n8175 , n8176 , n8177 , n8178 , n8179 , n8180 , n8181 , n8182 ,
     n8183 , n8184 , n8185 , n8186 , n8187 , n8188 , n8189 , n8190 , n8191 , n8192 ,
     n8193 , n8194 , n8195 , n8196 , n8197 , n8198 , n8199 , n8200 , n8201 , n8202 ,
     n8203 , n8204 , n8205 , n8206 , n8207 , n8208 , n8209 , n8210 , n8211 , n8212 ,
     n8213 , n8214 , n8215 , n8216 , n8217 , n8218 , n8219 , n8220 , n8221 , n8222 ,
     n8223 , n8224 , n8225 , n8226 , n8227 , n8228 , n8229 , n8230 , n8231 , n8232 ,
     n8233 , n8234 , n8235 , n8236 , n8237 , n8238 , n8239 , n8240 , n8241 , n8242 ,
     n8243 , n8244 , n8245 , n8246 , n8247 , n8248 , n8249 , n8250 , n8251 , n8252 ,
     n8253 , n8254 , n8255 , n8256 , n8257 , n8258 , n8259 , n8260 , n8261 , n8262 ,
     n8263 , n8264 , n8265 , n8266 , n8267 , n8268 , n8269 , n8270 , n8271 , n8272 ,
     n8273 , n8274 , n8275 , n8276 , n8277 , n8278 , n8279 , n8280 , n8281 , n8282 ,
     n8283 , n8284 , n8285 , n8286 , n8287 , n8288 , n8289 , n8290 , n8291 , n8292 ,
     n8293 , n8294 , n8295 , n8296 , n8297 , n8298 , n8299 , n8300 , n8301 , n8302 ,
     n8303 , n8304 , n8305 , n8306 , n8307 , n8308 , n8309 , n8310 , n8311 , n8312 ,
     n8313 , n8314 , n8315 , n8316 , n8317 , n8318 , n8319 , n8320 , n8321 , n8322 ,
     n8323 , n8324 , n8325 , n8326 , n8327 , n8328 , n8329 , n8330 , n8331 , n8332 ,
     n8333 , n8334 , n8335 , n8336 , n8337 , n8338 , n8339 , n8340 , n8341 , n8342 ,
     n8343 , n8344 , n8345 , n8346 , n8347 , n8348 , n8349 , n8350 , n8351 , n8352 ,
     n8353 , n8354 , n8355 , n8356 , n8357 , n8358 , n8359 , n8360 , n8361 , n8362 ,
     n8363 , n8364 , n8365 , n8366 , n8367 , n8368 , n8369 , n8370 , n8371 , n8372 ,
     n8373 , n8374 , n8375 , n8376 , n8377 , n8378 , n8379 , n8380 , n8381 , n8382 ,
     n8383 , n8384 , n8385 , n8386 , n8387 , n8388 , n8389 , n8390 , n8391 , n8392 ,
     n8393 , n8394 , n8395 , n8396 , n8397 , n8398 , n8399 , n8400 , n8401 , n8402 ,
     n8403 , n8404 , n8405 , n8406 , n8407 , n8408 , n8409 , n8410 , n8411 , n8412 ,
     n8413 , n8414 , n8415 , n8416 , n8417 , n8418 , n8419 , n8420 , n8421 , n8422 ,
     n8423 , n8424 , n8425 , n8426 , n8427 , n8428 , n8429 , n8430 , n8431 , n8432 ,
     n8433 , n8434 , n8435 , n8436 , n8437 , n8438 , n8439 , n8440 , n8441 , n8442 ,
     n8443 , n8444 , n8445 , n8446 , n8447 , n8448 , n8449 , n8450 , n8451 , n8452 ,
     n8453 , n8454 , n8455 , n8456 , n8457 , n8458 , n8459 , n8460 , n8461 , n8462 ,
     n8463 , n8464 , n8465 , n8466 , n8467 , n8468 , n8469 , n8470 , n8471 , n8472 ,
     n8473 , n8474 , n8475 , n8476 , n8477 , n8478 , n8479 , n8480 , n8481 , n8482 ,
     n8483 , n8484 , n8485 , n8486 , n8487 , n8488 , n8489 , n8490 , n8491 , n8492 ,
     n8493 , n8494 , n8495 , n8496 , n8497 , n8498 , n8499 , n8500 , n8501 , n8502 ,
     n8503 , n8504 , n8505 , n8506 , n8507 , n8508 , n8509 , n8510 , n8511 , n8512 ,
     n8513 , n8514 , n8515 , n8516 , n8517 , n8518 , n8519 , n8520 , n8521 , n8522 ,
     n8523 , n8524 , n8525 , n8526 , n8527 , n8528 , n8529 , n8530 , n8531 , n8532 ,
     n8533 , n8534 , n8535 , n8536 , n8537 , n8538 , n8539 , n8540 , n8541 , n8542 ,
     n8543 , n8544 , n8545 , n8546 , n8547 , n8548 , n8549 , n8550 , n8551 , n8552 ,
     n8553 , n8554 , n8555 , n8556 , n8557 , n8558 , n8559 , n8560 , n8561 , n8562 ,
     n8563 , n8564 , n8565 , n8566 , n8567 , n8568 , n8569 , n8570 , n8571 , n8572 ,
     n8573 , n8574 , n8575 , n8576 , n8577 , n8578 , n8579 , n8580 , n8581 , n8582 ,
     n8583 , n8584 , n8585 , n8586 , n8587 , n8588 , n8589 , n8590 , n8591 , n8592 ,
     n8593 , n8594 , n8595 , n8596 , n8597 , n8598 , n8599 , n8600 , n8601 , n8602 ,
     n8603 , n8604 , n8605 , n8606 , n8607 , n8608 , n8609 , n8610 , n8611 , n8612 ,
     n8613 , n8614 , n8615 , n8616 , n8617 , n8618 , n8619 , n8620 , n8621 , n8622 ,
     n8623 , n8624 , n8625 , n8626 , n8627 , n8628 , n8629 , n8630 , n8631 , n8632 ,
     n8633 , n8634 , n8635 , n8636 , n8637 , n8638 , n8639 , n8640 , n8641 , n8642 ,
     n8643 , n8644 , n8645 , n8646 , n8647 , n8648 , n8649 , n8650 , n8651 , n8652 ,
     n8653 , n8654 , n8655 , n8656 , n8657 , n8658 , n8659 , n8660 , n8661 , n8662 ,
     n8663 , n8664 , n8665 , n8666 , n8667 , n8668 , n8669 , n8670 , n8671 , n8672 ,
     n8673 , n8674 , n8675 , n8676 , n8677 , n8678 , n8679 , n8680 , n8681 , n8682 ,
     n8683 , n8684 , n8685 , n8686 , n8687 , n8688 , n8689 , n8690 , n8691 , n8692 ,
     n8693 , n8694 , n8695 , n8696 , n8697 , n8698 , n8699 , n8700 , n8701 , n8702 ,
     n8703 , n8704 , n8705 , n8706 , n8707 , n8708 , n8709 , n8710 , n8711 , n8712 ,
     n8713 , n8714 , n8715 , n8716 , n8717 , n8718 , n8719 , n8720 , n8721 , n8722 ,
     n8723 , n8724 , n8725 , n8726 , n8727 , n8728 , n8729 , n8730 , n8731 , n8732 ,
     n8733 , n8734 , n8735 , n8736 , n8737 , n8738 , n8739 , n8740 , n8741 , n8742 ,
     n8743 , n8744 , n8745 , n8746 , n8747 , n8748 , n8749 , n8750 , n8751 , n8752 ,
     n8753 , n8754 , n8755 , n8756 , n8757 , n8758 , n8759 , n8760 , n8761 , n8762 ,
     n8763 , n8764 , n8765 , n8766 , n8767 , n8768 , n8769 , n8770 , n8771 , n8772 ,
     n8773 , n8774 , n8775 , n8776 , n8777 , n8778 , n8779 , n8780 , n8781 , n8782 ,
     n8783 , n8784 , n8785 , n8786 , n8787 , n8788 , n8789 , n8790 , n8791 , n8792 ,
     n8793 , n8794 , n8795 , n8796 , n8797 , n8798 , n8799 , n8800 , n8801 , n8802 ,
     n8803 , n8804 , n8805 , n8806 , n8807 , n8808 , n8809 , n8810 , n8811 , n8812 ,
     n8813 , n8814 , n8815 , n8816 , n8817 , n8818 , n8819 , n8820 , n8821 , n8822 ,
     n8823 , n8824 , n8825 , n8826 , n8827 , n8828 , n8829 , n8830 , n8831 , n8832 ,
     n8833 , n8834 , n8835 , n8836 , n8837 , n8838 , n8839 , n8840 , n8841 , n8842 ,
     n8843 , n8844 , n8845 , n8846 , n8847 , n8848 , n8849 , n8850 , n8851 , n8852 ,
     n8853 , n8854 , n8855 , n8856 , n8857 , n8858 , n8859 , n8860 , n8861 , n8862 ,
     n8863 , n8864 , n8865 , n8866 , n8867 , n8868 , n8869 , n8870 , n8871 , n8872 ,
     n8873 , n8874 , n8875 , n8876 , n8877 , n8878 , n8879 , n8880 , n8881 , n8882 ,
     n8883 , n8884 , n8885 , n8886 , n8887 , n8888 , n8889 , n8890 , n8891 , n8892 ,
     n8893 , n8894 , n8895 , n8896 , n8897 , n8898 , n8899 , n8900 , n8901 , n8902 ,
     n8903 , n8904 , n8905 , n8906 , n8907 , n8908 , n8909 , n8910 , n8911 , n8912 ,
     n8913 , n8914 , n8915 , n8916 , n8917 , n8918 , n8919 , n8920 , n8921 , n8922 ,
     n8923 , n8924 , n8925 , n8926 , n8927 , n8928 , n8929 , n8930 , n8931 , n8932 ,
     n8933 , n8934 , n8935 , n8936 , n8937 , n8938 , n8939 , n8940 , n8941 , n8942 ,
     n8943 , n8944 , n8945 , n8946 , n8947 , n8948 , n8949 , n8950 , n8951 , n8952 ,
     n8953 , n8954 , n8955 , n8956 , n8957 , n8958 , n8959 , n8960 , n8961 , n8962 ,
     n8963 , n8964 , n8965 , n8966 , n8967 , n8968 , n8969 , n8970 , n8971 , n8972 ,
     n8973 , n8974 , n8975 , n8976 , n8977 , n8978 , n8979 , n8980 , n8981 , n8982 ,
     n8983 , n8984 , n8985 , n8986 , n8987 , n8988 , n8989 , n8990 , n8991 , n8992 ,
     n8993 , n8994 , n8995 , n8996 , n8997 , n8998 , n8999 , n9000 , n9001 , n9002 ,
     n9003 , n9004 , n9005 , n9006 , n9007 , n9008 , n9009 , n9010 , n9011 , n9012 ,
     n9013 , n9014 , n9015 , n9016 , n9017 , n9018 , n9019 , n9020 , n9021 , n9022 ,
     n9023 , n9024 , n9025 , n9026 , n9027 , n9028 , n9029 , n9030 , n9031 , n9032 ,
     n9033 , n9034 , n9035 , n9036 , n9037 , n9038 , n9039 , n9040 , n9041 , n9042 ,
     n9043 , n9044 , n9045 , n9046 , n9047 , n9048 , n9049 , n9050 , n9051 , n9052 ,
     n9053 , n9054 , n9055 , n9056 , n9057 , n9058 , n9059 , n9060 , n9061 , n9062 ,
     n9063 , n9064 , n9065 , n9066 , n9067 , n9068 , n9069 , n9070 , n9071 , n9072 ,
     n9073 , n9074 , n9075 , n9076 , n9077 , n9078 , n9079 , n9080 , n9081 , n9082 ,
     n9083 , n9084 , n9085 , n9086 , n9087 , n9088 , n9089 , n9090 , n9091 , n9092 ,
     n9093 , n9094 , n9095 , n9096 , n9097 , n9098 , n9099 , n9100 , n9101 , n9102 ,
     n9103 , n9104 , n9105 , n9106 , n9107 , n9108 , n9109 , n9110 , n9111 , n9112 ,
     n9113 , n9114 , n9115 , n9116 , n9117 , n9118 , n9119 , n9120 , n9121 , n9122 ,
     n9123 , n9124 , n9125 , n9126 , n9127 , n9128 , n9129 , n9130 , n9131 , n9132 ,
     n9133 , n9134 , n9135 , n9136 , n9137 , n9138 , n9139 , n9140 , n9141 , n9142 ,
     n9143 , n9144 , n9145 , n9146 , n9147 , n9148 , n9149 , n9150 , n9151 , n9152 ,
     n9153 , n9154 , n9155 , n9156 , n9157 , n9158 , n9159 , n9160 , n9161 , n9162 ,
     n9163 , n9164 , n9165 , n9166 , n9167 , n9168 , n9169 , n9170 , n9171 , n9172 ,
     n9173 , n9174 , n9175 , n9176 , n9177 , n9178 , n9179 , n9180 , n9181 , n9182 ,
     n9183 , n9184 , n9185 , n9186 , n9187 , n9188 , n9189 , n9190 , n9191 , n9192 ,
     n9193 , n9194 , n9195 , n9196 , n9197 , n9198 , n9199 , n9200 , n9201 , n9202 ,
     n9203 , n9204 , n9205 , n9206 , n9207 , n9208 , n9209 , n9210 , n9211 , n9212 ,
     n9213 , n9214 , n9215 , n9216 , n9217 , n9218 , n9219 , n9220 , n9221 , n9222 ,
     n9223 , n9224 , n9225 , n9226 , n9227 , n9228 , n9229 , n9230 , n9231 , n9232 ,
     n9233 , n9234 , n9235 , n9236 , n9237 , n9238 , n9239 , n9240 , n9241 , n9242 ,
     n9243 , n9244 , n9245 , n9246 , n9247 , n9248 , n9249 , n9250 , n9251 , n9252 ,
     n9253 , n9254 , n9255 , n9256 , n9257 , n9258 , n9259 , n9260 , n9261 , n9262 ,
     n9263 , n9264 , n9265 , n9266 , n9267 , n9268 , n9269 , n9270 , n9271 , n9272 ,
     n9273 , n9274 , n9275 , n9276 , n9277 , n9278 , n9279 , n9280 , n9281 , n9282 ,
     n9283 , n9284 , n9285 , n9286 , n9287 , n9288 , n9289 , n9290 , n9291 , n9292 ,
     n9293 , n9294 , n9295 , n9296 , n9297 , n9298 , n9299 , n9300 , n9301 , n9302 ,
     n9303 , n9304 , n9305 , n9306 , n9307 , n9308 , n9309 , n9310 , n9311 , n9312 ,
     n9313 , n9314 , n9315 , n9316 , n9317 , n9318 , n9319 , n9320 , n9321 , n9322 ,
     n9323 , n9324 , n9325 , n9326 , n9327 , n9328 , n9329 , n9330 , n9331 , n9332 ,
     n9333 , n9334 , n9335 , n9336 , n9337 , n9338 , n9339 , n9340 , n9341 , n9342 ,
     n9343 , n9344 , n9345 , n9346 , n9347 , n9348 , n9349 , n9350 , n9351 , n9352 ,
     n9353 , n9354 , n9355 , n9356 , n9357 , n9358 , n9359 , n9360 , n9361 , n9362 ,
     n9363 , n9364 , n9365 , n9366 , n9367 , n9368 , n9369 , n9370 , n9371 , n9372 ,
     n9373 , n9374 , n9375 , n9376 , n9377 , n9378 , n9379 , n9380 , n9381 , n9382 ,
     n9383 , n9384 , n9385 , n9386 , n9387 , n9388 , n9389 , n9390 , n9391 , n9392 ,
     n9393 , n9394 , n9395 , n9396 , n9397 , n9398 , n9399 , n9400 , n9401 , n9402 ,
     n9403 , n9404 , n9405 , n9406 , n9407 , n9408 , n9409 , n9410 , n9411 , n9412 ,
     n9413 , n9414 , n9415 , n9416 , n9417 , n9418 , n9419 , n9420 , n9421 , n9422 ,
     n9423 , n9424 , n9425 , n9426 , n9427 , n9428 , n9429 , n9430 , n9431 , n9432 ,
     n9433 , n9434 , n9435 , n9436 , n9437 , n9438 , n9439 , n9440 , n9441 , n9442 ,
     n9443 , n9444 , n9445 , n9446 , n9447 , n9448 , n9449 , n9450 , n9451 , n9452 ,
     n9453 , n9454 , n9455 , n9456 , n9457 , n9458 , n9459 , n9460 , n9461 , n9462 ,
     n9463 , n9464 , n9465 , n9466 , n9467 , n9468 , n9469 , n9470 , n9471 , n9472 ,
     n9473 , n9474 , n9475 , n9476 , n9477 , n9478 , n9479 , n9480 , n9481 , n9482 ,
     n9483 , n9484 , n9485 , n9486 , n9487 , n9488 , n9489 , n9490 , n9491 , n9492 ,
     n9493 , n9494 , n9495 , n9496 , n9497 , n9498 , n9499 , n9500 , n9501 , n9502 ,
     n9503 , n9504 , n9505 , n9506 , n9507 , n9508 , n9509 , n9510 , n9511 , n9512 ,
     n9513 , n9514 , n9515 , n9516 , n9517 , n9518 , n9519 , n9520 , n9521 , n9522 ,
     n9523 , n9524 , n9525 , n9526 , n9527 , n9528 , n9529 , n9530 , n9531 , n9532 ,
     n9533 , n9534 , n9535 , n9536 , n9537 , n9538 , n9539 , n9540 , n9541 , n9542 ,
     n9543 , n9544 , n9545 , n9546 , n9547 , n9548 , n9549 , n9550 , n9551 , n9552 ,
     n9553 , n9554 , n9555 , n9556 , n9557 , n9558 , n9559 , n9560 , n9561 , n9562 ,
     n9563 , n9564 , n9565 , n9566 , n9567 , n9568 , n9569 , n9570 , n9571 , n9572 ,
     n9573 , n9574 , n9575 , n9576 , n9577 , n9578 , n9579 , n9580 , n9581 , n9582 ,
     n9583 , n9584 , n9585 , n9586 , n9587 , n9588 , n9589 , n9590 , n9591 , n9592 ,
     n9593 , n9594 , n9595 , n9596 , n9597 , n9598 , n9599 , n9600 , n9601 , n9602 ,
     n9603 , n9604 , n9605 , n9606 , n9607 , n9608 , n9609 , n9610 , n9611 , n9612 ,
     n9613 , n9614 , n9615 , n9616 , n9617 , n9618 , n9619 , n9620 , n9621 , n9622 ,
     n9623 , n9624 , n9625 , n9626 , n9627 , n9628 , n9629 , n9630 , n9631 , n9632 ,
     n9633 , n9634 , n9635 , n9636 , n9637 , n9638 , n9639 , n9640 , n9641 , n9642 ,
     n9643 , n9644 , n9645 , n9646 , n9647 , n9648 , n9649 , n9650 , n9651 , n9652 ,
     n9653 , n9654 , n9655 , n9656 , n9657 , n9658 , n9659 , n9660 , n9661 , n9662 ,
     n9663 , n9664 , n9665 , n9666 , n9667 , n9668 , n9669 , n9670 , n9671 , n9672 ,
     n9673 , n9674 , n9675 , n9676 , n9677 , n9678 , n9679 , n9680 , n9681 , n9682 ,
     n9683 , n9684 , n9685 , n9686 , n9687 , n9688 , n9689 , n9690 , n9691 , n9692 ,
     n9693 , n9694 , n9695 , n9696 , n9697 , n9698 , n9699 , n9700 , n9701 , n9702 ,
     n9703 , n9704 , n9705 , n9706 , n9707 , n9708 , n9709 , n9710 , n9711 , n9712 ,
     n9713 , n9714 , n9715 , n9716 , n9717 , n9718 , n9719 , n9720 , n9721 , n9722 ,
     n9723 , n9724 , n9725 , n9726 , n9727 , n9728 , n9729 , n9730 , n9731 , n9732 ,
     n9733 , n9734 , n9735 , n9736 , n9737 , n9738 , n9739 , n9740 , n9741 , n9742 ,
     n9743 , n9744 , n9745 , n9746 , n9747 , n9748 , n9749 , n9750 , n9751 , n9752 ,
     n9753 , n9754 , n9755 , n9756 , n9757 , n9758 , n9759 , n9760 , n9761 , n9762 ,
     n9763 , n9764 , n9765 , n9766 , n9767 , n9768 , n9769 , n9770 , n9771 , n9772 ,
     n9773 , n9774 , n9775 , n9776 , n9777 , n9778 , n9779 , n9780 , n9781 , n9782 ,
     n9783 , n9784 , n9785 , n9786 , n9787 , n9788 , n9789 , n9790 , n9791 , n9792 ,
     n9793 , n9794 , n9795 , n9796 , n9797 , n9798 , n9799 , n9800 , n9801 , n9802 ,
     n9803 , n9804 , n9805 , n9806 , n9807 , n9808 , n9809 , n9810 , n9811 , n9812 ,
     n9813 , n9814 , n9815 , n9816 , n9817 , n9818 , n9819 , n9820 , n9821 , n9822 ,
     n9823 , n9824 , n9825 , n9826 , n9827 , n9828 , n9829 , n9830 , n9831 , n9832 ,
     n9833 , n9834 , n9835 , n9836 , n9837 , n9838 , n9839 , n9840 , n9841 , n9842 ,
     n9843 , n9844 , n9845 , n9846 , n9847 , n9848 , n9849 , n9850 , n9851 , n9852 ,
     n9853 , n9854 , n9855 , n9856 , n9857 , n9858 , n9859 , n9860 , n9861 , n9862 ,
     n9863 , n9864 , n9865 , n9866 , n9867 , n9868 , n9869 , n9870 , n9871 , n9872 ,
     n9873 , n9874 , n9875 , n9876 , n9877 , n9878 , n9879 , n9880 , n9881 , n9882 ,
     n9883 , n9884 , n9885 , n9886 , n9887 , n9888 , n9889 , n9890 , n9891 , n9892 ,
     n9893 , n9894 , n9895 , n9896 , n9897 , n9898 , n9899 , n9900 , n9901 , n9902 ,
     n9903 , n9904 , n9905 , n9906 , n9907 , n9908 , n9909 , n9910 , n9911 , n9912 ,
     n9913 , n9914 , n9915 , n9916 , n9917 , n9918 , n9919 , n9920 , n9921 , n9922 ,
     n9923 , n9924 , n9925 , n9926 , n9927 , n9928 , n9929 , n9930 , n9931 , n9932 ,
     n9933 , n9934 , n9935 , n9936 , n9937 , n9938 , n9939 , n9940 , n9941 , n9942 ,
     n9943 , n9944 , n9945 , n9946 , n9947 , n9948 , n9949 , n9950 , n9951 , n9952 ,
     n9953 , n9954 , n9955 , n9956 , n9957 , n9958 , n9959 , n9960 , n9961 , n9962 ,
     n9963 , n9964 , n9965 , n9966 , n9967 , n9968 , n9969 , n9970 , n9971 , n9972 ,
     n9973 , n9974 , n9975 , n9976 , n9977 , n9978 , n9979 , n9980 , n9981 , n9982 ,
     n9983 , n9984 , n9985 , n9986 , n9987 , n9988 , n9989 , n9990 , n9991 , n9992 ,
     n9993 , n9994 , n9995 , n9996 , n9997 , n9998 , n9999 , n10000 , n10001 , n10002 ,
     n10003 , n10004 , n10005 , n10006 , n10007 , n10008 , n10009 , n10010 , n10011 , n10012 ,
     n10013 , n10014 , n10015 , n10016 , n10017 , n10018 , n10019 , n10020 , n10021 , n10022 ,
     n10023 , n10024 , n10025 , n10026 , n10027 , n10028 , n10029 , n10030 , n10031 , n10032 ,
     n10033 , n10034 , n10035 , n10036 , n10037 , n10038 , n10039 , n10040 , n10041 , n10042 ,
     n10043 , n10044 , n10045 , n10046 , n10047 , n10048 , n10049 , n10050 , n10051 , n10052 ,
     n10053 , n10054 , n10055 , n10056 , n10057 , n10058 , n10059 , n10060 , n10061 , n10062 ,
     n10063 , n10064 , n10065 , n10066 , n10067 , n10068 , n10069 , n10070 , n10071 , n10072 ,
     n10073 , n10074 , n10075 , n10076 , n10077 , n10078 , n10079 , n10080 , n10081 , n10082 ,
     n10083 , n10084 , n10085 , n10086 , n10087 , n10088 , n10089 , n10090 , n10091 , n10092 ,
     n10093 , n10094 , n10095 , n10096 , n10097 , n10098 , n10099 , n10100 , n10101 , n10102 ,
     n10103 , n10104 , n10105 , n10106 , n10107 , n10108 , n10109 , n10110 , n10111 , n10112 ,
     n10113 , n10114 , n10115 , n10116 , n10117 , n10118 , n10119 , n10120 , n10121 , n10122 ,
     n10123 , n10124 , n10125 , n10126 , n10127 , n10128 , n10129 , n10130 , n10131 , n10132 ,
     n10133 , n10134 , n10135 , n10136 , n10137 , n10138 , n10139 , n10140 , n10141 , n10142 ,
     n10143 , n10144 , n10145 , n10146 , n10147 , n10148 , n10149 , n10150 , n10151 , n10152 ,
     n10153 , n10154 , n10155 , n10156 , n10157 , n10158 , n10159 , n10160 , n10161 , n10162 ,
     n10163 , n10164 , n10165 , n10166 , n10167 , n10168 , n10169 , n10170 , n10171 , n10172 ,
     n10173 , n10174 , n10175 , n10176 , n10177 , n10178 , n10179 , n10180 , n10181 , n10182 ,
     n10183 , n10184 , n10185 , n10186 , n10187 , n10188 , n10189 , n10190 , n10191 , n10192 ,
     n10193 , n10194 , n10195 , n10196 , n10197 , n10198 , n10199 , n10200 , n10201 , n10202 ,
     n10203 , n10204 , n10205 , n10206 , n10207 , n10208 , n10209 , n10210 , n10211 , n10212 ,
     n10213 , n10214 , n10215 , n10216 , n10217 , n10218 , n10219 , n10220 , n10221 , n10222 ,
     n10223 , n10224 , n10225 , n10226 , n10227 , n10228 , n10229 , n10230 , n10231 , n10232 ,
     n10233 , n10234 , n10235 , n10236 , n10237 , n10238 , n10239 , n10240 , n10241 , n10242 ,
     n10243 , n10244 , n10245 , n10246 , n10247 , n10248 , n10249 , n10250 , n10251 , n10252 ,
     n10253 , n10254 , n10255 , n10256 , n10257 , n10258 , n10259 , n10260 , n10261 , n10262 ,
     n10263 , n10264 , n10265 , n10266 , n10267 , n10268 , n10269 , n10270 , n10271 , n10272 ,
     n10273 , n10274 , n10275 , n10276 , n10277 , n10278 , n10279 , n10280 , n10281 , n10282 ,
     n10283 , n10284 , n10285 , n10286 , n10287 , n10288 , n10289 , n10290 , n10291 , n10292 ,
     n10293 , n10294 , n10295 , n10296 , n10297 , n10298 , n10299 , n10300 , n10301 , n10302 ,
     n10303 , n10304 , n10305 , n10306 , n10307 , n10308 , n10309 , n10310 , n10311 , n10312 ,
     n10313 , n10314 , n10315 , n10316 , n10317 , n10318 , n10319 , n10320 , n10321 , n10322 ,
     n10323 , n10324 , n10325 , n10326 , n10327 , n10328 , n10329 , n10330 , n10331 , n10332 ,
     n10333 , n10334 , n10335 , n10336 , n10337 , n10338 , n10339 , n10340 , n10341 , n10342 ,
     n10343 , n10344 , n10345 , n10346 , n10347 , n10348 , n10349 , n10350 , n10351 , n10352 ,
     n10353 , n10354 , n10355 , n10356 , n10357 , n10358 , n10359 , n10360 , n10361 , n10362 ,
     n10363 , n10364 , n10365 , n10366 , n10367 , n10368 , n10369 , n10370 , n10371 , n10372 ,
     n10373 , n10374 , n10375 , n10376 , n10377 , n10378 , n10379 , n10380 , n10381 , n10382 ,
     n10383 , n10384 , n10385 , n10386 , n10387 , n10388 , n10389 , n10390 , n10391 , n10392 ,
     n10393 , n10394 , n10395 , n10396 , n10397 , n10398 , n10399 , n10400 , n10401 , n10402 ,
     n10403 , n10404 , n10405 , n10406 , n10407 , n10408 , n10409 , n10410 , n10411 , n10412 ,
     n10413 , n10414 , n10415 , n10416 , n10417 , n10418 , n10419 , n10420 , n10421 , n10422 ,
     n10423 , n10424 , n10425 , n10426 , n10427 , n10428 , n10429 , n10430 , n10431 , n10432 ,
     n10433 , n10434 , n10435 , n10436 , n10437 , n10438 , n10439 , n10440 , n10441 , n10442 ,
     n10443 , n10444 , n10445 , n10446 , n10447 , n10448 , n10449 , n10450 , n10451 , n10452 ,
     n10453 , n10454 , n10455 , n10456 , n10457 , n10458 , n10459 , n10460 , n10461 , n10462 ,
     n10463 , n10464 , n10465 , n10466 , n10467 , n10468 , n10469 , n10470 , n10471 , n10472 ,
     n10473 , n10474 , n10475 , n10476 , n10477 , n10478 , n10479 , n10480 , n10481 , n10482 ,
     n10483 , n10484 , n10485 , n10486 , n10487 , n10488 , n10489 , n10490 , n10491 , n10492 ,
     n10493 , n10494 , n10495 , n10496 , n10497 , n10498 , n10499 , n10500 , n10501 , n10502 ,
     n10503 , n10504 , n10505 , n10506 , n10507 , n10508 , n10509 , n10510 , n10511 , n10512 ,
     n10513 , n10514 , n10515 , n10516 , n10517 , n10518 , n10519 , n10520 , n10521 , n10522 ,
     n10523 , n10524 , n10525 , n10526 , n10527 , n10528 , n10529 , n10530 , n10531 , n10532 ,
     n10533 , n10534 , n10535 , n10536 , n10537 , n10538 , n10539 , n10540 , n10541 , n10542 ,
     n10543 , n10544 , n10545 , n10546 , n10547 , n10548 , n10549 , n10550 , n10551 , n10552 ,
     n10553 , n10554 , n10555 , n10556 , n10557 , n10558 , n10559 , n10560 , n10561 , n10562 ,
     n10563 , n10564 , n10565 , n10566 , n10567 , n10568 , n10569 , n10570 , n10571 , n10572 ,
     n10573 , n10574 , n10575 , n10576 , n10577 , n10578 , n10579 , n10580 , n10581 , n10582 ,
     n10583 , n10584 , n10585 , n10586 , n10587 , n10588 , n10589 , n10590 , n10591 , n10592 ,
     n10593 , n10594 , n10595 , n10596 , n10597 , n10598 , n10599 , n10600 , n10601 , n10602 ,
     n10603 , n10604 , n10605 , n10606 , n10607 , n10608 , n10609 , n10610 , n10611 , n10612 ,
     n10613 , n10614 , n10615 , n10616 , n10617 , n10618 , n10619 , n10620 , n10621 , n10622 ,
     n10623 , n10624 , n10625 , n10626 , n10627 , n10628 , n10629 , n10630 , n10631 , n10632 ,
     n10633 , n10634 , n10635 , n10636 , n10637 , n10638 , n10639 , n10640 , n10641 , n10642 ,
     n10643 , n10644 , n10645 , n10646 , n10647 , n10648 , n10649 , n10650 , n10651 , n10652 ,
     n10653 , n10654 , n10655 , n10656 , n10657 , n10658 , n10659 , n10660 , n10661 , n10662 ,
     n10663 , n10664 , n10665 , n10666 , n10667 , n10668 , n10669 , n10670 , n10671 , n10672 ,
     n10673 , n10674 , n10675 , n10676 , n10677 , n10678 , n10679 , n10680 , n10681 , n10682 ,
     n10683 , n10684 , n10685 , n10686 , n10687 , n10688 , n10689 , n10690 , n10691 , n10692 ,
     n10693 , n10694 , n10695 , n10696 , n10697 , n10698 , n10699 , n10700 , n10701 , n10702 ,
     n10703 , n10704 , n10705 , n10706 , n10707 , n10708 , n10709 , n10710 , n10711 , n10712 ,
     n10713 , n10714 , n10715 , n10716 , n10717 , n10718 , n10719 , n10720 , n10721 , n10722 ,
     n10723 , n10724 , n10725 , n10726 , n10727 , n10728 , n10729 , n10730 , n10731 , n10732 ,
     n10733 , n10734 , n10735 , n10736 , n10737 , n10738 , n10739 , n10740 , n10741 , n10742 ,
     n10743 , n10744 , n10745 , n10746 , n10747 , n10748 , n10749 , n10750 , n10751 , n10752 ,
     n10753 , n10754 , n10755 , n10756 , n10757 , n10758 , n10759 , n10760 , n10761 , n10762 ,
     n10763 , n10764 , n10765 , n10766 , n10767 , n10768 , n10769 , n10770 , n10771 , n10772 ,
     n10773 , n10774 , n10775 , n10776 , n10777 , n10778 , n10779 , n10780 , n10781 , n10782 ,
     n10783 , n10784 , n10785 , n10786 , n10787 , n10788 , n10789 , n10790 , n10791 , n10792 ,
     n10793 , n10794 , n10795 , n10796 , n10797 , n10798 , n10799 , n10800 , n10801 , n10802 ,
     n10803 , n10804 , n10805 , n10806 , n10807 , n10808 , n10809 , n10810 , n10811 , n10812 ,
     n10813 , n10814 , n10815 , n10816 , n10817 , n10818 , n10819 , n10820 , n10821 , n10822 ,
     n10823 , n10824 , n10825 , n10826 , n10827 , n10828 , n10829 , n10830 , n10831 , n10832 ,
     n10833 , n10834 , n10835 , n10836 , n10837 , n10838 , n10839 , n10840 , n10841 , n10842 ,
     n10843 , n10844 , n10845 , n10846 , n10847 , n10848 , n10849 , n10850 , n10851 , n10852 ,
     n10853 , n10854 , n10855 , n10856 , n10857 , n10858 , n10859 , n10860 , n10861 , n10862 ,
     n10863 , n10864 , n10865 , n10866 , n10867 , n10868 , n10869 , n10870 , n10871 , n10872 ,
     n10873 , n10874 , n10875 , n10876 , n10877 , n10878 , n10879 , n10880 , n10881 , n10882 ,
     n10883 , n10884 , n10885 , n10886 , n10887 , n10888 , n10889 , n10890 , n10891 , n10892 ,
     n10893 , n10894 , n10895 , n10896 , n10897 , n10898 , n10899 , n10900 , n10901 , n10902 ,
     n10903 , n10904 , n10905 , n10906 , n10907 , n10908 , n10909 , n10910 , n10911 , n10912 ,
     n10913 , n10914 , n10915 , n10916 , n10917 , n10918 , n10919 , n10920 , n10921 , n10922 ,
     n10923 , n10924 , n10925 , n10926 , n10927 , n10928 , n10929 , n10930 , n10931 , n10932 ,
     n10933 , n10934 , n10935 , n10936 , n10937 , n10938 , n10939 , n10940 , n10941 , n10942 ,
     n10943 , n10944 , n10945 , n10946 , n10947 , n10948 , n10949 , n10950 , n10951 , n10952 ,
     n10953 , n10954 , n10955 , n10956 , n10957 , n10958 , n10959 , n10960 , n10961 , n10962 ,
     n10963 , n10964 , n10965 , n10966 , n10967 , n10968 , n10969 , n10970 , n10971 , n10972 ,
     n10973 , n10974 , n10975 , n10976 , n10977 , n10978 , n10979 , n10980 , n10981 , n10982 ,
     n10983 , n10984 , n10985 , n10986 , n10987 , n10988 , n10989 , n10990 , n10991 , n10992 ,
     n10993 , n10994 , n10995 , n10996 , n10997 , n10998 , n10999 , n11000 , n11001 , n11002 ,
     n11003 , n11004 , n11005 , n11006 , n11007 , n11008 , n11009 , n11010 , n11011 , n11012 ,
     n11013 , n11014 , n11015 , n11016 , n11017 , n11018 , n11019 , n11020 , n11021 , n11022 ,
     n11023 , n11024 , n11025 , n11026 , n11027 , n11028 , n11029 , n11030 , n11031 , n11032 ,
     n11033 , n11034 , n11035 , n11036 , n11037 , n11038 , n11039 , n11040 , n11041 , n11042 ,
     n11043 , n11044 , n11045 , n11046 , n11047 , n11048 , n11049 , n11050 , n11051 , n11052 ,
     n11053 , n11054 , n11055 , n11056 , n11057 , n11058 , n11059 , n11060 , n11061 , n11062 ,
     n11063 , n11064 , n11065 , n11066 , n11067 , n11068 , n11069 , n11070 , n11071 , n11072 ,
     n11073 , n11074 , n11075 , n11076 , n11077 , n11078 , n11079 , n11080 , n11081 , n11082 ,
     n11083 , n11084 , n11085 , n11086 , n11087 , n11088 , n11089 , n11090 , n11091 , n11092 ,
     n11093 , n11094 , n11095 , n11096 , n11097 , n11098 , n11099 , n11100 , n11101 , n11102 ,
     n11103 , n11104 , n11105 , n11106 , n11107 , n11108 , n11109 , n11110 , n11111 , n11112 ,
     n11113 , n11114 , n11115 , n11116 , n11117 , n11118 , n11119 , n11120 , n11121 , n11122 ,
     n11123 , n11124 , n11125 , n11126 , n11127 , n11128 , n11129 , n11130 , n11131 , n11132 ,
     n11133 , n11134 , n11135 , n11136 , n11137 , n11138 , n11139 , n11140 , n11141 , n11142 ,
     n11143 , n11144 , n11145 , n11146 , n11147 , n11148 , n11149 , n11150 , n11151 , n11152 ,
     n11153 , n11154 , n11155 , n11156 , n11157 , n11158 , n11159 , n11160 , n11161 , n11162 ,
     n11163 , n11164 , n11165 , n11166 , n11167 , n11168 , n11169 , n11170 , n11171 , n11172 ,
     n11173 , n11174 , n11175 , n11176 , n11177 , n11178 , n11179 , n11180 , n11181 , n11182 ,
     n11183 , n11184 , n11185 , n11186 , n11187 , n11188 , n11189 , n11190 , n11191 , n11192 ,
     n11193 , n11194 , n11195 , n11196 , n11197 , n11198 , n11199 , n11200 , n11201 , n11202 ,
     n11203 , n11204 , n11205 , n11206 , n11207 , n11208 , n11209 , n11210 , n11211 , n11212 ,
     n11213 , n11214 , n11215 , n11216 , n11217 , n11218 , n11219 , n11220 , n11221 , n11222 ,
     n11223 , n11224 , n11225 , n11226 , n11227 , n11228 , n11229 , n11230 , n11231 , n11232 ,
     n11233 , n11234 , n11235 , n11236 , n11237 , n11238 , n11239 , n11240 , n11241 , n11242 ,
     n11243 , n11244 , n11245 , n11246 , n11247 , n11248 , n11249 , n11250 , n11251 , n11252 ,
     n11253 , n11254 , n11255 , n11256 , n11257 , n11258 , n11259 , n11260 , n11261 , n11262 ,
     n11263 , n11264 , n11265 , n11266 , n11267 , n11268 , n11269 , n11270 , n11271 , n11272 ,
     n11273 , n11274 , n11275 , n11276 , n11277 , n11278 , n11279 , n11280 , n11281 , n11282 ,
     n11283 , n11284 , n11285 , n11286 , n11287 , n11288 , n11289 , n11290 , n11291 , n11292 ,
     n11293 , n11294 , n11295 , n11296 , n11297 , n11298 , n11299 , n11300 , n11301 , n11302 ,
     n11303 , n11304 , n11305 , n11306 , n11307 , n11308 , n11309 , n11310 , n11311 , n11312 ,
     n11313 , n11314 , n11315 , n11316 , n11317 , n11318 , n11319 , n11320 , n11321 , n11322 ,
     n11323 , n11324 , n11325 , n11326 , n11327 , n11328 , n11329 , n11330 , n11331 , n11332 ,
     n11333 , n11334 , n11335 , n11336 , n11337 , n11338 , n11339 , n11340 , n11341 , n11342 ,
     n11343 , n11344 , n11345 , n11346 , n11347 , n11348 , n11349 , n11350 , n11351 , n11352 ,
     n11353 , n11354 , n11355 , n11356 , n11357 , n11358 , n11359 , n11360 , n11361 , n11362 ,
     n11363 , n11364 , n11365 , n11366 , n11367 , n11368 , n11369 , n11370 , n11371 , n11372 ,
     n11373 , n11374 , n11375 , n11376 , n11377 , n11378 , n11379 , n11380 , n11381 , n11382 ,
     n11383 , n11384 , n11385 , n11386 , n11387 , n11388 , n11389 , n11390 , n11391 , n11392 ,
     n11393 , n11394 , n11395 , n11396 , n11397 , n11398 , n11399 , n11400 , n11401 , n11402 ,
     n11403 , n11404 , n11405 , n11406 , n11407 , n11408 , n11409 , n11410 , n11411 , n11412 ,
     n11413 , n11414 , n11415 , n11416 , n11417 , n11418 , n11419 , n11420 , n11421 , n11422 ,
     n11423 , n11424 , n11425 , n11426 , n11427 , n11428 , n11429 , n11430 , n11431 , n11432 ,
     n11433 , n11434 , n11435 , n11436 , n11437 , n11438 , n11439 , n11440 , n11441 , n11442 ,
     n11443 , n11444 , n11445 , n11446 , n11447 , n11448 , n11449 , n11450 , n11451 , n11452 ,
     n11453 , n11454 , n11455 , n11456 , n11457 , n11458 , n11459 , n11460 , n11461 , n11462 ,
     n11463 , n11464 , n11465 , n11466 , n11467 , n11468 , n11469 , n11470 , n11471 , n11472 ,
     n11473 , n11474 , n11475 , n11476 , n11477 , n11478 , n11479 , n11480 , n11481 , n11482 ,
     n11483 , n11484 , n11485 , n11486 , n11487 , n11488 , n11489 , n11490 , n11491 , n11492 ,
     n11493 , n11494 , n11495 , n11496 , n11497 , n11498 , n11499 , n11500 , n11501 , n11502 ,
     n11503 , n11504 , n11505 , n11506 , n11507 , n11508 , n11509 , n11510 , n11511 , n11512 ,
     n11513 , n11514 , n11515 , n11516 , n11517 , n11518 , n11519 , n11520 , n11521 , n11522 ,
     n11523 , n11524 , n11525 , n11526 , n11527 , n11528 , n11529 , n11530 , n11531 , n11532 ,
     n11533 , n11534 , n11535 , n11536 , n11537 , n11538 , n11539 , n11540 , n11541 , n11542 ,
     n11543 , n11544 , n11545 , n11546 , n11547 , n11548 , n11549 , n11550 , n11551 , n11552 ,
     n11553 , n11554 , n11555 , n11556 , n11557 , n11558 , n11559 , n11560 , n11561 , n11562 ,
     n11563 , n11564 , n11565 , n11566 , n11567 , n11568 , n11569 , n11570 , n11571 , n11572 ,
     n11573 , n11574 , n11575 , n11576 , n11577 , n11578 , n11579 , n11580 , n11581 , n11582 ,
     n11583 , n11584 , n11585 , n11586 , n11587 , n11588 , n11589 , n11590 , n11591 , n11592 ,
     n11593 , n11594 , n11595 , n11596 , n11597 , n11598 , n11599 , n11600 , n11601 , n11602 ,
     n11603 , n11604 , n11605 , n11606 , n11607 , n11608 , n11609 , n11610 , n11611 , n11612 ,
     n11613 , n11614 , n11615 , n11616 , n11617 , n11618 , n11619 , n11620 , n11621 , n11622 ,
     n11623 , n11624 , n11625 , n11626 , n11627 , n11628 , n11629 , n11630 , n11631 , n11632 ,
     n11633 , n11634 , n11635 , n11636 , n11637 , n11638 , n11639 , n11640 , n11641 , n11642 ,
     n11643 , n11644 , n11645 , n11646 , n11647 , n11648 , n11649 , n11650 , n11651 , n11652 ,
     n11653 , n11654 , n11655 , n11656 , n11657 , n11658 , n11659 , n11660 , n11661 , n11662 ,
     n11663 , n11664 , n11665 , n11666 , n11667 , n11668 , n11669 , n11670 , n11671 , n11672 ,
     n11673 , n11674 , n11675 , n11676 , n11677 , n11678 , n11679 , n11680 , n11681 , n11682 ,
     n11683 , n11684 , n11685 , n11686 , n11687 , n11688 , n11689 , n11690 , n11691 , n11692 ,
     n11693 , n11694 , n11695 , n11696 , n11697 , n11698 , n11699 , n11700 , n11701 , n11702 ,
     n11703 , n11704 , n11705 , n11706 , n11707 , n11708 , n11709 , n11710 , n11711 , n11712 ,
     n11713 , n11714 , n11715 , n11716 , n11717 , n11718 , n11719 , n11720 , n11721 , n11722 ,
     n11723 , n11724 , n11725 , n11726 , n11727 , n11728 , n11729 , n11730 , n11731 , n11732 ,
     n11733 , n11734 , n11735 , n11736 , n11737 , n11738 , n11739 , n11740 , n11741 , n11742 ,
     n11743 , n11744 , n11745 , n11746 , n11747 , n11748 , n11749 , n11750 , n11751 , n11752 ,
     n11753 , n11754 , n11755 , n11756 , n11757 , n11758 , n11759 , n11760 , n11761 , n11762 ,
     n11763 , n11764 , n11765 , n11766 , n11767 , n11768 , n11769 , n11770 , n11771 , n11772 ,
     n11773 , n11774 , n11775 , n11776 , n11777 , n11778 , n11779 , n11780 , n11781 , n11782 ,
     n11783 , n11784 , n11785 , n11786 , n11787 , n11788 , n11789 , n11790 , n11791 , n11792 ,
     n11793 , n11794 , n11795 , n11796 , n11797 , n11798 , n11799 , n11800 , n11801 , n11802 ,
     n11803 , n11804 , n11805 , n11806 , n11807 , n11808 , n11809 , n11810 , n11811 , n11812 ,
     n11813 , n11814 , n11815 , n11816 , n11817 , n11818 , n11819 , n11820 , n11821 , n11822 ,
     n11823 , n11824 , n11825 , n11826 , n11827 , n11828 , n11829 , n11830 , n11831 , n11832 ,
     n11833 , n11834 , n11835 , n11836 , n11837 , n11838 , n11839 , n11840 , n11841 , n11842 ,
     n11843 , n11844 , n11845 , n11846 , n11847 , n11848 , n11849 , n11850 , n11851 , n11852 ,
     n11853 , n11854 , n11855 , n11856 , n11857 , n11858 , n11859 , n11860 , n11861 , n11862 ,
     n11863 , n11864 , n11865 , n11866 , n11867 , n11868 , n11869 , n11870 , n11871 , n11872 ,
     n11873 , n11874 , n11875 , n11876 , n11877 , n11878 , n11879 , n11880 , n11881 , n11882 ,
     n11883 , n11884 , n11885 , n11886 , n11887 , n11888 , n11889 , n11890 , n11891 , n11892 ,
     n11893 , n11894 , n11895 , n11896 , n11897 , n11898 , n11899 , n11900 , n11901 , n11902 ,
     n11903 , n11904 , n11905 , n11906 , n11907 , n11908 , n11909 , n11910 , n11911 , n11912 ,
     n11913 , n11914 , n11915 , n11916 , n11917 , n11918 , n11919 , n11920 , n11921 , n11922 ,
     n11923 , n11924 , n11925 , n11926 , n11927 , n11928 , n11929 , n11930 , n11931 , n11932 ,
     n11933 , n11934 , n11935 , n11936 , n11937 , n11938 , n11939 , n11940 , n11941 , n11942 ,
     n11943 , n11944 , n11945 , n11946 , n11947 , n11948 , n11949 , n11950 , n11951 , n11952 ,
     n11953 , n11954 , n11955 , n11956 , n11957 , n11958 , n11959 , n11960 , n11961 , n11962 ,
     n11963 , n11964 , n11965 , n11966 , n11967 , n11968 , n11969 , n11970 , n11971 , n11972 ,
     n11973 , n11974 , n11975 , n11976 , n11977 , n11978 , n11979 , n11980 , n11981 , n11982 ,
     n11983 , n11984 , n11985 , n11986 , n11987 , n11988 , n11989 , n11990 , n11991 , n11992 ,
     n11993 , n11994 , n11995 , n11996 , n11997 , n11998 , n11999 , n12000 , n12001 , n12002 ,
     n12003 , n12004 , n12005 , n12006 , n12007 , n12008 , n12009 , n12010 , n12011 , n12012 ,
     n12013 , n12014 , n12015 , n12016 , n12017 , n12018 , n12019 , n12020 , n12021 , n12022 ,
     n12023 , n12024 , n12025 , n12026 , n12027 , n12028 , n12029 , n12030 , n12031 , n12032 ,
     n12033 , n12034 , n12035 , n12036 , n12037 , n12038 , n12039 , n12040 , n12041 , n12042 ,
     n12043 , n12044 , n12045 , n12046 , n12047 , n12048 , n12049 , n12050 , n12051 , n12052 ,
     n12053 , n12054 , n12055 , n12056 , n12057 , n12058 , n12059 , n12060 , n12061 , n12062 ,
     n12063 , n12064 , n12065 , n12066 , n12067 , n12068 , n12069 , n12070 , n12071 , n12072 ,
     n12073 , n12074 , n12075 , n12076 , n12077 , n12078 , n12079 , n12080 , n12081 , n12082 ,
     n12083 , n12084 , n12085 , n12086 , n12087 , n12088 , n12089 , n12090 , n12091 , n12092 ,
     n12093 , n12094 , n12095 , n12096 , n12097 , n12098 , n12099 , n12100 , n12101 , n12102 ,
     n12103 , n12104 , n12105 , n12106 , n12107 , n12108 , n12109 , n12110 , n12111 , n12112 ,
     n12113 , n12114 , n12115 , n12116 , n12117 , n12118 , n12119 , n12120 , n12121 , n12122 ,
     n12123 , n12124 , n12125 , n12126 , n12127 , n12128 , n12129 , n12130 , n12131 , n12132 ,
     n12133 , n12134 , n12135 , n12136 , n12137 , n12138 , n12139 , n12140 , n12141 , n12142 ,
     n12143 , n12144 , n12145 , n12146 , n12147 , n12148 , n12149 , n12150 , n12151 , n12152 ,
     n12153 , n12154 , n12155 , n12156 , n12157 , n12158 , n12159 , n12160 , n12161 , n12162 ,
     n12163 , n12164 , n12165 , n12166 , n12167 , n12168 , n12169 , n12170 , n12171 , n12172 ,
     n12173 , n12174 , n12175 , n12176 , n12177 , n12178 , n12179 , n12180 , n12181 , n12182 ,
     n12183 , n12184 , n12185 , n12186 , n12187 , n12188 , n12189 , n12190 , n12191 , n12192 ,
     n12193 , n12194 , n12195 , n12196 , n12197 , n12198 , n12199 , n12200 , n12201 , n12202 ,
     n12203 , n12204 , n12205 , n12206 , n12207 , n12208 , n12209 , n12210 , n12211 , n12212 ,
     n12213 , n12214 , n12215 , n12216 , n12217 , n12218 , n12219 , n12220 , n12221 , n12222 ,
     n12223 , n12224 , n12225 , n12226 , n12227 , n12228 , n12229 , n12230 , n12231 , n12232 ,
     n12233 , n12234 , n12235 , n12236 , n12237 , n12238 , n12239 , n12240 , n12241 , n12242 ,
     n12243 , n12244 , n12245 , n12246 , n12247 , n12248 , n12249 , n12250 , n12251 , n12252 ,
     n12253 , n12254 , n12255 , n12256 , n12257 , n12258 , n12259 , n12260 , n12261 , n12262 ,
     n12263 , n12264 , n12265 , n12266 , n12267 , n12268 , n12269 , n12270 , n12271 , n12272 ,
     n12273 , n12274 , n12275 , n12276 , n12277 , n12278 , n12279 , n12280 , n12281 , n12282 ,
     n12283 , n12284 , n12285 , n12286 , n12287 , n12288 , n12289 , n12290 , n12291 , n12292 ,
     n12293 , n12294 , n12295 , n12296 , n12297 , n12298 , n12299 , n12300 , n12301 , n12302 ,
     n12303 , n12304 , n12305 , n12306 , n12307 , n12308 , n12309 , n12310 , n12311 , n12312 ,
     n12313 , n12314 , n12315 , n12316 , n12317 , n12318 , n12319 , n12320 , n12321 , n12322 ,
     n12323 , n12324 , n12325 , n12326 , n12327 , n12328 , n12329 , n12330 , n12331 , n12332 ,
     n12333 , n12334 , n12335 , n12336 , n12337 , n12338 , n12339 , n12340 , n12341 , n12342 ,
     n12343 , n12344 , n12345 , n12346 , n12347 , n12348 , n12349 , n12350 , n12351 , n12352 ,
     n12353 , n12354 , n12355 , n12356 , n12357 , n12358 , n12359 , n12360 , n12361 , n12362 ,
     n12363 , n12364 , n12365 , n12366 , n12367 , n12368 , n12369 , n12370 , n12371 , n12372 ,
     n12373 , n12374 , n12375 , n12376 , n12377 , n12378 , n12379 , n12380 , n12381 , n12382 ,
     n12383 , n12384 , n12385 , n12386 , n12387 , n12388 , n12389 , n12390 , n12391 , n12392 ,
     n12393 , n12394 , n12395 , n12396 , n12397 , n12398 , n12399 , n12400 , n12401 , n12402 ,
     n12403 , n12404 , n12405 , n12406 , n12407 , n12408 , n12409 , n12410 , n12411 , n12412 ,
     n12413 , n12414 , n12415 , n12416 , n12417 , n12418 , n12419 , n12420 , n12421 , n12422 ,
     n12423 , n12424 , n12425 , n12426 , n12427 , n12428 , n12429 , n12430 , n12431 , n12432 ,
     n12433 , n12434 , n12435 , n12436 , n12437 , n12438 , n12439 , n12440 , n12441 , n12442 ,
     n12443 , n12444 , n12445 , n12446 , n12447 , n12448 , n12449 , n12450 , n12451 , n12452 ,
     n12453 , n12454 , n12455 , n12456 , n12457 , n12458 , n12459 , n12460 , n12461 , n12462 ,
     n12463 , n12464 , n12465 , n12466 , n12467 , n12468 , n12469 , n12470 , n12471 , n12472 ,
     n12473 , n12474 , n12475 , n12476 , n12477 , n12478 , n12479 , n12480 , n12481 , n12482 ,
     n12483 , n12484 , n12485 , n12486 , n12487 , n12488 , n12489 , n12490 , n12491 , n12492 ,
     n12493 , n12494 , n12495 , n12496 , n12497 , n12498 , n12499 , n12500 , n12501 , n12502 ,
     n12503 , n12504 , n12505 , n12506 , n12507 , n12508 , n12509 , n12510 , n12511 , n12512 ,
     n12513 , n12514 , n12515 , n12516 , n12517 , n12518 , n12519 , n12520 , n12521 , n12522 ,
     n12523 , n12524 , n12525 , n12526 , n12527 , n12528 , n12529 , n12530 , n12531 , n12532 ,
     n12533 , n12534 , n12535 , n12536 , n12537 , n12538 , n12539 , n12540 , n12541 , n12542 ,
     n12543 , n12544 , n12545 , n12546 , n12547 , n12548 , n12549 , n12550 , n12551 , n12552 ,
     n12553 , n12554 , n12555 , n12556 , n12557 , n12558 , n12559 , n12560 , n12561 , n12562 ,
     n12563 , n12564 , n12565 , n12566 , n12567 , n12568 , n12569 , n12570 , n12571 , n12572 ,
     n12573 , n12574 , n12575 , n12576 , n12577 , n12578 , n12579 , n12580 , n12581 , n12582 ,
     n12583 , n12584 , n12585 , n12586 , n12587 , n12588 , n12589 , n12590 , n12591 , n12592 ,
     n12593 , n12594 , n12595 , n12596 , n12597 , n12598 , n12599 , n12600 , n12601 , n12602 ,
     n12603 , n12604 , n12605 , n12606 , n12607 , n12608 , n12609 , n12610 , n12611 , n12612 ,
     n12613 , n12614 , n12615 , n12616 , n12617 , n12618 , n12619 , n12620 , n12621 , n12622 ,
     n12623 , n12624 , n12625 , n12626 , n12627 , n12628 , n12629 , n12630 , n12631 , n12632 ,
     n12633 , n12634 , n12635 , n12636 , n12637 , n12638 , n12639 , n12640 , n12641 , n12642 ,
     n12643 , n12644 , n12645 , n12646 , n12647 , n12648 , n12649 , n12650 , n12651 , n12652 ,
     n12653 , n12654 , n12655 , n12656 , n12657 , n12658 , n12659 , n12660 , n12661 , n12662 ,
     n12663 , n12664 , n12665 , n12666 , n12667 , n12668 , n12669 , n12670 , n12671 , n12672 ,
     n12673 , n12674 , n12675 , n12676 , n12677 , n12678 , n12679 , n12680 , n12681 , n12682 ,
     n12683 , n12684 , n12685 , n12686 , n12687 , n12688 , n12689 , n12690 , n12691 , n12692 ,
     n12693 , n12694 , n12695 , n12696 , n12697 , n12698 , n12699 , n12700 , n12701 , n12702 ,
     n12703 , n12704 , n12705 , n12706 , n12707 , n12708 , n12709 , n12710 , n12711 , n12712 ,
     n12713 , n12714 , n12715 , n12716 , n12717 , n12718 , n12719 , n12720 , n12721 , n12722 ,
     n12723 , n12724 , n12725 , n12726 , n12727 , n12728 , n12729 , n12730 , n12731 , n12732 ,
     n12733 , n12734 , n12735 , n12736 , n12737 , n12738 , n12739 , n12740 , n12741 , n12742 ,
     n12743 , n12744 , n12745 , n12746 , n12747 , n12748 , n12749 , n12750 , n12751 , n12752 ,
     n12753 , n12754 , n12755 , n12756 , n12757 , n12758 , n12759 , n12760 , n12761 , n12762 ,
     n12763 , n12764 , n12765 , n12766 , n12767 , n12768 , n12769 , n12770 , n12771 , n12772 ,
     n12773 , n12774 , n12775 , n12776 , n12777 , n12778 , n12779 , n12780 , n12781 , n12782 ,
     n12783 , n12784 , n12785 , n12786 , n12787 , n12788 , n12789 , n12790 , n12791 , n12792 ,
     n12793 , n12794 , n12795 , n12796 , n12797 , n12798 , n12799 , n12800 , n12801 , n12802 ,
     n12803 , n12804 , n12805 , n12806 , n12807 , n12808 , n12809 , n12810 , n12811 , n12812 ,
     n12813 , n12814 , n12815 , n12816 , n12817 , n12818 , n12819 , n12820 , n12821 , n12822 ,
     n12823 , n12824 , n12825 , n12826 , n12827 , n12828 , n12829 , n12830 , n12831 , n12832 ,
     n12833 , n12834 , n12835 , n12836 , n12837 , n12838 , n12839 , n12840 , n12841 , n12842 ,
     n12843 , n12844 , n12845 , n12846 , n12847 , n12848 , n12849 , n12850 , n12851 , n12852 ,
     n12853 , n12854 , n12855 , n12856 , n12857 , n12858 , n12859 , n12860 , n12861 , n12862 ,
     n12863 , n12864 , n12865 , n12866 , n12867 , n12868 , n12869 , n12870 , n12871 , n12872 ,
     n12873 , n12874 , n12875 , n12876 , n12877 , n12878 , n12879 , n12880 , n12881 , n12882 ,
     n12883 , n12884 , n12885 , n12886 , n12887 , n12888 , n12889 , n12890 , n12891 , n12892 ,
     n12893 , n12894 , n12895 , n12896 , n12897 , n12898 , n12899 , n12900 , n12901 , n12902 ,
     n12903 , n12904 , n12905 , n12906 , n12907 , n12908 , n12909 , n12910 , n12911 , n12912 ,
     n12913 , n12914 , n12915 , n12916 , n12917 , n12918 , n12919 , n12920 , n12921 , n12922 ,
     n12923 , n12924 , n12925 , n12926 , n12927 , n12928 , n12929 , n12930 , n12931 , n12932 ,
     n12933 , n12934 , n12935 , n12936 , n12937 , n12938 , n12939 , n12940 , n12941 , n12942 ,
     n12943 , n12944 , n12945 , n12946 , n12947 , n12948 , n12949 , n12950 , n12951 , n12952 ,
     n12953 , n12954 , n12955 , n12956 , n12957 , n12958 , n12959 , n12960 , n12961 , n12962 ,
     n12963 , n12964 , n12965 , n12966 , n12967 , n12968 , n12969 , n12970 , n12971 , n12972 ,
     n12973 , n12974 , n12975 , n12976 , n12977 , n12978 , n12979 , n12980 , n12981 , n12982 ,
     n12983 , n12984 , n12985 , n12986 , n12987 , n12988 , n12989 , n12990 , n12991 , n12992 ,
     n12993 , n12994 , n12995 , n12996 , n12997 , n12998 , n12999 , n13000 , n13001 , n13002 ,
     n13003 , n13004 , n13005 , n13006 , n13007 , n13008 , n13009 , n13010 , n13011 , n13012 ,
     n13013 , n13014 , n13015 , n13016 , n13017 , n13018 , n13019 , n13020 , n13021 , n13022 ,
     n13023 , n13024 , n13025 , n13026 , n13027 , n13028 , n13029 , n13030 , n13031 , n13032 ,
     n13033 , n13034 , n13035 , n13036 , n13037 , n13038 , n13039 , n13040 , n13041 , n13042 ,
     n13043 , n13044 , n13045 , n13046 , n13047 , n13048 , n13049 , n13050 , n13051 , n13052 ,
     n13053 , n13054 , n13055 , n13056 , n13057 , n13058 , n13059 , n13060 , n13061 , n13062 ,
     n13063 , n13064 , n13065 , n13066 , n13067 , n13068 , n13069 , n13070 , n13071 , n13072 ,
     n13073 , n13074 , n13075 , n13076 , n13077 , n13078 , n13079 , n13080 , n13081 , n13082 ,
     n13083 , n13084 , n13085 , n13086 , n13087 , n13088 , n13089 , n13090 , n13091 , n13092 ,
     n13093 , n13094 , n13095 , n13096 , n13097 , n13098 , n13099 , n13100 , n13101 , n13102 ,
     n13103 , n13104 , n13105 , n13106 , n13107 , n13108 , n13109 , n13110 , n13111 , n13112 ,
     n13113 , n13114 , n13115 , n13116 , n13117 , n13118 , n13119 , n13120 , n13121 , n13122 ,
     n13123 , n13124 , n13125 , n13126 , n13127 , n13128 , n13129 , n13130 , n13131 , n13132 ,
     n13133 , n13134 , n13135 , n13136 , n13137 , n13138 , n13139 , n13140 , n13141 , n13142 ,
     n13143 , n13144 , n13145 , n13146 , n13147 , n13148 , n13149 , n13150 , n13151 , n13152 ,
     n13153 , n13154 , n13155 , n13156 , n13157 , n13158 , n13159 , n13160 , n13161 , n13162 ,
     n13163 , n13164 , n13165 , n13166 , n13167 , n13168 , n13169 , n13170 , n13171 , n13172 ,
     n13173 , n13174 , n13175 , n13176 , n13177 , n13178 , n13179 , n13180 , n13181 , n13182 ,
     n13183 , n13184 , n13185 , n13186 , n13187 , n13188 , n13189 , n13190 , n13191 , n13192 ,
     n13193 , n13194 , n13195 , n13196 , n13197 , n13198 , n13199 , n13200 , n13201 , n13202 ,
     n13203 , n13204 , n13205 , n13206 , n13207 , n13208 , n13209 , n13210 , n13211 , n13212 ,
     n13213 , n13214 , n13215 , n13216 , n13217 , n13218 , n13219 , n13220 , n13221 , n13222 ,
     n13223 , n13224 , n13225 , n13226 , n13227 , n13228 , n13229 , n13230 , n13231 , n13232 ,
     n13233 , n13234 , n13235 , n13236 , n13237 , n13238 , n13239 , n13240 , n13241 , n13242 ,
     n13243 , n13244 , n13245 , n13246 , n13247 , n13248 , n13249 , n13250 , n13251 , n13252 ,
     n13253 , n13254 , n13255 , n13256 , n13257 , n13258 , n13259 , n13260 , n13261 , n13262 ,
     n13263 , n13264 , n13265 , n13266 , n13267 , n13268 , n13269 , n13270 , n13271 , n13272 ,
     n13273 , n13274 , n13275 , n13276 , n13277 , n13278 , n13279 , n13280 , n13281 , n13282 ,
     n13283 , n13284 , n13285 , n13286 , n13287 , n13288 , n13289 , n13290 , n13291 , n13292 ,
     n13293 , n13294 , n13295 , n13296 , n13297 , n13298 , n13299 , n13300 , n13301 , n13302 ,
     n13303 , n13304 , n13305 , n13306 , n13307 , n13308 , n13309 , n13310 , n13311 , n13312 ,
     n13313 , n13314 , n13315 , n13316 , n13317 , n13318 , n13319 , n13320 , n13321 , n13322 ,
     n13323 , n13324 , n13325 , n13326 , n13327 , n13328 , n13329 , n13330 , n13331 , n13332 ,
     n13333 , n13334 , n13335 , n13336 , n13337 , n13338 , n13339 , n13340 , n13341 , n13342 ,
     n13343 , n13344 , n13345 , n13346 , n13347 , n13348 , n13349 , n13350 , n13351 , n13352 ,
     n13353 , n13354 , n13355 , n13356 , n13357 , n13358 , n13359 , n13360 , n13361 , n13362 ,
     n13363 , n13364 , n13365 , n13366 , n13367 , n13368 , n13369 , n13370 , n13371 , n13372 ,
     n13373 , n13374 , n13375 , n13376 , n13377 , n13378 , n13379 , n13380 , n13381 , n13382 ,
     n13383 , n13384 , n13385 , n13386 , n13387 , n13388 , n13389 , n13390 , n13391 , n13392 ,
     n13393 , n13394 , n13395 , n13396 , n13397 , n13398 , n13399 , n13400 , n13401 , n13402 ,
     n13403 , n13404 , n13405 , n13406 , n13407 , n13408 , n13409 , n13410 , n13411 , n13412 ,
     n13413 , n13414 , n13415 , n13416 , n13417 , n13418 , n13419 , n13420 , n13421 , n13422 ,
     n13423 , n13424 , n13425 , n13426 , n13427 , n13428 , n13429 , n13430 , n13431 , n13432 ,
     n13433 , n13434 , n13435 , n13436 , n13437 , n13438 , n13439 , n13440 , n13441 , n13442 ,
     n13443 , n13444 , n13445 , n13446 , n13447 , n13448 , n13449 , n13450 , n13451 , n13452 ,
     n13453 , n13454 , n13455 , n13456 , n13457 , n13458 , n13459 , n13460 , n13461 , n13462 ,
     n13463 , n13464 , n13465 , n13466 , n13467 , n13468 , n13469 , n13470 , n13471 , n13472 ,
     n13473 , n13474 , n13475 , n13476 , n13477 , n13478 , n13479 , n13480 , n13481 , n13482 ,
     n13483 , n13484 , n13485 , n13486 , n13487 , n13488 , n13489 , n13490 , n13491 , n13492 ,
     n13493 , n13494 , n13495 , n13496 , n13497 , n13498 , n13499 , n13500 , n13501 , n13502 ,
     n13503 , n13504 , n13505 , n13506 , n13507 , n13508 , n13509 , n13510 , n13511 , n13512 ,
     n13513 , n13514 , n13515 , n13516 , n13517 , n13518 , n13519 , n13520 , n13521 , n13522 ,
     n13523 , n13524 , n13525 , n13526 , n13527 , n13528 , n13529 , n13530 , n13531 , n13532 ,
     n13533 , n13534 , n13535 , n13536 , n13537 , n13538 , n13539 , n13540 , n13541 , n13542 ,
     n13543 , n13544 , n13545 , n13546 , n13547 , n13548 , n13549 , n13550 , n13551 , n13552 ,
     n13553 , n13554 , n13555 , n13556 , n13557 , n13558 , n13559 , n13560 , n13561 , n13562 ,
     n13563 , n13564 , n13565 , n13566 , n13567 , n13568 , n13569 , n13570 , n13571 , n13572 ,
     n13573 , n13574 , n13575 , n13576 , n13577 , n13578 , n13579 , n13580 , n13581 , n13582 ,
     n13583 , n13584 , n13585 , n13586 , n13587 , n13588 , n13589 , n13590 , n13591 , n13592 ,
     n13593 , n13594 , n13595 , n13596 , n13597 , n13598 , n13599 , n13600 , n13601 , n13602 ,
     n13603 , n13604 , n13605 , n13606 , n13607 , n13608 , n13609 , n13610 , n13611 , n13612 ,
     n13613 , n13614 , n13615 , n13616 , n13617 , n13618 , n13619 , n13620 , n13621 , n13622 ,
     n13623 , n13624 , n13625 , n13626 , n13627 , n13628 , n13629 , n13630 , n13631 , n13632 ,
     n13633 , n13634 , n13635 , n13636 , n13637 , n13638 , n13639 , n13640 , n13641 , n13642 ,
     n13643 , n13644 , n13645 , n13646 , n13647 , n13648 , n13649 , n13650 , n13651 , n13652 ,
     n13653 , n13654 , n13655 , n13656 , n13657 , n13658 , n13659 , n13660 , n13661 , n13662 ,
     n13663 , n13664 , n13665 , n13666 , n13667 , n13668 , n13669 , n13670 , n13671 , n13672 ,
     n13673 , n13674 , n13675 , n13676 , n13677 , n13678 , n13679 , n13680 , n13681 , n13682 ,
     n13683 , n13684 , n13685 , n13686 , n13687 , n13688 , n13689 , n13690 , n13691 , n13692 ,
     n13693 , n13694 , n13695 , n13696 , n13697 , n13698 , n13699 , n13700 , n13701 , n13702 ,
     n13703 , n13704 , n13705 , n13706 , n13707 , n13708 , n13709 , n13710 , n13711 , n13712 ,
     n13713 , n13714 , n13715 , n13716 , n13717 , n13718 , n13719 , n13720 , n13721 , n13722 ,
     n13723 , n13724 , n13725 , n13726 , n13727 , n13728 , n13729 , n13730 , n13731 , n13732 ,
     n13733 , n13734 , n13735 , n13736 , n13737 , n13738 , n13739 , n13740 , n13741 , n13742 ,
     n13743 , n13744 , n13745 , n13746 , n13747 , n13748 , n13749 , n13750 , n13751 , n13752 ,
     n13753 , n13754 , n13755 , n13756 , n13757 , n13758 , n13759 , n13760 , n13761 , n13762 ,
     n13763 , n13764 , n13765 , n13766 , n13767 , n13768 , n13769 , n13770 , n13771 , n13772 ,
     n13773 , n13774 , n13775 , n13776 , n13777 , n13778 , n13779 , n13780 , n13781 , n13782 ,
     n13783 , n13784 , n13785 , n13786 , n13787 , n13788 , n13789 , n13790 , n13791 , n13792 ,
     n13793 , n13794 , n13795 , n13796 , n13797 , n13798 , n13799 , n13800 , n13801 , n13802 ,
     n13803 , n13804 , n13805 , n13806 , n13807 , n13808 , n13809 , n13810 , n13811 , n13812 ,
     n13813 , n13814 , n13815 , n13816 , n13817 , n13818 , n13819 , n13820 , n13821 , n13822 ,
     n13823 , n13824 , n13825 , n13826 , n13827 , n13828 , n13829 , n13830 , n13831 , n13832 ,
     n13833 , n13834 , n13835 , n13836 , n13837 , n13838 , n13839 , n13840 , n13841 , n13842 ,
     n13843 , n13844 , n13845 , n13846 , n13847 , n13848 , n13849 , n13850 , n13851 , n13852 ,
     n13853 , n13854 , n13855 , n13856 , n13857 , n13858 , n13859 , n13860 , n13861 , n13862 ,
     n13863 , n13864 , n13865 , n13866 , n13867 , n13868 , n13869 , n13870 , n13871 , n13872 ,
     n13873 , n13874 , n13875 , n13876 , n13877 , n13878 , n13879 , n13880 , n13881 , n13882 ,
     n13883 , n13884 , n13885 , n13886 , n13887 , n13888 , n13889 , n13890 , n13891 , n13892 ,
     n13893 , n13894 , n13895 , n13896 , n13897 , n13898 , n13899 , n13900 , n13901 , n13902 ,
     n13903 , n13904 , n13905 , n13906 , n13907 , n13908 , n13909 , n13910 , n13911 , n13912 ,
     n13913 , n13914 , n13915 , n13916 , n13917 , n13918 , n13919 , n13920 , n13921 , n13922 ,
     n13923 , n13924 , n13925 , n13926 , n13927 , n13928 , n13929 , n13930 , n13931 , n13932 ,
     n13933 , n13934 , n13935 , n13936 , n13937 , n13938 , n13939 , n13940 , n13941 , n13942 ,
     n13943 , n13944 , n13945 , n13946 , n13947 , n13948 , n13949 , n13950 , n13951 , n13952 ,
     n13953 , n13954 , n13955 , n13956 , n13957 , n13958 , n13959 , n13960 , n13961 , n13962 ,
     n13963 , n13964 , n13965 , n13966 , n13967 , n13968 , n13969 , n13970 , n13971 , n13972 ,
     n13973 , n13974 , n13975 , n13976 , n13977 , n13978 , n13979 , n13980 , n13981 , n13982 ,
     n13983 , n13984 , n13985 , n13986 , n13987 , n13988 , n13989 , n13990 , n13991 , n13992 ,
     n13993 , n13994 , n13995 , n13996 , n13997 , n13998 , n13999 , n14000 , n14001 , n14002 ,
     n14003 , n14004 , n14005 , n14006 , n14007 , n14008 , n14009 , n14010 , n14011 , n14012 ,
     n14013 , n14014 , n14015 , n14016 , n14017 , n14018 , n14019 , n14020 , n14021 , n14022 ,
     n14023 , n14024 , n14025 , n14026 , n14027 , n14028 , n14029 , n14030 , n14031 , n14032 ,
     n14033 , n14034 , n14035 , n14036 , n14037 , n14038 , n14039 , n14040 , n14041 , n14042 ,
     n14043 , n14044 , n14045 , n14046 , n14047 , n14048 , n14049 , n14050 , n14051 , n14052 ,
     n14053 , n14054 , n14055 , n14056 , n14057 , n14058 , n14059 , n14060 , n14061 , n14062 ,
     n14063 , n14064 , n14065 , n14066 , n14067 , n14068 , n14069 , n14070 , n14071 , n14072 ,
     n14073 , n14074 , n14075 , n14076 , n14077 , n14078 , n14079 , n14080 , n14081 , n14082 ,
     n14083 , n14084 , n14085 , n14086 , n14087 , n14088 , n14089 , n14090 , n14091 , n14092 ,
     n14093 , n14094 , n14095 , n14096 , n14097 , n14098 , n14099 , n14100 , n14101 , n14102 ,
     n14103 , n14104 , n14105 , n14106 , n14107 , n14108 , n14109 , n14110 , n14111 , n14112 ,
     n14113 , n14114 , n14115 , n14116 , n14117 , n14118 , n14119 , n14120 , n14121 , n14122 ,
     n14123 , n14124 , n14125 , n14126 , n14127 , n14128 , n14129 , n14130 , n14131 , n14132 ,
     n14133 , n14134 , n14135 , n14136 , n14137 , n14138 , n14139 , n14140 , n14141 , n14142 ,
     n14143 , n14144 , n14145 , n14146 , n14147 , n14148 , n14149 , n14150 , n14151 , n14152 ,
     n14153 , n14154 , n14155 , n14156 , n14157 , n14158 , n14159 , n14160 , n14161 , n14162 ,
     n14163 , n14164 , n14165 , n14166 , n14167 , n14168 , n14169 , n14170 , n14171 , n14172 ,
     n14173 , n14174 , n14175 , n14176 , n14177 , n14178 , n14179 , n14180 , n14181 , n14182 ,
     n14183 , n14184 , n14185 , n14186 , n14187 , n14188 , n14189 , n14190 , n14191 , n14192 ,
     n14193 , n14194 , n14195 , n14196 , n14197 , n14198 , n14199 , n14200 , n14201 , n14202 ,
     n14203 , n14204 , n14205 , n14206 , n14207 , n14208 , n14209 , n14210 , n14211 , n14212 ,
     n14213 , n14214 , n14215 , n14216 , n14217 , n14218 , n14219 , n14220 , n14221 , n14222 ,
     n14223 , n14224 , n14225 , n14226 , n14227 , n14228 , n14229 , n14230 , n14231 , n14232 ,
     n14233 , n14234 , n14235 , n14236 , n14237 , n14238 , n14239 , n14240 , n14241 , n14242 ,
     n14243 , n14244 , n14245 , n14246 , n14247 , n14248 , n14249 , n14250 , n14251 , n14252 ,
     n14253 , n14254 , n14255 , n14256 , n14257 , n14258 , n14259 , n14260 , n14261 , n14262 ,
     n14263 , n14264 , n14265 , n14266 , n14267 , n14268 , n14269 , n14270 , n14271 , n14272 ,
     n14273 , n14274 , n14275 , n14276 , n14277 , n14278 , n14279 , n14280 , n14281 , n14282 ,
     n14283 , n14284 , n14285 , n14286 , n14287 , n14288 , n14289 , n14290 , n14291 , n14292 ,
     n14293 , n14294 , n14295 , n14296 , n14297 , n14298 , n14299 , n14300 , n14301 , n14302 ,
     n14303 , n14304 , n14305 , n14306 , n14307 , n14308 , n14309 , n14310 , n14311 , n14312 ,
     n14313 , n14314 , n14315 , n14316 , n14317 , n14318 , n14319 , n14320 , n14321 , n14322 ,
     n14323 , n14324 , n14325 , n14326 , n14327 , n14328 , n14329 , n14330 , n14331 , n14332 ,
     n14333 , n14334 , n14335 , n14336 , n14337 , n14338 , n14339 , n14340 , n14341 , n14342 ,
     n14343 , n14344 , n14345 , n14346 , n14347 , n14348 , n14349 , n14350 , n14351 , n14352 ,
     n14353 , n14354 , n14355 , n14356 , n14357 , n14358 , n14359 , n14360 , n14361 , n14362 ,
     n14363 , n14364 , n14365 , n14366 , n14367 , n14368 , n14369 , n14370 , n14371 , n14372 ,
     n14373 , n14374 , n14375 , n14376 , n14377 , n14378 , n14379 , n14380 , n14381 , n14382 ,
     n14383 , n14384 , n14385 , n14386 , n14387 , n14388 , n14389 , n14390 , n14391 , n14392 ,
     n14393 , n14394 , n14395 , n14396 , n14397 , n14398 , n14399 , n14400 , n14401 , n14402 ,
     n14403 , n14404 , n14405 , n14406 , n14407 , n14408 , n14409 , n14410 , n14411 , n14412 ,
     n14413 , n14414 , n14415 , n14416 , n14417 , n14418 , n14419 , n14420 , n14421 , n14422 ,
     n14423 , n14424 , n14425 , n14426 , n14427 , n14428 , n14429 , n14430 , n14431 , n14432 ,
     n14433 , n14434 , n14435 , n14436 , n14437 , n14438 , n14439 , n14440 , n14441 , n14442 ,
     n14443 , n14444 , n14445 , n14446 , n14447 , n14448 , n14449 , n14450 , n14451 , n14452 ,
     n14453 , n14454 , n14455 , n14456 , n14457 , n14458 , n14459 , n14460 , n14461 , n14462 ,
     n14463 , n14464 , n14465 , n14466 , n14467 , n14468 , n14469 , n14470 , n14471 , n14472 ,
     n14473 , n14474 , n14475 , n14476 , n14477 , n14478 , n14479 , n14480 , n14481 , n14482 ,
     n14483 , n14484 , n14485 , n14486 , n14487 , n14488 , n14489 , n14490 , n14491 , n14492 ,
     n14493 , n14494 , n14495 , n14496 , n14497 , n14498 , n14499 , n14500 , n14501 , n14502 ,
     n14503 , n14504 , n14505 , n14506 , n14507 , n14508 , n14509 , n14510 , n14511 , n14512 ,
     n14513 , n14514 , n14515 , n14516 , n14517 , n14518 , n14519 , n14520 , n14521 , n14522 ,
     n14523 , n14524 , n14525 , n14526 , n14527 , n14528 , n14529 , n14530 , n14531 , n14532 ,
     n14533 , n14534 , n14535 , n14536 , n14537 , n14538 , n14539 , n14540 , n14541 , n14542 ,
     n14543 , n14544 , n14545 , n14546 , n14547 , n14548 , n14549 , n14550 , n14551 , n14552 ,
     n14553 , n14554 , n14555 , n14556 , n14557 , n14558 , n14559 , n14560 , n14561 , n14562 ,
     n14563 , n14564 , n14565 , n14566 , n14567 , n14568 , n14569 , n14570 , n14571 , n14572 ,
     n14573 , n14574 , n14575 , n14576 , n14577 , n14578 , n14579 , n14580 , n14581 , n14582 ,
     n14583 , n14584 , n14585 , n14586 , n14587 , n14588 , n14589 , n14590 , n14591 , n14592 ,
     n14593 , n14594 , n14595 , n14596 , n14597 , n14598 , n14599 , n14600 , n14601 , n14602 ,
     n14603 , n14604 , n14605 , n14606 , n14607 , n14608 , n14609 , n14610 , n14611 , n14612 ,
     n14613 , n14614 , n14615 , n14616 , n14617 , n14618 , n14619 , n14620 , n14621 , n14622 ,
     n14623 , n14624 , n14625 , n14626 , n14627 , n14628 , n14629 , n14630 , n14631 , n14632 ,
     n14633 , n14634 , n14635 , n14636 , n14637 , n14638 , n14639 , n14640 , n14641 , n14642 ,
     n14643 , n14644 , n14645 , n14646 , n14647 , n14648 , n14649 , n14650 , n14651 , n14652 ,
     n14653 , n14654 , n14655 , n14656 , n14657 , n14658 , n14659 , n14660 , n14661 , n14662 ,
     n14663 , n14664 , n14665 , n14666 , n14667 , n14668 , n14669 , n14670 , n14671 , n14672 ,
     n14673 , n14674 , n14675 , n14676 , n14677 , n14678 , n14679 , n14680 , n14681 , n14682 ,
     n14683 , n14684 , n14685 , n14686 , n14687 , n14688 , n14689 , n14690 , n14691 , n14692 ,
     n14693 , n14694 , n14695 , n14696 , n14697 , n14698 , n14699 , n14700 , n14701 , n14702 ,
     n14703 , n14704 , n14705 , n14706 , n14707 , n14708 , n14709 , n14710 , n14711 , n14712 ,
     n14713 , n14714 , n14715 , n14716 , n14717 , n14718 , n14719 , n14720 , n14721 , n14722 ,
     n14723 , n14724 , n14725 , n14726 , n14727 , n14728 , n14729 , n14730 , n14731 , n14732 ,
     n14733 , n14734 , n14735 , n14736 , n14737 , n14738 , n14739 , n14740 , n14741 , n14742 ,
     n14743 , n14744 , n14745 , n14746 , n14747 , n14748 , n14749 , n14750 , n14751 , n14752 ,
     n14753 , n14754 , n14755 , n14756 , n14757 , n14758 , n14759 , n14760 , n14761 , n14762 ,
     n14763 , n14764 , n14765 , n14766 , n14767 , n14768 , n14769 , n14770 , n14771 , n14772 ,
     n14773 , n14774 , n14775 , n14776 , n14777 , n14778 , n14779 , n14780 , n14781 , n14782 ,
     n14783 , n14784 , n14785 , n14786 , n14787 , n14788 , n14789 , n14790 , n14791 , n14792 ,
     n14793 , n14794 , n14795 , n14796 , n14797 , n14798 , n14799 , n14800 , n14801 , n14802 ,
     n14803 , n14804 , n14805 , n14806 , n14807 , n14808 , n14809 , n14810 , n14811 , n14812 ,
     n14813 , n14814 , n14815 , n14816 , n14817 , n14818 , n14819 , n14820 , n14821 , n14822 ,
     n14823 , n14824 , n14825 , n14826 , n14827 , n14828 , n14829 , n14830 , n14831 , n14832 ,
     n14833 , n14834 , n14835 , n14836 , n14837 , n14838 , n14839 , n14840 , n14841 , n14842 ,
     n14843 , n14844 , n14845 , n14846 , n14847 , n14848 , n14849 , n14850 , n14851 , n14852 ,
     n14853 , n14854 , n14855 , n14856 , n14857 , n14858 , n14859 , n14860 , n14861 , n14862 ,
     n14863 , n14864 , n14865 , n14866 , n14867 , n14868 , n14869 , n14870 , n14871 , n14872 ,
     n14873 , n14874 , n14875 , n14876 , n14877 , n14878 , n14879 , n14880 , n14881 , n14882 ,
     n14883 , n14884 , n14885 , n14886 , n14887 , n14888 , n14889 , n14890 , n14891 , n14892 ,
     n14893 , n14894 , n14895 , n14896 , n14897 , n14898 , n14899 , n14900 , n14901 , n14902 ,
     n14903 , n14904 , n14905 , n14906 , n14907 , n14908 , n14909 , n14910 , n14911 , n14912 ,
     n14913 , n14914 , n14915 , n14916 , n14917 , n14918 , n14919 , n14920 , n14921 , n14922 ,
     n14923 , n14924 , n14925 , n14926 , n14927 , n14928 , n14929 , n14930 , n14931 , n14932 ,
     n14933 , n14934 , n14935 , n14936 , n14937 , n14938 , n14939 , n14940 , n14941 , n14942 ,
     n14943 , n14944 , n14945 , n14946 , n14947 , n14948 , n14949 , n14950 , n14951 , n14952 ,
     n14953 , n14954 , n14955 , n14956 , n14957 , n14958 , n14959 , n14960 , n14961 , n14962 ,
     n14963 , n14964 , n14965 , n14966 , n14967 , n14968 , n14969 , n14970 , n14971 , n14972 ,
     n14973 , n14974 , n14975 , n14976 , n14977 , n14978 , n14979 , n14980 , n14981 , n14982 ,
     n14983 , n14984 , n14985 , n14986 , n14987 , n14988 , n14989 , n14990 , n14991 , n14992 ,
     n14993 , n14994 , n14995 , n14996 , n14997 , n14998 , n14999 , n15000 , n15001 , n15002 ,
     n15003 , n15004 , n15005 , n15006 , n15007 , n15008 , n15009 , n15010 , n15011 , n15012 ,
     n15013 , n15014 , n15015 , n15016 , n15017 , n15018 , n15019 , n15020 , n15021 , n15022 ,
     n15023 , n15024 , n15025 , n15026 , n15027 , n15028 , n15029 , n15030 , n15031 , n15032 ,
     n15033 , n15034 , n15035 , n15036 , n15037 , n15038 , n15039 , n15040 , n15041 , n15042 ,
     n15043 , n15044 , n15045 , n15046 , n15047 , n15048 , n15049 , n15050 , n15051 , n15052 ,
     n15053 , n15054 , n15055 , n15056 , n15057 , n15058 , n15059 , n15060 , n15061 , n15062 ,
     n15063 , n15064 , n15065 , n15066 , n15067 , n15068 , n15069 , n15070 , n15071 , n15072 ,
     n15073 , n15074 , n15075 , n15076 , n15077 , n15078 , n15079 , n15080 , n15081 , n15082 ,
     n15083 , n15084 , n15085 , n15086 , n15087 , n15088 , n15089 , n15090 , n15091 , n15092 ,
     n15093 , n15094 , n15095 , n15096 , n15097 , n15098 , n15099 , n15100 , n15101 , n15102 ,
     n15103 , n15104 , n15105 , n15106 , n15107 , n15108 , n15109 , n15110 , n15111 , n15112 ,
     n15113 , n15114 , n15115 , n15116 , n15117 , n15118 , n15119 , n15120 , n15121 , n15122 ,
     n15123 , n15124 , n15125 , n15126 , n15127 , n15128 , n15129 , n15130 , n15131 , n15132 ,
     n15133 , n15134 , n15135 , n15136 , n15137 , n15138 , n15139 , n15140 , n15141 , n15142 ,
     n15143 , n15144 , n15145 , n15146 , n15147 , n15148 , n15149 , n15150 , n15151 , n15152 ,
     n15153 , n15154 , n15155 , n15156 , n15157 , n15158 , n15159 , n15160 , n15161 , n15162 ,
     n15163 , n15164 , n15165 , n15166 , n15167 , n15168 , n15169 , n15170 , n15171 , n15172 ,
     n15173 , n15174 , n15175 , n15176 , n15177 , n15178 , n15179 , n15180 , n15181 , n15182 ,
     n15183 , n15184 , n15185 , n15186 , n15187 , n15188 , n15189 , n15190 , n15191 , n15192 ,
     n15193 , n15194 , n15195 , n15196 , n15197 , n15198 , n15199 , n15200 , n15201 , n15202 ,
     n15203 , n15204 , n15205 , n15206 , n15207 , n15208 , n15209 , n15210 , n15211 , n15212 ,
     n15213 , n15214 , n15215 , n15216 , n15217 , n15218 , n15219 , n15220 , n15221 , n15222 ,
     n15223 , n15224 , n15225 , n15226 , n15227 , n15228 , n15229 , n15230 , n15231 , n15232 ,
     n15233 , n15234 , n15235 , n15236 , n15237 , n15238 , n15239 , n15240 , n15241 , n15242 ,
     n15243 , n15244 , n15245 , n15246 , n15247 , n15248 , n15249 , n15250 , n15251 , n15252 ,
     n15253 , n15254 , n15255 , n15256 , n15257 , n15258 , n15259 , n15260 , n15261 , n15262 ,
     n15263 , n15264 , n15265 , n15266 , n15267 , n15268 , n15269 , n15270 , n15271 , n15272 ,
     n15273 , n15274 , n15275 , n15276 , n15277 , n15278 , n15279 , n15280 , n15281 , n15282 ,
     n15283 , n15284 , n15285 , n15286 , n15287 , n15288 , n15289 , n15290 , n15291 , n15292 ,
     n15293 , n15294 , n15295 , n15296 , n15297 , n15298 , n15299 , n15300 , n15301 , n15302 ,
     n15303 , n15304 , n15305 , n15306 , n15307 , n15308 , n15309 , n15310 , n15311 , n15312 ,
     n15313 , n15314 , n15315 , n15316 , n15317 , n15318 , n15319 , n15320 , n15321 , n15322 ,
     n15323 , n15324 , n15325 , n15326 , n15327 , n15328 , n15329 , n15330 , n15331 , n15332 ,
     n15333 , n15334 , n15335 , n15336 , n15337 , n15338 , n15339 , n15340 , n15341 , n15342 ,
     n15343 , n15344 , n15345 , n15346 , n15347 , n15348 , n15349 , n15350 , n15351 , n15352 ,
     n15353 , n15354 , n15355 , n15356 , n15357 , n15358 , n15359 , n15360 , n15361 , n15362 ,
     n15363 , n15364 , n15365 , n15366 , n15367 , n15368 , n15369 , n15370 , n15371 , n15372 ,
     n15373 , n15374 , n15375 , n15376 , n15377 , n15378 , n15379 , n15380 , n15381 , n15382 ,
     n15383 , n15384 , n15385 , n15386 , n15387 , n15388 , n15389 , n15390 , n15391 , n15392 ,
     n15393 , n15394 , n15395 , n15396 , n15397 , n15398 , n15399 , n15400 , n15401 , n15402 ,
     n15403 , n15404 , n15405 , n15406 , n15407 , n15408 , n15409 , n15410 , n15411 , n15412 ,
     n15413 , n15414 , n15415 , n15416 , n15417 , n15418 , n15419 , n15420 , n15421 , n15422 ,
     n15423 , n15424 , n15425 , n15426 , n15427 , n15428 , n15429 , n15430 , n15431 , n15432 ,
     n15433 , n15434 , n15435 , n15436 , n15437 , n15438 , n15439 , n15440 , n15441 , n15442 ,
     n15443 , n15444 , n15445 , n15446 , n15447 , n15448 , n15449 , n15450 , n15451 , n15452 ,
     n15453 , n15454 , n15455 , n15456 , n15457 , n15458 , n15459 , n15460 , n15461 , n15462 ,
     n15463 , n15464 , n15465 , n15466 , n15467 , n15468 , n15469 , n15470 , n15471 , n15472 ,
     n15473 , n15474 , n15475 , n15476 , n15477 , n15478 , n15479 , n15480 , n15481 , n15482 ,
     n15483 , n15484 , n15485 , n15486 , n15487 , n15488 , n15489 , n15490 , n15491 , n15492 ,
     n15493 , n15494 , n15495 , n15496 , n15497 , n15498 , n15499 , n15500 , n15501 , n15502 ,
     n15503 , n15504 , n15505 , n15506 , n15507 , n15508 , n15509 , n15510 , n15511 , n15512 ,
     n15513 , n15514 , n15515 , n15516 , n15517 , n15518 , n15519 , n15520 , n15521 , n15522 ,
     n15523 , n15524 , n15525 , n15526 , n15527 , n15528 , n15529 , n15530 , n15531 , n15532 ,
     n15533 , n15534 , n15535 , n15536 , n15537 , n15538 , n15539 , n15540 , n15541 , n15542 ,
     n15543 , n15544 , n15545 , n15546 , n15547 , n15548 , n15549 , n15550 , n15551 , n15552 ,
     n15553 , n15554 , n15555 , n15556 , n15557 , n15558 , n15559 , n15560 , n15561 , n15562 ,
     n15563 , n15564 , n15565 , n15566 , n15567 , n15568 , n15569 , n15570 , n15571 , n15572 ,
     n15573 , n15574 , n15575 , n15576 , n15577 , n15578 , n15579 , n15580 , n15581 , n15582 ,
     n15583 , n15584 , n15585 , n15586 , n15587 , n15588 , n15589 , n15590 , n15591 , n15592 ,
     n15593 , n15594 , n15595 , n15596 , n15597 , n15598 , n15599 , n15600 , n15601 , n15602 ,
     n15603 , n15604 , n15605 , n15606 , n15607 , n15608 , n15609 , n15610 , n15611 , n15612 ,
     n15613 , n15614 , n15615 , n15616 , n15617 , n15618 , n15619 , n15620 , n15621 , n15622 ,
     n15623 , n15624 , n15625 , n15626 , n15627 , n15628 , n15629 , n15630 , n15631 , n15632 ,
     n15633 , n15634 , n15635 , n15636 , n15637 , n15638 , n15639 , n15640 , n15641 , n15642 ,
     n15643 , n15644 , n15645 , n15646 , n15647 , n15648 , n15649 , n15650 , n15651 , n15652 ,
     n15653 , n15654 , n15655 , n15656 , n15657 , n15658 , n15659 , n15660 , n15661 , n15662 ,
     n15663 , n15664 , n15665 , n15666 , n15667 , n15668 , n15669 , n15670 , n15671 , n15672 ,
     n15673 , n15674 , n15675 , n15676 , n15677 , n15678 , n15679 , n15680 , n15681 , n15682 ,
     n15683 , n15684 , n15685 , n15686 , n15687 , n15688 , n15689 , n15690 , n15691 , n15692 ,
     n15693 , n15694 , n15695 , n15696 , n15697 , n15698 , n15699 , n15700 , n15701 , n15702 ,
     n15703 , n15704 , n15705 , n15706 , n15707 , n15708 , n15709 , n15710 , n15711 , n15712 ,
     n15713 , n15714 , n15715 , n15716 , n15717 , n15718 , n15719 , n15720 , n15721 , n15722 ,
     n15723 , n15724 , n15725 , n15726 , n15727 , n15728 , n15729 , n15730 , n15731 , n15732 ,
     n15733 , n15734 , n15735 , n15736 , n15737 , n15738 , n15739 , n15740 , n15741 , n15742 ,
     n15743 , n15744 , n15745 , n15746 , n15747 , n15748 , n15749 , n15750 , n15751 , n15752 ,
     n15753 , n15754 , n15755 , n15756 , n15757 , n15758 , n15759 , n15760 , n15761 , n15762 ,
     n15763 , n15764 , n15765 , n15766 , n15767 , n15768 , n15769 , n15770 , n15771 , n15772 ,
     n15773 , n15774 , n15775 , n15776 , n15777 , n15778 , n15779 , n15780 , n15781 , n15782 ,
     n15783 , n15784 , n15785 , n15786 , n15787 , n15788 , n15789 , n15790 , n15791 , n15792 ,
     n15793 , n15794 , n15795 , n15796 , n15797 , n15798 , n15799 , n15800 , n15801 , n15802 ,
     n15803 , n15804 , n15805 , n15806 , n15807 , n15808 , n15809 , n15810 , n15811 , n15812 ,
     n15813 , n15814 , n15815 , n15816 , n15817 , n15818 , n15819 , n15820 , n15821 , n15822 ,
     n15823 , n15824 , n15825 , n15826 , n15827 , n15828 , n15829 , n15830 , n15831 , n15832 ,
     n15833 , n15834 , n15835 , n15836 , n15837 , n15838 , n15839 , n15840 , n15841 , n15842 ,
     n15843 , n15844 , n15845 , n15846 , n15847 , n15848 , n15849 , n15850 , n15851 , n15852 ,
     n15853 , n15854 , n15855 , n15856 , n15857 , n15858 , n15859 , n15860 , n15861 , n15862 ,
     n15863 , n15864 , n15865 , n15866 , n15867 , n15868 , n15869 , n15870 , n15871 , n15872 ,
     n15873 , n15874 , n15875 , n15876 , n15877 , n15878 , n15879 , n15880 , n15881 , n15882 ,
     n15883 , n15884 , n15885 , n15886 , n15887 , n15888 , n15889 , n15890 , n15891 , n15892 ,
     n15893 , n15894 , n15895 , n15896 , n15897 , n15898 , n15899 , n15900 , n15901 , n15902 ,
     n15903 , n15904 , n15905 , n15906 , n15907 , n15908 , n15909 , n15910 , n15911 , n15912 ,
     n15913 , n15914 , n15915 , n15916 , n15917 , n15918 , n15919 , n15920 , n15921 , n15922 ,
     n15923 , n15924 , n15925 , n15926 , n15927 , n15928 , n15929 , n15930 , n15931 , n15932 ,
     n15933 , n15934 , n15935 , n15936 , n15937 , n15938 , n15939 , n15940 , n15941 , n15942 ,
     n15943 , n15944 , n15945 , n15946 , n15947 , n15948 , n15949 , n15950 , n15951 , n15952 ,
     n15953 , n15954 , n15955 , n15956 , n15957 , n15958 , n15959 , n15960 , n15961 , n15962 ,
     n15963 , n15964 , n15965 , n15966 , n15967 , n15968 , n15969 , n15970 , n15971 , n15972 ,
     n15973 , n15974 , n15975 , n15976 , n15977 , n15978 , n15979 , n15980 , n15981 , n15982 ,
     n15983 , n15984 , n15985 , n15986 , n15987 , n15988 , n15989 , n15990 , n15991 , n15992 ,
     n15993 , n15994 , n15995 , n15996 , n15997 , n15998 , n15999 , n16000 , n16001 , n16002 ,
     n16003 , n16004 , n16005 , n16006 , n16007 , n16008 , n16009 , n16010 , n16011 , n16012 ,
     n16013 , n16014 , n16015 , n16016 , n16017 , n16018 , n16019 , n16020 , n16021 , n16022 ,
     n16023 , n16024 , n16025 , n16026 , n16027 , n16028 , n16029 , n16030 , n16031 , n16032 ,
     n16033 , n16034 , n16035 , n16036 , n16037 , n16038 , n16039 , n16040 , n16041 , n16042 ,
     n16043 , n16044 , n16045 , n16046 , n16047 , n16048 , n16049 , n16050 , n16051 , n16052 ,
     n16053 , n16054 , n16055 , n16056 , n16057 , n16058 , n16059 , n16060 , n16061 , n16062 ,
     n16063 , n16064 , n16065 , n16066 , n16067 , n16068 , n16069 , n16070 , n16071 , n16072 ,
     n16073 , n16074 , n16075 , n16076 , n16077 , n16078 , n16079 , n16080 , n16081 , n16082 ,
     n16083 , n16084 , n16085 , n16086 , n16087 , n16088 , n16089 , n16090 , n16091 , n16092 ,
     n16093 , n16094 , n16095 , n16096 , n16097 , n16098 , n16099 , n16100 , n16101 , n16102 ,
     n16103 , n16104 , n16105 , n16106 , n16107 , n16108 , n16109 , n16110 , n16111 , n16112 ,
     n16113 , n16114 , n16115 , n16116 , n16117 , n16118 , n16119 , n16120 , n16121 , n16122 ,
     n16123 , n16124 , n16125 , n16126 , n16127 , n16128 , n16129 , n16130 , n16131 , n16132 ,
     n16133 , n16134 , n16135 , n16136 , n16137 , n16138 , n16139 , n16140 , n16141 , n16142 ,
     n16143 , n16144 , n16145 , n16146 , n16147 , n16148 , n16149 , n16150 , n16151 , n16152 ,
     n16153 , n16154 , n16155 , n16156 , n16157 , n16158 , n16159 , n16160 , n16161 , n16162 ,
     n16163 , n16164 , n16165 , n16166 , n16167 , n16168 , n16169 , n16170 , n16171 , n16172 ,
     n16173 , n16174 , n16175 , n16176 , n16177 , n16178 , n16179 , n16180 , n16181 , n16182 ,
     n16183 , n16184 , n16185 , n16186 , n16187 , n16188 , n16189 , n16190 , n16191 , n16192 ,
     n16193 , n16194 , n16195 , n16196 , n16197 , n16198 , n16199 , n16200 , n16201 , n16202 ,
     n16203 , n16204 , n16205 , n16206 , n16207 , n16208 , n16209 , n16210 , n16211 , n16212 ,
     n16213 , n16214 , n16215 , n16216 , n16217 , n16218 , n16219 , n16220 , n16221 , n16222 ,
     n16223 , n16224 , n16225 , n16226 , n16227 , n16228 , n16229 , n16230 , n16231 , n16232 ,
     n16233 , n16234 , n16235 , n16236 , n16237 , n16238 , n16239 , n16240 , n16241 , n16242 ,
     n16243 , n16244 , n16245 , n16246 , n16247 , n16248 , n16249 , n16250 , n16251 , n16252 ,
     n16253 , n16254 , n16255 , n16256 , n16257 , n16258 , n16259 , n16260 , n16261 , n16262 ,
     n16263 , n16264 , n16265 , n16266 , n16267 , n16268 , n16269 , n16270 , n16271 , n16272 ,
     n16273 , n16274 , n16275 , n16276 , n16277 , n16278 , n16279 , n16280 , n16281 , n16282 ,
     n16283 , n16284 , n16285 , n16286 , n16287 , n16288 , n16289 , n16290 , n16291 , n16292 ,
     n16293 , n16294 , n16295 , n16296 , n16297 , n16298 , n16299 , n16300 , n16301 , n16302 ,
     n16303 , n16304 , n16305 , n16306 , n16307 , n16308 , n16309 , n16310 , n16311 , n16312 ,
     n16313 , n16314 , n16315 , n16316 , n16317 , n16318 , n16319 , n16320 , n16321 , n16322 ,
     n16323 , n16324 , n16325 , n16326 , n16327 , n16328 , n16329 , n16330 , n16331 , n16332 ,
     n16333 , n16334 , n16335 , n16336 , n16337 , n16338 , n16339 , n16340 , n16341 , n16342 ,
     n16343 , n16344 , n16345 , n16346 , n16347 , n16348 , n16349 , n16350 , n16351 , n16352 ,
     n16353 , n16354 , n16355 , n16356 , n16357 , n16358 , n16359 , n16360 , n16361 , n16362 ,
     n16363 , n16364 , n16365 , n16366 , n16367 , n16368 , n16369 , n16370 , n16371 , n16372 ,
     n16373 , n16374 , n16375 , n16376 , n16377 , n16378 , n16379 , n16380 , n16381 , n16382 ,
     n16383 , n16384 , n16385 , n16386 , n16387 , n16388 , n16389 , n16390 , n16391 , n16392 ,
     n16393 , n16394 , n16395 , n16396 , n16397 , n16398 , n16399 , n16400 , n16401 , n16402 ,
     n16403 , n16404 , n16405 , n16406 , n16407 , n16408 , n16409 , n16410 , n16411 , n16412 ,
     n16413 , n16414 , n16415 , n16416 , n16417 , n16418 , n16419 , n16420 , n16421 , n16422 ,
     n16423 , n16424 , n16425 , n16426 , n16427 , n16428 , n16429 , n16430 , n16431 , n16432 ,
     n16433 , n16434 , n16435 , n16436 , n16437 , n16438 , n16439 , n16440 , n16441 , n16442 ,
     n16443 , n16444 , n16445 , n16446 , n16447 , n16448 , n16449 , n16450 , n16451 , n16452 ,
     n16453 , n16454 , n16455 , n16456 , n16457 , n16458 , n16459 , n16460 , n16461 , n16462 ,
     n16463 , n16464 , n16465 , n16466 , n16467 , n16468 , n16469 , n16470 , n16471 , n16472 ,
     n16473 , n16474 , n16475 , n16476 , n16477 , n16478 , n16479 , n16480 , n16481 , n16482 ,
     n16483 , n16484 , n16485 , n16486 , n16487 , n16488 , n16489 , n16490 , n16491 , n16492 ,
     n16493 , n16494 , n16495 , n16496 , n16497 , n16498 , n16499 , n16500 , n16501 , n16502 ,
     n16503 , n16504 , n16505 , n16506 , n16507 , n16508 , n16509 , n16510 , n16511 , n16512 ,
     n16513 , n16514 , n16515 , n16516 , n16517 , n16518 , n16519 , n16520 , n16521 , n16522 ,
     n16523 , n16524 , n16525 , n16526 , n16527 , n16528 , n16529 , n16530 , n16531 , n16532 ,
     n16533 , n16534 , n16535 , n16536 , n16537 , n16538 , n16539 , n16540 , n16541 , n16542 ,
     n16543 , n16544 , n16545 , n16546 , n16547 , n16548 , n16549 , n16550 , n16551 , n16552 ,
     n16553 , n16554 , n16555 , n16556 , n16557 , n16558 , n16559 , n16560 , n16561 , n16562 ,
     n16563 , n16564 , n16565 , n16566 , n16567 , n16568 , n16569 , n16570 , n16571 , n16572 ,
     n16573 , n16574 , n16575 , n16576 , n16577 , n16578 , n16579 , n16580 , n16581 , n16582 ,
     n16583 , n16584 , n16585 , n16586 , n16587 , n16588 , n16589 , n16590 , n16591 , n16592 ,
     n16593 , n16594 , n16595 , n16596 , n16597 , n16598 , n16599 , n16600 , n16601 , n16602 ,
     n16603 , n16604 , n16605 , n16606 , n16607 , n16608 , n16609 , n16610 , n16611 , n16612 ,
     n16613 , n16614 , n16615 , n16616 , n16617 , n16618 , n16619 , n16620 , n16621 , n16622 ,
     n16623 , n16624 , n16625 , n16626 , n16627 , n16628 , n16629 , n16630 , n16631 , n16632 ,
     n16633 , n16634 , n16635 , n16636 , n16637 , n16638 , n16639 , n16640 , n16641 , n16642 ,
     n16643 , n16644 , n16645 , n16646 , n16647 , n16648 , n16649 , n16650 , n16651 , n16652 ,
     n16653 , n16654 , n16655 , n16656 , n16657 , n16658 , n16659 , n16660 , n16661 , n16662 ,
     n16663 , n16664 , n16665 , n16666 , n16667 , n16668 , n16669 , n16670 , n16671 , n16672 ,
     n16673 , n16674 , n16675 , n16676 , n16677 , n16678 , n16679 , n16680 , n16681 , n16682 ,
     n16683 , n16684 , n16685 , n16686 , n16687 , n16688 , n16689 , n16690 , n16691 , n16692 ,
     n16693 , n16694 , n16695 , n16696 , n16697 , n16698 , n16699 , n16700 , n16701 , n16702 ,
     n16703 , n16704 , n16705 , n16706 , n16707 , n16708 , n16709 , n16710 , n16711 , n16712 ,
     n16713 , n16714 , n16715 , n16716 , n16717 , n16718 , n16719 , n16720 , n16721 , n16722 ,
     n16723 , n16724 , n16725 , n16726 , n16727 , n16728 , n16729 , n16730 , n16731 , n16732 ,
     n16733 , n16734 , n16735 , n16736 , n16737 , n16738 , n16739 , n16740 , n16741 , n16742 ,
     n16743 , n16744 , n16745 , n16746 , n16747 , n16748 , n16749 , n16750 , n16751 , n16752 ,
     n16753 , n16754 , n16755 , n16756 , n16757 , n16758 , n16759 , n16760 , n16761 , n16762 ,
     n16763 , n16764 , n16765 , n16766 , n16767 , n16768 , n16769 , n16770 , n16771 , n16772 ,
     n16773 , n16774 , n16775 , n16776 , n16777 , n16778 , n16779 , n16780 , n16781 , n16782 ,
     n16783 , n16784 , n16785 , n16786 , n16787 , n16788 , n16789 , n16790 , n16791 , n16792 ,
     n16793 , n16794 , n16795 , n16796 , n16797 , n16798 , n16799 , n16800 , n16801 , n16802 ,
     n16803 , n16804 , n16805 , n16806 , n16807 , n16808 , n16809 , n16810 , n16811 , n16812 ,
     n16813 , n16814 , n16815 , n16816 , n16817 , n16818 , n16819 , n16820 , n16821 , n16822 ,
     n16823 , n16824 , n16825 , n16826 , n16827 , n16828 , n16829 , n16830 , n16831 , n16832 ,
     n16833 , n16834 , n16835 , n16836 , n16837 , n16838 , n16839 , n16840 , n16841 , n16842 ,
     n16843 , n16844 , n16845 , n16846 , n16847 , n16848 , n16849 , n16850 , n16851 , n16852 ,
     n16853 , n16854 , n16855 , n16856 , n16857 , n16858 , n16859 , n16860 , n16861 , n16862 ,
     n16863 , n16864 , n16865 , n16866 , n16867 , n16868 , n16869 , n16870 , n16871 , n16872 ,
     n16873 , n16874 , n16875 , n16876 , n16877 , n16878 , n16879 , n16880 , n16881 , n16882 ,
     n16883 , n16884 , n16885 , n16886 , n16887 , n16888 , n16889 , n16890 , n16891 , n16892 ,
     n16893 , n16894 , n16895 , n16896 , n16897 , n16898 , n16899 , n16900 , n16901 , n16902 ,
     n16903 , n16904 , n16905 , n16906 , n16907 , n16908 , n16909 , n16910 , n16911 , n16912 ,
     n16913 , n16914 , n16915 , n16916 , n16917 , n16918 , n16919 , n16920 , n16921 , n16922 ,
     n16923 , n16924 , n16925 , n16926 , n16927 , n16928 , n16929 , n16930 , n16931 , n16932 ,
     n16933 , n16934 , n16935 , n16936 , n16937 , n16938 , n16939 , n16940 , n16941 , n16942 ,
     n16943 , n16944 , n16945 , n16946 , n16947 , n16948 , n16949 , n16950 , n16951 , n16952 ,
     n16953 , n16954 , n16955 , n16956 , n16957 , n16958 , n16959 , n16960 , n16961 , n16962 ,
     n16963 , n16964 , n16965 , n16966 , n16967 , n16968 , n16969 , n16970 , n16971 , n16972 ,
     n16973 , n16974 , n16975 , n16976 , n16977 , n16978 , n16979 , n16980 , n16981 , n16982 ,
     n16983 , n16984 , n16985 , n16986 , n16987 , n16988 , n16989 , n16990 , n16991 , n16992 ,
     n16993 , n16994 , n16995 , n16996 , n16997 , n16998 , n16999 , n17000 , n17001 , n17002 ,
     n17003 , n17004 , n17005 , n17006 , n17007 , n17008 , n17009 , n17010 , n17011 , n17012 ,
     n17013 , n17014 , n17015 , n17016 , n17017 , n17018 , n17019 , n17020 , n17021 , n17022 ,
     n17023 , n17024 , n17025 , n17026 , n17027 , n17028 , n17029 , n17030 , n17031 , n17032 ,
     n17033 , n17034 , n17035 , n17036 , n17037 , n17038 , n17039 , n17040 , n17041 , n17042 ,
     n17043 , n17044 , n17045 , n17046 , n17047 , n17048 , n17049 , n17050 , n17051 , n17052 ,
     n17053 , n17054 , n17055 , n17056 , n17057 , n17058 , n17059 , n17060 , n17061 , n17062 ,
     n17063 , n17064 , n17065 , n17066 , n17067 , n17068 , n17069 , n17070 , n17071 , n17072 ,
     n17073 , n17074 , n17075 , n17076 , n17077 , n17078 , n17079 , n17080 , n17081 , n17082 ,
     n17083 , n17084 , n17085 , n17086 , n17087 , n17088 , n17089 , n17090 , n17091 , n17092 ,
     n17093 , n17094 , n17095 , n17096 , n17097 , n17098 , n17099 , n17100 , n17101 , n17102 ,
     n17103 , n17104 , n17105 , n17106 , n17107 , n17108 , n17109 , n17110 , n17111 , n17112 ,
     n17113 , n17114 , n17115 , n17116 , n17117 , n17118 , n17119 , n17120 , n17121 , n17122 ,
     n17123 , n17124 , n17125 , n17126 , n17127 , n17128 , n17129 , n17130 , n17131 , n17132 ,
     n17133 , n17134 , n17135 , n17136 , n17137 , n17138 , n17139 , n17140 , n17141 , n17142 ,
     n17143 , n17144 , n17145 , n17146 , n17147 , n17148 , n17149 , n17150 , n17151 , n17152 ,
     n17153 , n17154 , n17155 , n17156 , n17157 , n17158 , n17159 , n17160 , n17161 , n17162 ,
     n17163 , n17164 , n17165 , n17166 , n17167 , n17168 , n17169 , n17170 , n17171 , n17172 ,
     n17173 , n17174 , n17175 , n17176 , n17177 , n17178 , n17179 , n17180 , n17181 , n17182 ,
     n17183 , n17184 , n17185 , n17186 , n17187 , n17188 , n17189 , n17190 , n17191 , n17192 ,
     n17193 , n17194 , n17195 , n17196 , n17197 , n17198 , n17199 , n17200 , n17201 , n17202 ,
     n17203 , n17204 , n17205 , n17206 , n17207 , n17208 , n17209 , n17210 , n17211 , n17212 ,
     n17213 , n17214 , n17215 , n17216 , n17217 , n17218 , n17219 , n17220 , n17221 , n17222 ,
     n17223 , n17224 , n17225 , n17226 , n17227 , n17228 , n17229 , n17230 , n17231 , n17232 ,
     n17233 , n17234 , n17235 , n17236 , n17237 , n17238 , n17239 , n17240 , n17241 , n17242 ,
     n17243 , n17244 , n17245 , n17246 , n17247 , n17248 , n17249 , n17250 , n17251 , n17252 ,
     n17253 , n17254 , n17255 , n17256 , n17257 , n17258 , n17259 , n17260 , n17261 , n17262 ,
     n17263 , n17264 , n17265 , n17266 , n17267 , n17268 , n17269 , n17270 , n17271 , n17272 ,
     n17273 , n17274 , n17275 , n17276 , n17277 , n17278 , n17279 , n17280 , n17281 , n17282 ,
     n17283 , n17284 , n17285 , n17286 , n17287 , n17288 , n17289 , n17290 , n17291 , n17292 ,
     n17293 , n17294 , n17295 , n17296 , n17297 , n17298 , n17299 , n17300 , n17301 , n17302 ,
     n17303 , n17304 , n17305 , n17306 , n17307 , n17308 , n17309 , n17310 , n17311 , n17312 ,
     n17313 , n17314 , n17315 , n17316 , n17317 , n17318 , n17319 , n17320 , n17321 , n17322 ,
     n17323 , n17324 , n17325 , n17326 , n17327 , n17328 , n17329 , n17330 , n17331 , n17332 ,
     n17333 , n17334 , n17335 , n17336 , n17337 , n17338 , n17339 , n17340 , n17341 , n17342 ,
     n17343 , n17344 , n17345 , n17346 , n17347 , n17348 , n17349 , n17350 , n17351 , n17352 ,
     n17353 , n17354 , n17355 , n17356 , n17357 , n17358 , n17359 , n17360 , n17361 , n17362 ,
     n17363 , n17364 , n17365 , n17366 , n17367 , n17368 , n17369 , n17370 , n17371 , n17372 ,
     n17373 , n17374 , n17375 , n17376 , n17377 , n17378 , n17379 , n17380 , n17381 , n17382 ,
     n17383 , n17384 , n17385 , n17386 , n17387 , n17388 , n17389 , n17390 , n17391 , n17392 ,
     n17393 , n17394 , n17395 , n17396 , n17397 , n17398 , n17399 , n17400 , n17401 , n17402 ,
     n17403 , n17404 , n17405 , n17406 , n17407 , n17408 , n17409 , n17410 , n17411 , n17412 ,
     n17413 , n17414 , n17415 , n17416 , n17417 , n17418 , n17419 , n17420 , n17421 , n17422 ,
     n17423 , n17424 , n17425 , n17426 , n17427 , n17428 , n17429 , n17430 , n17431 , n17432 ,
     n17433 , n17434 , n17435 , n17436 , n17437 , n17438 , n17439 , n17440 , n17441 , n17442 ,
     n17443 , n17444 , n17445 , n17446 , n17447 , n17448 , n17449 , n17450 , n17451 , n17452 ,
     n17453 , n17454 , n17455 , n17456 , n17457 , n17458 , n17459 , n17460 , n17461 , n17462 ,
     n17463 , n17464 , n17465 , n17466 , n17467 , n17468 , n17469 , n17470 , n17471 , n17472 ,
     n17473 , n17474 , n17475 , n17476 , n17477 , n17478 , n17479 , n17480 , n17481 , n17482 ,
     n17483 , n17484 , n17485 , n17486 , n17487 , n17488 , n17489 , n17490 , n17491 , n17492 ,
     n17493 , n17494 , n17495 , n17496 , n17497 , n17498 , n17499 , n17500 , n17501 , n17502 ,
     n17503 , n17504 , n17505 , n17506 , n17507 , n17508 , n17509 , n17510 , n17511 , n17512 ,
     n17513 , n17514 , n17515 , n17516 , n17517 , n17518 , n17519 , n17520 , n17521 , n17522 ,
     n17523 , n17524 , n17525 , n17526 , n17527 , n17528 , n17529 , n17530 , n17531 , n17532 ,
     n17533 , n17534 , n17535 , n17536 , n17537 , n17538 , n17539 , n17540 , n17541 , n17542 ,
     n17543 , n17544 , n17545 , n17546 , n17547 , n17548 , n17549 , n17550 , n17551 , n17552 ,
     n17553 , n17554 , n17555 , n17556 , n17557 , n17558 , n17559 , n17560 , n17561 , n17562 ,
     n17563 , n17564 , n17565 , n17566 , n17567 , n17568 , n17569 , n17570 , n17571 , n17572 ,
     n17573 , n17574 , n17575 , n17576 , n17577 , n17578 , n17579 , n17580 , n17581 , n17582 ,
     n17583 , n17584 , n17585 , n17586 , n17587 , n17588 , n17589 , n17590 , n17591 , n17592 ,
     n17593 , n17594 , n17595 , n17596 , n17597 , n17598 , n17599 , n17600 , n17601 , n17602 ,
     n17603 , n17604 , n17605 , n17606 , n17607 , n17608 , n17609 , n17610 , n17611 , n17612 ,
     n17613 , n17614 , n17615 , n17616 , n17617 , n17618 , n17619 , n17620 , n17621 , n17622 ,
     n17623 , n17624 , n17625 , n17626 , n17627 , n17628 , n17629 , n17630 , n17631 , n17632 ,
     n17633 , n17634 , n17635 , n17636 , n17637 , n17638 , n17639 , n17640 , n17641 , n17642 ,
     n17643 , n17644 , n17645 , n17646 , n17647 , n17648 , n17649 , n17650 , n17651 , n17652 ,
     n17653 , n17654 , n17655 , n17656 , n17657 , n17658 , n17659 , n17660 , n17661 , n17662 ,
     n17663 , n17664 , n17665 , n17666 , n17667 , n17668 , n17669 , n17670 , n17671 , n17672 ,
     n17673 , n17674 , n17675 , n17676 , n17677 , n17678 , n17679 , n17680 , n17681 , n17682 ,
     n17683 , n17684 , n17685 , n17686 , n17687 , n17688 , n17689 , n17690 , n17691 , n17692 ,
     n17693 , n17694 , n17695 , n17696 , n17697 , n17698 , n17699 , n17700 , n17701 , n17702 ,
     n17703 , n17704 , n17705 , n17706 , n17707 , n17708 , n17709 , n17710 , n17711 , n17712 ,
     n17713 , n17714 , n17715 , n17716 , n17717 , n17718 , n17719 , n17720 , n17721 , n17722 ,
     n17723 , n17724 , n17725 , n17726 , n17727 , n17728 , n17729 , n17730 , n17731 , n17732 ,
     n17733 , n17734 , n17735 , n17736 , n17737 , n17738 , n17739 , n17740 , n17741 , n17742 ,
     n17743 , n17744 , n17745 , n17746 , n17747 , n17748 , n17749 , n17750 , n17751 , n17752 ,
     n17753 , n17754 , n17755 , n17756 , n17757 , n17758 , n17759 , n17760 , n17761 , n17762 ,
     n17763 , n17764 , n17765 , n17766 , n17767 , n17768 , n17769 , n17770 , n17771 , n17772 ,
     n17773 , n17774 , n17775 , n17776 , n17777 , n17778 , n17779 , n17780 , n17781 , n17782 ,
     n17783 , n17784 , n17785 , n17786 , n17787 , n17788 , n17789 , n17790 , n17791 , n17792 ,
     n17793 , n17794 , n17795 , n17796 , n17797 , n17798 , n17799 , n17800 , n17801 , n17802 ,
     n17803 , n17804 , n17805 , n17806 , n17807 , n17808 , n17809 , n17810 , n17811 , n17812 ,
     n17813 , n17814 , n17815 , n17816 , n17817 , n17818 , n17819 , n17820 , n17821 , n17822 ,
     n17823 , n17824 , n17825 , n17826 , n17827 , n17828 , n17829 , n17830 , n17831 , n17832 ,
     n17833 , n17834 , n17835 , n17836 , n17837 , n17838 , n17839 , n17840 , n17841 , n17842 ,
     n17843 , n17844 , n17845 , n17846 , n17847 , n17848 , n17849 , n17850 , n17851 , n17852 ,
     n17853 , n17854 , n17855 , n17856 , n17857 , n17858 , n17859 , n17860 , n17861 , n17862 ,
     n17863 , n17864 , n17865 , n17866 , n17867 , n17868 , n17869 , n17870 , n17871 , n17872 ,
     n17873 , n17874 , n17875 , n17876 , n17877 , n17878 , n17879 , n17880 , n17881 , n17882 ,
     n17883 , n17884 , n17885 , n17886 , n17887 , n17888 , n17889 , n17890 , n17891 , n17892 ,
     n17893 , n17894 , n17895 , n17896 , n17897 , n17898 , n17899 , n17900 , n17901 , n17902 ,
     n17903 , n17904 , n17905 , n17906 , n17907 , n17908 , n17909 , n17910 , n17911 , n17912 ,
     n17913 , n17914 , n17915 , n17916 , n17917 , n17918 , n17919 , n17920 , n17921 , n17922 ,
     n17923 , n17924 , n17925 , n17926 , n17927 , n17928 , n17929 , n17930 , n17931 , n17932 ,
     n17933 , n17934 , n17935 , n17936 , n17937 , n17938 , n17939 , n17940 , n17941 , n17942 ,
     n17943 , n17944 , n17945 , n17946 , n17947 , n17948 , n17949 , n17950 , n17951 , n17952 ,
     n17953 , n17954 , n17955 , n17956 , n17957 , n17958 , n17959 , n17960 , n17961 , n17962 ,
     n17963 , n17964 , n17965 , n17966 , n17967 , n17968 , n17969 , n17970 , n17971 , n17972 ,
     n17973 , n17974 , n17975 , n17976 , n17977 , n17978 , n17979 , n17980 , n17981 , n17982 ,
     n17983 , n17984 , n17985 , n17986 , n17987 , n17988 , n17989 , n17990 , n17991 , n17992 ,
     n17993 , n17994 , n17995 , n17996 , n17997 , n17998 , n17999 , n18000 , n18001 , n18002 ,
     n18003 , n18004 , n18005 , n18006 , n18007 , n18008 , n18009 , n18010 , n18011 , n18012 ,
     n18013 , n18014 , n18015 , n18016 , n18017 , n18018 , n18019 , n18020 , n18021 , n18022 ,
     n18023 , n18024 , n18025 , n18026 , n18027 , n18028 , n18029 , n18030 , n18031 , n18032 ,
     n18033 , n18034 , n18035 , n18036 , n18037 , n18038 , n18039 , n18040 , n18041 , n18042 ,
     n18043 , n18044 , n18045 , n18046 , n18047 , n18048 , n18049 , n18050 , n18051 , n18052 ,
     n18053 , n18054 , n18055 , n18056 , n18057 , n18058 , n18059 , n18060 , n18061 , n18062 ,
     n18063 , n18064 , n18065 , n18066 , n18067 , n18068 , n18069 , n18070 , n18071 , n18072 ,
     n18073 , n18074 , n18075 , n18076 , n18077 , n18078 , n18079 , n18080 , n18081 , n18082 ,
     n18083 , n18084 , n18085 , n18086 , n18087 , n18088 , n18089 , n18090 , n18091 , n18092 ,
     n18093 , n18094 , n18095 , n18096 , n18097 , n18098 , n18099 , n18100 , n18101 , n18102 ,
     n18103 , n18104 , n18105 , n18106 , n18107 , n18108 , n18109 , n18110 , n18111 , n18112 ,
     n18113 , n18114 , n18115 , n18116 , n18117 , n18118 , n18119 , n18120 , n18121 , n18122 ,
     n18123 , n18124 , n18125 , n18126 , n18127 , n18128 , n18129 , n18130 , n18131 , n18132 ,
     n18133 , n18134 , n18135 , n18136 , n18137 , n18138 , n18139 , n18140 , n18141 , n18142 ,
     n18143 , n18144 , n18145 , n18146 , n18147 , n18148 , n18149 , n18150 , n18151 , n18152 ,
     n18153 , n18154 , n18155 , n18156 , n18157 , n18158 , n18159 , n18160 , n18161 , n18162 ,
     n18163 , n18164 , n18165 , n18166 , n18167 , n18168 , n18169 , n18170 , n18171 , n18172 ,
     n18173 , n18174 , n18175 , n18176 , n18177 , n18178 , n18179 , n18180 , n18181 , n18182 ,
     n18183 , n18184 , n18185 , n18186 , n18187 , n18188 , n18189 , n18190 , n18191 , n18192 ,
     n18193 , n18194 , n18195 , n18196 , n18197 , n18198 , n18199 , n18200 , n18201 , n18202 ,
     n18203 , n18204 , n18205 , n18206 , n18207 , n18208 , n18209 , n18210 , n18211 , n18212 ,
     n18213 , n18214 , n18215 , n18216 , n18217 , n18218 , n18219 , n18220 , n18221 , n18222 ,
     n18223 , n18224 , n18225 , n18226 , n18227 , n18228 , n18229 , n18230 , n18231 , n18232 ,
     n18233 , n18234 , n18235 , n18236 , n18237 , n18238 , n18239 , n18240 , n18241 , n18242 ,
     n18243 , n18244 , n18245 , n18246 , n18247 , n18248 , n18249 , n18250 , n18251 , n18252 ,
     n18253 , n18254 , n18255 , n18256 , n18257 , n18258 , n18259 , n18260 , n18261 , n18262 ,
     n18263 , n18264 , n18265 , n18266 , n18267 , n18268 , n18269 , n18270 , n18271 , n18272 ,
     n18273 , n18274 , n18275 , n18276 , n18277 , n18278 , n18279 , n18280 , n18281 , n18282 ,
     n18283 , n18284 , n18285 , n18286 , n18287 , n18288 , n18289 , n18290 , n18291 , n18292 ,
     n18293 , n18294 , n18295 , n18296 , n18297 , n18298 , n18299 , n18300 , n18301 , n18302 ,
     n18303 , n18304 , n18305 , n18306 , n18307 , n18308 , n18309 , n18310 , n18311 , n18312 ,
     n18313 , n18314 , n18315 , n18316 , n18317 , n18318 , n18319 , n18320 , n18321 , n18322 ,
     n18323 , n18324 , n18325 , n18326 , n18327 , n18328 , n18329 , n18330 , n18331 , n18332 ,
     n18333 , n18334 , n18335 , n18336 , n18337 , n18338 , n18339 , n18340 , n18341 , n18342 ,
     n18343 , n18344 , n18345 , n18346 , n18347 , n18348 , n18349 , n18350 , n18351 , n18352 ,
     n18353 , n18354 , n18355 , n18356 , n18357 , n18358 , n18359 , n18360 , n18361 , n18362 ,
     n18363 , n18364 , n18365 , n18366 , n18367 , n18368 , n18369 , n18370 , n18371 , n18372 ,
     n18373 , n18374 , n18375 , n18376 , n18377 , n18378 , n18379 , n18380 , n18381 , n18382 ,
     n18383 , n18384 , n18385 , n18386 , n18387 , n18388 , n18389 , n18390 , n18391 , n18392 ,
     n18393 , n18394 , n18395 , n18396 , n18397 , n18398 , n18399 , n18400 , n18401 , n18402 ,
     n18403 , n18404 , n18405 , n18406 , n18407 , n18408 , n18409 , n18410 , n18411 , n18412 ,
     n18413 , n18414 , n18415 , n18416 , n18417 , n18418 , n18419 , n18420 , n18421 , n18422 ,
     n18423 , n18424 , n18425 , n18426 , n18427 , n18428 , n18429 , n18430 , n18431 , n18432 ,
     n18433 , n18434 , n18435 , n18436 , n18437 , n18438 , n18439 , n18440 , n18441 , n18442 ,
     n18443 , n18444 , n18445 , n18446 , n18447 , n18448 , n18449 , n18450 , n18451 , n18452 ,
     n18453 , n18454 , n18455 , n18456 , n18457 , n18458 , n18459 , n18460 , n18461 , n18462 ,
     n18463 , n18464 , n18465 , n18466 , n18467 , n18468 , n18469 , n18470 , n18471 , n18472 ,
     n18473 , n18474 , n18475 , n18476 , n18477 , n18478 , n18479 , n18480 , n18481 , n18482 ,
     n18483 , n18484 , n18485 , n18486 , n18487 , n18488 , n18489 , n18490 , n18491 , n18492 ,
     n18493 , n18494 , n18495 , n18496 , n18497 , n18498 , n18499 , n18500 , n18501 , n18502 ,
     n18503 , n18504 , n18505 , n18506 , n18507 , n18508 , n18509 , n18510 , n18511 , n18512 ,
     n18513 , n18514 , n18515 , n18516 , n18517 , n18518 , n18519 , n18520 , n18521 , n18522 ,
     n18523 , n18524 , n18525 , n18526 , n18527 , n18528 , n18529 , n18530 , n18531 , n18532 ,
     n18533 , n18534 , n18535 , n18536 , n18537 , n18538 , n18539 , n18540 , n18541 , n18542 ,
     n18543 , n18544 , n18545 , n18546 , n18547 , n18548 , n18549 , n18550 , n18551 , n18552 ,
     n18553 , n18554 , n18555 , n18556 , n18557 , n18558 , n18559 , n18560 , n18561 , n18562 ,
     n18563 , n18564 , n18565 , n18566 , n18567 , n18568 , n18569 , n18570 , n18571 , n18572 ,
     n18573 , n18574 , n18575 , n18576 , n18577 , n18578 , n18579 , n18580 , n18581 , n18582 ,
     n18583 , n18584 , n18585 , n18586 , n18587 , n18588 , n18589 , n18590 , n18591 , n18592 ,
     n18593 , n18594 , n18595 , n18596 , n18597 , n18598 , n18599 , n18600 , n18601 , n18602 ,
     n18603 , n18604 , n18605 , n18606 , n18607 , n18608 , n18609 , n18610 , n18611 , n18612 ,
     n18613 , n18614 , n18615 , n18616 , n18617 , n18618 , n18619 , n18620 , n18621 , n18622 ,
     n18623 , n18624 , n18625 , n18626 , n18627 , n18628 , n18629 , n18630 , n18631 , n18632 ,
     n18633 , n18634 , n18635 , n18636 , n18637 , n18638 , n18639 , n18640 , n18641 , n18642 ,
     n18643 , n18644 , n18645 , n18646 , n18647 , n18648 , n18649 , n18650 , n18651 , n18652 ,
     n18653 , n18654 , n18655 , n18656 , n18657 , n18658 , n18659 , n18660 , n18661 , n18662 ,
     n18663 , n18664 , n18665 , n18666 , n18667 , n18668 , n18669 , n18670 , n18671 , n18672 ,
     n18673 , n18674 , n18675 , n18676 , n18677 , n18678 , n18679 , n18680 , n18681 , n18682 ,
     n18683 , n18684 , n18685 , n18686 , n18687 , n18688 , n18689 , n18690 , n18691 , n18692 ,
     n18693 , n18694 , n18695 , n18696 , n18697 , n18698 , n18699 , n18700 , n18701 , n18702 ,
     n18703 , n18704 , n18705 , n18706 , n18707 , n18708 , n18709 , n18710 , n18711 , n18712 ,
     n18713 , n18714 , n18715 , n18716 , n18717 , n18718 , n18719 , n18720 , n18721 , n18722 ,
     n18723 , n18724 , n18725 , n18726 , n18727 , n18728 , n18729 , n18730 , n18731 , n18732 ,
     n18733 , n18734 , n18735 , n18736 , n18737 , n18738 , n18739 , n18740 , n18741 , n18742 ,
     n18743 , n18744 , n18745 , n18746 , n18747 , n18748 , n18749 , n18750 , n18751 , n18752 ,
     n18753 , n18754 , n18755 , n18756 , n18757 , n18758 , n18759 , n18760 , n18761 , n18762 ,
     n18763 , n18764 , n18765 , n18766 , n18767 , n18768 , n18769 , n18770 , n18771 , n18772 ,
     n18773 , n18774 , n18775 , n18776 , n18777 , n18778 , n18779 , n18780 , n18781 , n18782 ,
     n18783 , n18784 , n18785 , n18786 , n18787 , n18788 , n18789 , n18790 , n18791 , n18792 ,
     n18793 , n18794 , n18795 , n18796 , n18797 , n18798 , n18799 , n18800 , n18801 , n18802 ,
     n18803 , n18804 , n18805 , n18806 , n18807 , n18808 , n18809 , n18810 , n18811 , n18812 ,
     n18813 , n18814 , n18815 , n18816 , n18817 , n18818 , n18819 , n18820 , n18821 , n18822 ,
     n18823 , n18824 , n18825 , n18826 , n18827 , n18828 , n18829 , n18830 , n18831 , n18832 ,
     n18833 , n18834 , n18835 , n18836 , n18837 , n18838 , n18839 , n18840 , n18841 , n18842 ,
     n18843 , n18844 , n18845 , n18846 , n18847 , n18848 , n18849 , n18850 , n18851 , n18852 ,
     n18853 , n18854 , n18855 , n18856 , n18857 , n18858 , n18859 , n18860 , n18861 , n18862 ,
     n18863 , n18864 , n18865 , n18866 , n18867 , n18868 , n18869 , n18870 , n18871 , n18872 ,
     n18873 , n18874 , n18875 , n18876 , n18877 , n18878 , n18879 , n18880 , n18881 , n18882 ,
     n18883 , n18884 , n18885 , n18886 , n18887 , n18888 , n18889 , n18890 , n18891 , n18892 ,
     n18893 , n18894 , n18895 , n18896 , n18897 , n18898 , n18899 , n18900 , n18901 , n18902 ,
     n18903 , n18904 , n18905 , n18906 , n18907 , n18908 , n18909 , n18910 , n18911 , n18912 ,
     n18913 , n18914 , n18915 , n18916 , n18917 , n18918 , n18919 , n18920 , n18921 , n18922 ,
     n18923 , n18924 , n18925 , n18926 , n18927 , n18928 , n18929 , n18930 , n18931 , n18932 ,
     n18933 , n18934 , n18935 , n18936 , n18937 , n18938 , n18939 , n18940 , n18941 , n18942 ,
     n18943 , n18944 , n18945 , n18946 , n18947 , n18948 , n18949 , n18950 , n18951 , n18952 ,
     n18953 , n18954 , n18955 , n18956 , n18957 , n18958 , n18959 , n18960 , n18961 , n18962 ,
     n18963 , n18964 , n18965 , n18966 , n18967 , n18968 , n18969 , n18970 , n18971 , n18972 ,
     n18973 , n18974 , n18975 , n18976 , n18977 , n18978 , n18979 , n18980 , n18981 , n18982 ,
     n18983 , n18984 , n18985 , n18986 , n18987 , n18988 , n18989 , n18990 , n18991 , n18992 ,
     n18993 , n18994 , n18995 , n18996 , n18997 , n18998 , n18999 , n19000 , n19001 , n19002 ,
     n19003 , n19004 , n19005 , n19006 , n19007 , n19008 , n19009 , n19010 , n19011 , n19012 ,
     n19013 , n19014 , n19015 , n19016 , n19017 , n19018 , n19019 , n19020 , n19021 , n19022 ,
     n19023 , n19024 , n19025 , n19026 , n19027 , n19028 , n19029 , n19030 , n19031 , n19032 ,
     n19033 , n19034 , n19035 , n19036 , n19037 , n19038 , n19039 , n19040 , n19041 , n19042 ,
     n19043 , n19044 , n19045 , n19046 , n19047 , n19048 , n19049 , n19050 , n19051 , n19052 ,
     n19053 , n19054 , n19055 , n19056 , n19057 , n19058 , n19059 , n19060 , n19061 , n19062 ,
     n19063 , n19064 , n19065 , n19066 , n19067 , n19068 , n19069 , n19070 , n19071 , n19072 ,
     n19073 , n19074 , n19075 , n19076 , n19077 , n19078 , n19079 , n19080 , n19081 , n19082 ,
     n19083 , n19084 , n19085 , n19086 , n19087 , n19088 , n19089 , n19090 , n19091 , n19092 ,
     n19093 , n19094 , n19095 , n19096 , n19097 , n19098 , n19099 , n19100 , n19101 , n19102 ,
     n19103 , n19104 , n19105 , n19106 , n19107 , n19108 , n19109 , n19110 , n19111 , n19112 ,
     n19113 , n19114 , n19115 , n19116 , n19117 , n19118 , n19119 , n19120 , n19121 , n19122 ,
     n19123 , n19124 , n19125 , n19126 , n19127 , n19128 , n19129 , n19130 , n19131 , n19132 ,
     n19133 , n19134 , n19135 , n19136 , n19137 , n19138 , n19139 , n19140 , n19141 , n19142 ,
     n19143 , n19144 , n19145 , n19146 , n19147 , n19148 , n19149 , n19150 , n19151 , n19152 ,
     n19153 , n19154 , n19155 , n19156 , n19157 , n19158 , n19159 , n19160 , n19161 , n19162 ,
     n19163 , n19164 , n19165 , n19166 , n19167 , n19168 , n19169 , n19170 , n19171 , n19172 ,
     n19173 , n19174 , n19175 , n19176 , n19177 , n19178 , n19179 , n19180 , n19181 , n19182 ,
     n19183 , n19184 , n19185 , n19186 , n19187 , n19188 , n19189 , n19190 , n19191 , n19192 ,
     n19193 , n19194 , n19195 , n19196 , n19197 , n19198 , n19199 , n19200 , n19201 , n19202 ,
     n19203 , n19204 , n19205 , n19206 , n19207 , n19208 , n19209 , n19210 , n19211 , n19212 ,
     n19213 , n19214 , n19215 , n19216 , n19217 , n19218 , n19219 , n19220 , n19221 , n19222 ,
     n19223 , n19224 , n19225 , n19226 , n19227 , n19228 , n19229 , n19230 , n19231 , n19232 ,
     n19233 , n19234 , n19235 , n19236 , n19237 , n19238 , n19239 , n19240 , n19241 , n19242 ,
     n19243 , n19244 , n19245 , n19246 , n19247 , n19248 , n19249 , n19250 , n19251 , n19252 ,
     n19253 , n19254 , n19255 , n19256 , n19257 , n19258 , n19259 , n19260 , n19261 , n19262 ,
     n19263 , n19264 , n19265 , n19266 , n19267 , n19268 , n19269 , n19270 , n19271 , n19272 ,
     n19273 , n19274 , n19275 , n19276 , n19277 , n19278 , n19279 , n19280 , n19281 , n19282 ,
     n19283 , n19284 , n19285 , n19286 , n19287 , n19288 , n19289 , n19290 , n19291 , n19292 ,
     n19293 , n19294 , n19295 , n19296 , n19297 , n19298 , n19299 , n19300 , n19301 , n19302 ,
     n19303 , n19304 , n19305 , n19306 , n19307 , n19308 , n19309 , n19310 , n19311 , n19312 ,
     n19313 , n19314 , n19315 , n19316 , n19317 , n19318 , n19319 , n19320 , n19321 , n19322 ,
     n19323 , n19324 , n19325 , n19326 , n19327 , n19328 , n19329 , n19330 , n19331 , n19332 ,
     n19333 , n19334 , n19335 , n19336 , n19337 , n19338 , n19339 , n19340 , n19341 , n19342 ,
     n19343 , n19344 , n19345 , n19346 , n19347 , n19348 , n19349 , n19350 , n19351 , n19352 ,
     n19353 , n19354 , n19355 , n19356 , n19357 , n19358 , n19359 , n19360 , n19361 , n19362 ,
     n19363 , n19364 , n19365 , n19366 , n19367 , n19368 , n19369 , n19370 , n19371 , n19372 ,
     n19373 , n19374 , n19375 , n19376 , n19377 , n19378 , n19379 , n19380 , n19381 , n19382 ,
     n19383 , n19384 , n19385 , n19386 , n19387 , n19388 , n19389 , n19390 , n19391 , n19392 ,
     n19393 , n19394 , n19395 , n19396 , n19397 , n19398 , n19399 , n19400 , n19401 , n19402 ,
     n19403 , n19404 , n19405 , n19406 , n19407 , n19408 , n19409 , n19410 , n19411 , n19412 ,
     n19413 , n19414 , n19415 , n19416 , n19417 , n19418 , n19419 , n19420 , n19421 , n19422 ,
     n19423 , n19424 , n19425 , n19426 , n19427 , n19428 , n19429 , n19430 , n19431 , n19432 ,
     n19433 , n19434 , n19435 , n19436 , n19437 , n19438 , n19439 , n19440 , n19441 , n19442 ,
     n19443 , n19444 , n19445 , n19446 , n19447 , n19448 , n19449 , n19450 , n19451 , n19452 ,
     n19453 , n19454 , n19455 , n19456 , n19457 , n19458 , n19459 , n19460 , n19461 , n19462 ,
     n19463 , n19464 , n19465 , n19466 , n19467 , n19468 , n19469 , n19470 , n19471 , n19472 ,
     n19473 , n19474 , n19475 , n19476 , n19477 , n19478 , n19479 , n19480 , n19481 , n19482 ,
     n19483 , n19484 , n19485 , n19486 , n19487 , n19488 , n19489 , n19490 , n19491 , n19492 ,
     n19493 , n19494 , n19495 , n19496 , n19497 , n19498 , n19499 , n19500 , n19501 , n19502 ,
     n19503 , n19504 , n19505 , n19506 , n19507 , n19508 , n19509 , n19510 , n19511 , n19512 ,
     n19513 , n19514 , n19515 , n19516 , n19517 , n19518 , n19519 , n19520 , n19521 , n19522 ,
     n19523 , n19524 , n19525 , n19526 , n19527 , n19528 , n19529 , n19530 , n19531 , n19532 ,
     n19533 , n19534 , n19535 , n19536 , n19537 , n19538 , n19539 , n19540 , n19541 , n19542 ,
     n19543 , n19544 , n19545 , n19546 , n19547 , n19548 , n19549 , n19550 , n19551 , n19552 ,
     n19553 , n19554 , n19555 , n19556 , n19557 , n19558 , n19559 , n19560 , n19561 , n19562 ,
     n19563 , n19564 , n19565 , n19566 , n19567 , n19568 , n19569 , n19570 , n19571 , n19572 ,
     n19573 , n19574 , n19575 , n19576 , n19577 , n19578 , n19579 , n19580 , n19581 , n19582 ,
     n19583 , n19584 , n19585 , n19586 , n19587 , n19588 , n19589 , n19590 , n19591 , n19592 ,
     n19593 , n19594 , n19595 , n19596 , n19597 , n19598 , n19599 , n19600 , n19601 , n19602 ,
     n19603 , n19604 , n19605 , n19606 , n19607 , n19608 , n19609 , n19610 , n19611 , n19612 ,
     n19613 , n19614 , n19615 , n19616 , n19617 , n19618 , n19619 , n19620 , n19621 , n19622 ,
     n19623 , n19624 , n19625 , n19626 , n19627 , n19628 , n19629 , n19630 , n19631 , n19632 ,
     n19633 , n19634 , n19635 , n19636 , n19637 , n19638 , n19639 , n19640 , n19641 , n19642 ,
     n19643 , n19644 , n19645 , n19646 , n19647 , n19648 , n19649 , n19650 , n19651 , n19652 ,
     n19653 , n19654 , n19655 , n19656 , n19657 , n19658 , n19659 , n19660 , n19661 , n19662 ,
     n19663 , n19664 , n19665 , n19666 , n19667 , n19668 , n19669 , n19670 , n19671 , n19672 ,
     n19673 , n19674 , n19675 , n19676 , n19677 , n19678 , n19679 , n19680 , n19681 , n19682 ,
     n19683 , n19684 , n19685 , n19686 , n19687 , n19688 , n19689 , n19690 , n19691 , n19692 ,
     n19693 , n19694 , n19695 , n19696 , n19697 , n19698 , n19699 , n19700 , n19701 , n19702 ,
     n19703 , n19704 , n19705 , n19706 , n19707 , n19708 , n19709 , n19710 , n19711 , n19712 ,
     n19713 , n19714 , n19715 , n19716 , n19717 , n19718 , n19719 , n19720 , n19721 , n19722 ,
     n19723 , n19724 , n19725 , n19726 , n19727 , n19728 , n19729 , n19730 , n19731 , n19732 ,
     n19733 , n19734 , n19735 , n19736 , n19737 , n19738 , n19739 , n19740 , n19741 , n19742 ,
     n19743 , n19744 , n19745 , n19746 , n19747 , n19748 , n19749 , n19750 , n19751 , n19752 ,
     n19753 , n19754 , n19755 , n19756 , n19757 , n19758 , n19759 , n19760 , n19761 , n19762 ,
     n19763 , n19764 , n19765 , n19766 , n19767 , n19768 , n19769 , n19770 , n19771 , n19772 ,
     n19773 , n19774 , n19775 , n19776 , n19777 , n19778 , n19779 , n19780 , n19781 , n19782 ,
     n19783 , n19784 , n19785 , n19786 , n19787 , n19788 , n19789 , n19790 , n19791 , n19792 ,
     n19793 , n19794 , n19795 , n19796 , n19797 , n19798 , n19799 , n19800 , n19801 , n19802 ,
     n19803 , n19804 , n19805 , n19806 , n19807 , n19808 , n19809 , n19810 , n19811 , n19812 ,
     n19813 , n19814 , n19815 , n19816 , n19817 , n19818 , n19819 , n19820 , n19821 , n19822 ,
     n19823 , n19824 , n19825 , n19826 , n19827 , n19828 , n19829 , n19830 , n19831 , n19832 ,
     n19833 , n19834 , n19835 , n19836 , n19837 , n19838 , n19839 , n19840 , n19841 , n19842 ,
     n19843 , n19844 , n19845 , n19846 , n19847 , n19848 , n19849 , n19850 , n19851 , n19852 ,
     n19853 , n19854 , n19855 , n19856 , n19857 , n19858 , n19859 , n19860 , n19861 , n19862 ,
     n19863 , n19864 , n19865 , n19866 , n19867 , n19868 , n19869 , n19870 , n19871 , n19872 ,
     n19873 , n19874 , n19875 , n19876 , n19877 , n19878 , n19879 , n19880 , n19881 , n19882 ,
     n19883 , n19884 , n19885 , n19886 , n19887 , n19888 , n19889 , n19890 , n19891 , n19892 ,
     n19893 , n19894 , n19895 , n19896 , n19897 , n19898 , n19899 , n19900 , n19901 , n19902 ,
     n19903 , n19904 , n19905 , n19906 , n19907 , n19908 , n19909 , n19910 , n19911 , n19912 ,
     n19913 , n19914 , n19915 , n19916 , n19917 , n19918 , n19919 , n19920 , n19921 , n19922 ,
     n19923 , n19924 , n19925 , n19926 , n19927 , n19928 , n19929 , n19930 , n19931 , n19932 ,
     n19933 , n19934 , n19935 , n19936 , n19937 , n19938 , n19939 , n19940 , n19941 , n19942 ,
     n19943 , n19944 , n19945 , n19946 , n19947 , n19948 , n19949 , n19950 , n19951 , n19952 ,
     n19953 , n19954 , n19955 , n19956 , n19957 , n19958 , n19959 , n19960 , n19961 , n19962 ,
     n19963 , n19964 , n19965 , n19966 , n19967 , n19968 , n19969 , n19970 , n19971 , n19972 ,
     n19973 , n19974 , n19975 , n19976 , n19977 , n19978 , n19979 , n19980 , n19981 , n19982 ,
     n19983 , n19984 , n19985 , n19986 , n19987 , n19988 , n19989 , n19990 , n19991 , n19992 ,
     n19993 , n19994 , n19995 , n19996 , n19997 , n19998 , n19999 , n20000 , n20001 , n20002 ,
     n20003 , n20004 , n20005 , n20006 , n20007 , n20008 , n20009 , n20010 , n20011 , n20012 ,
     n20013 , n20014 , n20015 , n20016 , n20017 , n20018 , n20019 , n20020 , n20021 , n20022 ,
     n20023 , n20024 , n20025 , n20026 , n20027 , n20028 , n20029 , n20030 , n20031 , n20032 ,
     n20033 , n20034 , n20035 , n20036 , n20037 , n20038 , n20039 , n20040 , n20041 , n20042 ,
     n20043 , n20044 , n20045 , n20046 , n20047 , n20048 , n20049 , n20050 , n20051 , n20052 ,
     n20053 , n20054 , n20055 , n20056 , n20057 , n20058 , n20059 , n20060 , n20061 , n20062 ,
     n20063 , n20064 , n20065 , n20066 , n20067 , n20068 , n20069 , n20070 , n20071 , n20072 ,
     n20073 , n20074 , n20075 , n20076 , n20077 , n20078 , n20079 , n20080 , n20081 , n20082 ,
     n20083 , n20084 , n20085 , n20086 , n20087 , n20088 , n20089 , n20090 , n20091 , n20092 ,
     n20093 , n20094 , n20095 , n20096 , n20097 , n20098 , n20099 , n20100 , n20101 , n20102 ,
     n20103 , n20104 , n20105 , n20106 , n20107 , n20108 , n20109 , n20110 , n20111 , n20112 ,
     n20113 , n20114 , n20115 , n20116 , n20117 , n20118 , n20119 , n20120 , n20121 , n20122 ,
     n20123 , n20124 , n20125 , n20126 , n20127 , n20128 , n20129 , n20130 , n20131 , n20132 ,
     n20133 , n20134 , n20135 , n20136 , n20137 , n20138 , n20139 , n20140 , n20141 , n20142 ,
     n20143 , n20144 , n20145 , n20146 , n20147 , n20148 , n20149 , n20150 , n20151 , n20152 ,
     n20153 , n20154 , n20155 , n20156 , n20157 , n20158 , n20159 , n20160 , n20161 , n20162 ,
     n20163 , n20164 , n20165 , n20166 , n20167 , n20168 , n20169 , n20170 , n20171 , n20172 ,
     n20173 , n20174 , n20175 , n20176 , n20177 , n20178 , n20179 , n20180 , n20181 , n20182 ,
     n20183 , n20184 , n20185 , n20186 , n20187 , n20188 , n20189 , n20190 , n20191 , n20192 ,
     n20193 , n20194 , n20195 , n20196 , n20197 , n20198 , n20199 , n20200 , n20201 , n20202 ,
     n20203 , n20204 , n20205 , n20206 , n20207 , n20208 , n20209 , n20210 , n20211 , n20212 ,
     n20213 , n20214 , n20215 , n20216 , n20217 , n20218 , n20219 , n20220 , n20221 , n20222 ,
     n20223 , n20224 , n20225 , n20226 , n20227 , n20228 , n20229 , n20230 , n20231 , n20232 ,
     n20233 , n20234 , n20235 , n20236 , n20237 , n20238 , n20239 , n20240 , n20241 , n20242 ,
     n20243 , n20244 , n20245 , n20246 , n20247 , n20248 , n20249 , n20250 , n20251 , n20252 ,
     n20253 , n20254 , n20255 , n20256 , n20257 , n20258 , n20259 , n20260 , n20261 , n20262 ,
     n20263 , n20264 , n20265 , n20266 , n20267 , n20268 , n20269 , n20270 , n20271 , n20272 ,
     n20273 , n20274 , n20275 , n20276 , n20277 , n20278 , n20279 , n20280 , n20281 , n20282 ,
     n20283 , n20284 , n20285 , n20286 , n20287 , n20288 , n20289 , n20290 , n20291 , n20292 ,
     n20293 , n20294 , n20295 , n20296 , n20297 , n20298 , n20299 , n20300 , n20301 , n20302 ,
     n20303 , n20304 , n20305 , n20306 , n20307 , n20308 , n20309 , n20310 , n20311 , n20312 ,
     n20313 , n20314 , n20315 , n20316 , n20317 , n20318 , n20319 , n20320 , n20321 , n20322 ,
     n20323 , n20324 , n20325 , n20326 , n20327 , n20328 , n20329 , n20330 , n20331 , n20332 ,
     n20333 , n20334 , n20335 , n20336 , n20337 , n20338 , n20339 , n20340 , n20341 , n20342 ,
     n20343 , n20344 , n20345 , n20346 , n20347 , n20348 , n20349 , n20350 , n20351 , n20352 ,
     n20353 , n20354 , n20355 , n20356 , n20357 , n20358 , n20359 , n20360 , n20361 , n20362 ,
     n20363 , n20364 , n20365 , n20366 , n20367 , n20368 , n20369 , n20370 , n20371 , n20372 ,
     n20373 , n20374 , n20375 , n20376 , n20377 , n20378 , n20379 , n20380 , n20381 , n20382 ,
     n20383 , n20384 , n20385 , n20386 , n20387 , n20388 , n20389 , n20390 , n20391 , n20392 ,
     n20393 , n20394 , n20395 , n20396 , n20397 , n20398 , n20399 , n20400 , n20401 , n20402 ,
     n20403 , n20404 , n20405 , n20406 , n20407 , n20408 , n20409 , n20410 , n20411 , n20412 ,
     n20413 , n20414 , n20415 , n20416 , n20417 , n20418 , n20419 , n20420 , n20421 , n20422 ,
     n20423 , n20424 , n20425 , n20426 , n20427 , n20428 , n20429 , n20430 , n20431 , n20432 ,
     n20433 , n20434 , n20435 , n20436 , n20437 , n20438 , n20439 , n20440 , n20441 , n20442 ,
     n20443 , n20444 , n20445 , n20446 , n20447 , n20448 , n20449 , n20450 , n20451 , n20452 ,
     n20453 , n20454 , n20455 , n20456 , n20457 , n20458 , n20459 , n20460 , n20461 , n20462 ,
     n20463 , n20464 , n20465 , n20466 , n20467 , n20468 , n20469 , n20470 , n20471 , n20472 ,
     n20473 , n20474 , n20475 , n20476 , n20477 , n20478 , n20479 , n20480 , n20481 , n20482 ,
     n20483 , n20484 , n20485 , n20486 , n20487 , n20488 , n20489 , n20490 , n20491 , n20492 ,
     n20493 , n20494 , n20495 , n20496 , n20497 , n20498 , n20499 , n20500 , n20501 , n20502 ,
     n20503 , n20504 , n20505 , n20506 , n20507 , n20508 , n20509 , n20510 , n20511 , n20512 ,
     n20513 , n20514 , n20515 , n20516 , n20517 , n20518 , n20519 , n20520 , n20521 , n20522 ,
     n20523 , n20524 , n20525 , n20526 , n20527 , n20528 , n20529 , n20530 , n20531 , n20532 ,
     n20533 , n20534 , n20535 , n20536 , n20537 , n20538 , n20539 , n20540 , n20541 , n20542 ,
     n20543 , n20544 , n20545 , n20546 , n20547 , n20548 , n20549 , n20550 , n20551 , n20552 ,
     n20553 , n20554 , n20555 , n20556 , n20557 , n20558 , n20559 , n20560 , n20561 , n20562 ,
     n20563 , n20564 , n20565 , n20566 , n20567 , n20568 , n20569 , n20570 , n20571 , n20572 ,
     n20573 , n20574 , n20575 , n20576 , n20577 , n20578 , n20579 , n20580 , n20581 , n20582 ,
     n20583 , n20584 , n20585 , n20586 , n20587 , n20588 , n20589 , n20590 , n20591 , n20592 ,
     n20593 , n20594 , n20595 , n20596 , n20597 , n20598 , n20599 , n20600 , n20601 , n20602 ,
     n20603 , n20604 , n20605 , n20606 , n20607 , n20608 , n20609 , n20610 , n20611 , n20612 ,
     n20613 , n20614 , n20615 , n20616 , n20617 , n20618 , n20619 , n20620 , n20621 , n20622 ,
     n20623 , n20624 , n20625 , n20626 , n20627 , n20628 , n20629 , n20630 , n20631 , n20632 ,
     n20633 , n20634 , n20635 , n20636 , n20637 , n20638 , n20639 , n20640 , n20641 , n20642 ,
     n20643 , n20644 , n20645 , n20646 , n20647 , n20648 , n20649 , n20650 , n20651 , n20652 ,
     n20653 , n20654 , n20655 , n20656 , n20657 , n20658 , n20659 , n20660 , n20661 , n20662 ,
     n20663 , n20664 , n20665 , n20666 , n20667 , n20668 , n20669 , n20670 , n20671 , n20672 ,
     n20673 , n20674 , n20675 , n20676 , n20677 , n20678 , n20679 , n20680 , n20681 , n20682 ,
     n20683 , n20684 , n20685 , n20686 , n20687 , n20688 , n20689 , n20690 , n20691 , n20692 ,
     n20693 , n20694 , n20695 , n20696 , n20697 , n20698 , n20699 , n20700 , n20701 , n20702 ,
     n20703 , n20704 , n20705 , n20706 , n20707 , n20708 , n20709 , n20710 , n20711 , n20712 ,
     n20713 , n20714 , n20715 , n20716 , n20717 , n20718 , n20719 , n20720 , n20721 , n20722 ,
     n20723 , n20724 , n20725 , n20726 , n20727 , n20728 , n20729 , n20730 , n20731 , n20732 ,
     n20733 , n20734 , n20735 , n20736 , n20737 , n20738 , n20739 , n20740 , n20741 , n20742 ,
     n20743 , n20744 , n20745 , n20746 , n20747 , n20748 , n20749 , n20750 , n20751 , n20752 ,
     n20753 , n20754 , n20755 , n20756 , n20757 , n20758 , n20759 , n20760 , n20761 , n20762 ,
     n20763 , n20764 , n20765 , n20766 , n20767 , n20768 , n20769 , n20770 , n20771 , n20772 ,
     n20773 , n20774 , n20775 , n20776 , n20777 , n20778 , n20779 , n20780 , n20781 , n20782 ,
     n20783 , n20784 , n20785 , n20786 , n20787 , n20788 , n20789 , n20790 , n20791 , n20792 ,
     n20793 , n20794 , n20795 , n20796 , n20797 , n20798 , n20799 , n20800 , n20801 , n20802 ,
     n20803 , n20804 , n20805 , n20806 , n20807 , n20808 , n20809 , n20810 , n20811 , n20812 ,
     n20813 , n20814 , n20815 , n20816 , n20817 , n20818 , n20819 , n20820 , n20821 , n20822 ,
     n20823 , n20824 , n20825 , n20826 , n20827 , n20828 , n20829 , n20830 , n20831 , n20832 ,
     n20833 , n20834 , n20835 , n20836 , n20837 , n20838 , n20839 , n20840 , n20841 , n20842 ,
     n20843 , n20844 , n20845 , n20846 , n20847 , n20848 , n20849 , n20850 , n20851 , n20852 ,
     n20853 , n20854 , n20855 , n20856 , n20857 , n20858 , n20859 , n20860 , n20861 , n20862 ,
     n20863 , n20864 , n20865 , n20866 , n20867 , n20868 , n20869 , n20870 , n20871 , n20872 ,
     n20873 , n20874 , n20875 , n20876 , n20877 , n20878 , n20879 , n20880 , n20881 , n20882 ,
     n20883 , n20884 , n20885 , n20886 , n20887 , n20888 , n20889 , n20890 , n20891 , n20892 ,
     n20893 , n20894 , n20895 , n20896 , n20897 , n20898 , n20899 , n20900 , n20901 , n20902 ,
     n20903 , n20904 , n20905 , n20906 , n20907 , n20908 , n20909 , n20910 , n20911 , n20912 ,
     n20913 , n20914 , n20915 , n20916 , n20917 , n20918 , n20919 , n20920 , n20921 , n20922 ,
     n20923 , n20924 , n20925 , n20926 , n20927 , n20928 , n20929 , n20930 , n20931 , n20932 ,
     n20933 , n20934 , n20935 , n20936 , n20937 , n20938 , n20939 , n20940 , n20941 , n20942 ,
     n20943 , n20944 , n20945 , n20946 , n20947 , n20948 , n20949 , n20950 , n20951 , n20952 ,
     n20953 , n20954 , n20955 , n20956 , n20957 , n20958 , n20959 , n20960 , n20961 , n20962 ,
     n20963 , n20964 , n20965 , n20966 , n20967 , n20968 , n20969 , n20970 , n20971 , n20972 ,
     n20973 , n20974 , n20975 , n20976 , n20977 , n20978 , n20979 , n20980 , n20981 , n20982 ,
     n20983 , n20984 , n20985 , n20986 , n20987 , n20988 , n20989 , n20990 , n20991 , n20992 ,
     n20993 , n20994 , n20995 , n20996 , n20997 , n20998 , n20999 , n21000 , n21001 , n21002 ,
     n21003 , n21004 , n21005 , n21006 , n21007 , n21008 , n21009 , n21010 , n21011 , n21012 ,
     n21013 , n21014 , n21015 , n21016 , n21017 , n21018 , n21019 , n21020 , n21021 , n21022 ,
     n21023 , n21024 , n21025 , n21026 , n21027 , n21028 , n21029 , n21030 , n21031 , n21032 ,
     n21033 , n21034 , n21035 , n21036 , n21037 , n21038 , n21039 , n21040 , n21041 , n21042 ,
     n21043 , n21044 , n21045 , n21046 , n21047 , n21048 , n21049 , n21050 , n21051 , n21052 ,
     n21053 , n21054 , n21055 , n21056 , n21057 , n21058 , n21059 , n21060 , n21061 , n21062 ,
     n21063 , n21064 , n21065 , n21066 , n21067 , n21068 , n21069 , n21070 , n21071 , n21072 ,
     n21073 , n21074 , n21075 , n21076 , n21077 , n21078 , n21079 , n21080 , n21081 , n21082 ,
     n21083 , n21084 , n21085 , n21086 , n21087 , n21088 , n21089 , n21090 , n21091 , n21092 ,
     n21093 , n21094 , n21095 , n21096 , n21097 , n21098 , n21099 , n21100 , n21101 , n21102 ,
     n21103 , n21104 , n21105 , n21106 , n21107 , n21108 , n21109 , n21110 , n21111 , n21112 ,
     n21113 , n21114 , n21115 , n21116 , n21117 , n21118 , n21119 , n21120 , n21121 , n21122 ,
     n21123 , n21124 , n21125 , n21126 , n21127 , n21128 , n21129 , n21130 , n21131 , n21132 ,
     n21133 , n21134 , n21135 , n21136 , n21137 , n21138 , n21139 , n21140 , n21141 , n21142 ,
     n21143 , n21144 , n21145 , n21146 , n21147 , n21148 , n21149 , n21150 , n21151 , n21152 ,
     n21153 , n21154 , n21155 , n21156 , n21157 , n21158 , n21159 , n21160 , n21161 , n21162 ,
     n21163 , n21164 , n21165 , n21166 , n21167 , n21168 , n21169 , n21170 , n21171 , n21172 ,
     n21173 , n21174 , n21175 , n21176 , n21177 , n21178 , n21179 , n21180 , n21181 , n21182 ,
     n21183 , n21184 , n21185 , n21186 , n21187 , n21188 , n21189 , n21190 , n21191 , n21192 ,
     n21193 , n21194 , n21195 , n21196 , n21197 , n21198 , n21199 , n21200 , n21201 , n21202 ,
     n21203 , n21204 , n21205 , n21206 , n21207 , n21208 , n21209 , n21210 , n21211 , n21212 ,
     n21213 , n21214 , n21215 , n21216 , n21217 , n21218 , n21219 , n21220 , n21221 , n21222 ,
     n21223 , n21224 , n21225 , n21226 , n21227 , n21228 , n21229 , n21230 , n21231 , n21232 ,
     n21233 , n21234 , n21235 , n21236 , n21237 , n21238 , n21239 , n21240 , n21241 , n21242 ,
     n21243 , n21244 , n21245 , n21246 , n21247 , n21248 , n21249 , n21250 , n21251 , n21252 ,
     n21253 , n21254 , n21255 , n21256 , n21257 , n21258 , n21259 , n21260 , n21261 , n21262 ,
     n21263 , n21264 , n21265 , n21266 , n21267 , n21268 , n21269 , n21270 , n21271 , n21272 ,
     n21273 , n21274 , n21275 , n21276 , n21277 , n21278 , n21279 , n21280 , n21281 , n21282 ,
     n21283 , n21284 , n21285 , n21286 , n21287 , n21288 , n21289 , n21290 , n21291 , n21292 ,
     n21293 , n21294 , n21295 , n21296 , n21297 , n21298 , n21299 , n21300 , n21301 , n21302 ,
     n21303 , n21304 , n21305 , n21306 , n21307 , n21308 , n21309 , n21310 , n21311 , n21312 ,
     n21313 , n21314 , n21315 , n21316 , n21317 , n21318 , n21319 , n21320 , n21321 , n21322 ,
     n21323 , n21324 , n21325 , n21326 , n21327 , n21328 , n21329 , n21330 , n21331 , n21332 ,
     n21333 , n21334 , n21335 , n21336 , n21337 , n21338 , n21339 , n21340 , n21341 , n21342 ,
     n21343 , n21344 , n21345 , n21346 , n21347 , n21348 , n21349 , n21350 , n21351 , n21352 ,
     n21353 , n21354 , n21355 , n21356 , n21357 , n21358 , n21359 , n21360 , n21361 , n21362 ,
     n21363 , n21364 , n21365 , n21366 , n21367 , n21368 , n21369 , n21370 , n21371 , n21372 ,
     n21373 , n21374 , n21375 , n21376 , n21377 , n21378 , n21379 , n21380 , n21381 , n21382 ,
     n21383 , n21384 , n21385 , n21386 , n21387 , n21388 , n21389 , n21390 , n21391 , n21392 ,
     n21393 , n21394 , n21395 , n21396 , n21397 , n21398 , n21399 , n21400 , n21401 , n21402 ,
     n21403 , n21404 , n21405 , n21406 , n21407 , n21408 , n21409 , n21410 , n21411 , n21412 ,
     n21413 , n21414 , n21415 , n21416 , n21417 , n21418 , n21419 , n21420 , n21421 , n21422 ,
     n21423 , n21424 , n21425 , n21426 , n21427 , n21428 , n21429 , n21430 , n21431 , n21432 ,
     n21433 , n21434 , n21435 , n21436 , n21437 , n21438 , n21439 , n21440 , n21441 , n21442 ,
     n21443 , n21444 , n21445 , n21446 , n21447 , n21448 , n21449 , n21450 , n21451 , n21452 ,
     n21453 , n21454 , n21455 , n21456 , n21457 , n21458 , n21459 , n21460 , n21461 , n21462 ,
     n21463 , n21464 , n21465 , n21466 , n21467 , n21468 , n21469 , n21470 , n21471 , n21472 ,
     n21473 , n21474 , n21475 , n21476 , n21477 , n21478 , n21479 , n21480 , n21481 , n21482 ,
     n21483 , n21484 , n21485 , n21486 , n21487 , n21488 , n21489 , n21490 , n21491 , n21492 ,
     n21493 , n21494 , n21495 , n21496 , n21497 , n21498 , n21499 , n21500 , n21501 , n21502 ,
     n21503 , n21504 , n21505 , n21506 , n21507 , n21508 , n21509 , n21510 , n21511 , n21512 ,
     n21513 , n21514 , n21515 , n21516 , n21517 , n21518 , n21519 , n21520 , n21521 , n21522 ,
     n21523 , n21524 , n21525 , n21526 , n21527 , n21528 , n21529 , n21530 , n21531 , n21532 ,
     n21533 , n21534 , n21535 , n21536 , n21537 , n21538 , n21539 , n21540 , n21541 , n21542 ,
     n21543 , n21544 , n21545 , n21546 , n21547 , n21548 , n21549 , n21550 , n21551 , n21552 ,
     n21553 , n21554 , n21555 , n21556 , n21557 , n21558 , n21559 , n21560 , n21561 , n21562 ,
     n21563 , n21564 , n21565 , n21566 , n21567 , n21568 , n21569 , n21570 , n21571 , n21572 ,
     n21573 , n21574 , n21575 , n21576 , n21577 , n21578 , n21579 , n21580 , n21581 , n21582 ,
     n21583 , n21584 , n21585 , n21586 , n21587 , n21588 , n21589 , n21590 , n21591 , n21592 ,
     n21593 , n21594 , n21595 , n21596 , n21597 , n21598 , n21599 , n21600 , n21601 , n21602 ,
     n21603 , n21604 , n21605 , n21606 , n21607 , n21608 , n21609 , n21610 , n21611 , n21612 ,
     n21613 , n21614 , n21615 , n21616 , n21617 , n21618 , n21619 , n21620 , n21621 , n21622 ,
     n21623 , n21624 , n21625 , n21626 , n21627 , n21628 , n21629 , n21630 , n21631 , n21632 ,
     n21633 , n21634 , n21635 , n21636 , n21637 , n21638 , n21639 , n21640 , n21641 , n21642 ,
     n21643 , n21644 , n21645 , n21646 , n21647 , n21648 , n21649 , n21650 , n21651 , n21652 ,
     n21653 , n21654 , n21655 , n21656 , n21657 , n21658 , n21659 , n21660 , n21661 , n21662 ,
     n21663 , n21664 , n21665 , n21666 , n21667 , n21668 , n21669 , n21670 , n21671 , n21672 ,
     n21673 , n21674 , n21675 , n21676 , n21677 , n21678 , n21679 , n21680 , n21681 , n21682 ,
     n21683 , n21684 , n21685 , n21686 , n21687 , n21688 , n21689 , n21690 , n21691 , n21692 ,
     n21693 , n21694 , n21695 , n21696 , n21697 , n21698 , n21699 , n21700 , n21701 , n21702 ,
     n21703 , n21704 , n21705 , n21706 , n21707 , n21708 , n21709 , n21710 , n21711 , n21712 ,
     n21713 , n21714 , n21715 , n21716 , n21717 , n21718 , n21719 , n21720 , n21721 , n21722 ,
     n21723 , n21724 , n21725 , n21726 , n21727 , n21728 , n21729 , n21730 , n21731 , n21732 ,
     n21733 , n21734 , n21735 , n21736 , n21737 , n21738 , n21739 , n21740 , n21741 , n21742 ,
     n21743 , n21744 , n21745 , n21746 , n21747 , n21748 , n21749 , n21750 , n21751 , n21752 ,
     n21753 , n21754 , n21755 , n21756 , n21757 , n21758 , n21759 , n21760 , n21761 , n21762 ,
     n21763 , n21764 , n21765 , n21766 , n21767 , n21768 , n21769 , n21770 , n21771 , n21772 ,
     n21773 , n21774 , n21775 , n21776 , n21777 , n21778 , n21779 , n21780 , n21781 , n21782 ,
     n21783 , n21784 , n21785 , n21786 , n21787 , n21788 , n21789 , n21790 , n21791 , n21792 ,
     n21793 , n21794 , n21795 , n21796 , n21797 , n21798 , n21799 , n21800 , n21801 , n21802 ,
     n21803 , n21804 , n21805 , n21806 , n21807 , n21808 , n21809 , n21810 , n21811 , n21812 ,
     n21813 , n21814 , n21815 , n21816 , n21817 , n21818 , n21819 , n21820 , n21821 , n21822 ,
     n21823 , n21824 , n21825 , n21826 , n21827 , n21828 , n21829 , n21830 , n21831 , n21832 ,
     n21833 , n21834 , n21835 , n21836 , n21837 , n21838 , n21839 , n21840 , n21841 , n21842 ,
     n21843 , n21844 , n21845 , n21846 , n21847 , n21848 , n21849 , n21850 , n21851 , n21852 ,
     n21853 , n21854 , n21855 , n21856 , n21857 , n21858 , n21859 , n21860 , n21861 , n21862 ,
     n21863 , n21864 , n21865 , n21866 , n21867 , n21868 , n21869 , n21870 , n21871 , n21872 ,
     n21873 , n21874 , n21875 , n21876 , n21877 , n21878 , n21879 , n21880 , n21881 , n21882 ,
     n21883 , n21884 , n21885 , n21886 , n21887 , n21888 , n21889 , n21890 , n21891 , n21892 ,
     n21893 , n21894 , n21895 , n21896 , n21897 , n21898 , n21899 , n21900 , n21901 , n21902 ,
     n21903 , n21904 , n21905 , n21906 , n21907 , n21908 , n21909 , n21910 , n21911 , n21912 ,
     n21913 , n21914 , n21915 , n21916 , n21917 , n21918 , n21919 , n21920 , n21921 , n21922 ,
     n21923 , n21924 , n21925 , n21926 , n21927 , n21928 , n21929 , n21930 , n21931 , n21932 ,
     n21933 , n21934 , n21935 , n21936 , n21937 , n21938 , n21939 , n21940 , n21941 , n21942 ,
     n21943 , n21944 , n21945 , n21946 , n21947 , n21948 , n21949 , n21950 , n21951 , n21952 ,
     n21953 , n21954 , n21955 , n21956 , n21957 , n21958 , n21959 , n21960 , n21961 , n21962 ,
     n21963 , n21964 , n21965 , n21966 , n21967 , n21968 , n21969 , n21970 , n21971 , n21972 ,
     n21973 , n21974 , n21975 , n21976 , n21977 , n21978 , n21979 , n21980 , n21981 , n21982 ,
     n21983 , n21984 , n21985 , n21986 , n21987 , n21988 , n21989 , n21990 , n21991 , n21992 ,
     n21993 , n21994 , n21995 , n21996 , n21997 , n21998 , n21999 , n22000 , n22001 , n22002 ,
     n22003 , n22004 , n22005 , n22006 , n22007 , n22008 , n22009 , n22010 , n22011 , n22012 ,
     n22013 , n22014 , n22015 , n22016 , n22017 , n22018 , n22019 , n22020 , n22021 , n22022 ,
     n22023 , n22024 , n22025 , n22026 , n22027 , n22028 , n22029 , n22030 , n22031 , n22032 ,
     n22033 , n22034 , n22035 , n22036 , n22037 , n22038 , n22039 , n22040 , n22041 , n22042 ,
     n22043 , n22044 , n22045 , n22046 , n22047 , n22048 , n22049 , n22050 , n22051 , n22052 ,
     n22053 , n22054 , n22055 , n22056 , n22057 , n22058 , n22059 , n22060 , n22061 , n22062 ,
     n22063 , n22064 , n22065 , n22066 , n22067 , n22068 , n22069 , n22070 , n22071 , n22072 ,
     n22073 , n22074 , n22075 , n22076 , n22077 , n22078 , n22079 , n22080 , n22081 , n22082 ,
     n22083 , n22084 , n22085 , n22086 , n22087 , n22088 , n22089 , n22090 , n22091 , n22092 ,
     n22093 , n22094 , n22095 , n22096 , n22097 , n22098 , n22099 , n22100 , n22101 , n22102 ,
     n22103 , n22104 , n22105 , n22106 , n22107 , n22108 , n22109 , n22110 , n22111 , n22112 ,
     n22113 , n22114 , n22115 , n22116 , n22117 , n22118 , n22119 , n22120 , n22121 , n22122 ,
     n22123 , n22124 , n22125 , n22126 , n22127 , n22128 , n22129 , n22130 , n22131 , n22132 ,
     n22133 , n22134 , n22135 , n22136 , n22137 , n22138 , n22139 , n22140 , n22141 , n22142 ,
     n22143 , n22144 , n22145 , n22146 , n22147 , n22148 , n22149 , n22150 , n22151 , n22152 ,
     n22153 , n22154 , n22155 , n22156 , n22157 , n22158 , n22159 , n22160 , n22161 , n22162 ,
     n22163 , n22164 , n22165 , n22166 , n22167 , n22168 , n22169 , n22170 , n22171 , n22172 ,
     n22173 , n22174 , n22175 , n22176 , n22177 , n22178 , n22179 , n22180 , n22181 , n22182 ,
     n22183 , n22184 , n22185 , n22186 , n22187 , n22188 , n22189 , n22190 , n22191 , n22192 ,
     n22193 , n22194 , n22195 , n22196 , n22197 , n22198 , n22199 , n22200 , n22201 , n22202 ,
     n22203 , n22204 , n22205 , n22206 , n22207 , n22208 , n22209 , n22210 , n22211 , n22212 ,
     n22213 , n22214 , n22215 , n22216 , n22217 , n22218 , n22219 , n22220 , n22221 , n22222 ,
     n22223 , n22224 , n22225 , n22226 , n22227 , n22228 , n22229 , n22230 , n22231 , n22232 ,
     n22233 , n22234 , n22235 , n22236 , n22237 , n22238 , n22239 , n22240 , n22241 , n22242 ,
     n22243 , n22244 , n22245 , n22246 , n22247 , n22248 , n22249 , n22250 , n22251 , n22252 ,
     n22253 , n22254 , n22255 , n22256 , n22257 , n22258 , n22259 , n22260 , n22261 , n22262 ,
     n22263 , n22264 , n22265 , n22266 , n22267 , n22268 , n22269 , n22270 , n22271 , n22272 ,
     n22273 , n22274 , n22275 , n22276 , n22277 , n22278 , n22279 , n22280 , n22281 , n22282 ,
     n22283 , n22284 , n22285 , n22286 , n22287 , n22288 , n22289 , n22290 , n22291 , n22292 ,
     n22293 , n22294 , n22295 , n22296 , n22297 , n22298 , n22299 , n22300 , n22301 , n22302 ,
     n22303 , n22304 , n22305 , n22306 , n22307 , n22308 , n22309 , n22310 , n22311 , n22312 ,
     n22313 , n22314 , n22315 , n22316 , n22317 , n22318 , n22319 , n22320 , n22321 , n22322 ,
     n22323 , n22324 , n22325 , n22326 , n22327 , n22328 , n22329 , n22330 , n22331 , n22332 ,
     n22333 , n22334 , n22335 , n22336 , n22337 , n22338 , n22339 , n22340 , n22341 , n22342 ,
     n22343 , n22344 , n22345 , n22346 , n22347 , n22348 , n22349 , n22350 , n22351 , n22352 ,
     n22353 , n22354 , n22355 , n22356 , n22357 , n22358 , n22359 , n22360 , n22361 , n22362 ,
     n22363 , n22364 , n22365 , n22366 , n22367 , n22368 , n22369 , n22370 , n22371 , n22372 ,
     n22373 , n22374 , n22375 , n22376 , n22377 , n22378 , n22379 , n22380 , n22381 , n22382 ,
     n22383 , n22384 , n22385 , n22386 , n22387 , n22388 , n22389 , n22390 , n22391 , n22392 ,
     n22393 , n22394 , n22395 , n22396 , n22397 , n22398 , n22399 , n22400 , n22401 , n22402 ,
     n22403 , n22404 , n22405 , n22406 , n22407 , n22408 , n22409 , n22410 , n22411 , n22412 ,
     n22413 , n22414 , n22415 , n22416 , n22417 , n22418 , n22419 , n22420 , n22421 , n22422 ,
     n22423 , n22424 , n22425 , n22426 , n22427 , n22428 , n22429 , n22430 , n22431 , n22432 ,
     n22433 , n22434 , n22435 , n22436 , n22437 , n22438 , n22439 , n22440 , n22441 , n22442 ,
     n22443 , n22444 , n22445 , n22446 , n22447 , n22448 , n22449 , n22450 , n22451 , n22452 ,
     n22453 , n22454 , n22455 , n22456 , n22457 , n22458 , n22459 , n22460 , n22461 , n22462 ,
     n22463 , n22464 , n22465 , n22466 , n22467 , n22468 , n22469 , n22470 , n22471 , n22472 ,
     n22473 , n22474 , n22475 , n22476 , n22477 , n22478 , n22479 , n22480 , n22481 , n22482 ,
     n22483 , n22484 , n22485 , n22486 , n22487 , n22488 , n22489 , n22490 , n22491 , n22492 ,
     n22493 , n22494 , n22495 , n22496 , n22497 , n22498 , n22499 , n22500 , n22501 , n22502 ,
     n22503 , n22504 , n22505 , n22506 , n22507 , n22508 , n22509 , n22510 , n22511 , n22512 ,
     n22513 , n22514 , n22515 , n22516 , n22517 , n22518 , n22519 , n22520 , n22521 , n22522 ,
     n22523 , n22524 , n22525 , n22526 , n22527 , n22528 , n22529 , n22530 , n22531 , n22532 ,
     n22533 , n22534 , n22535 , n22536 , n22537 , n22538 , n22539 , n22540 , n22541 , n22542 ,
     n22543 , n22544 , n22545 , n22546 , n22547 , n22548 , n22549 , n22550 , n22551 , n22552 ,
     n22553 , n22554 , n22555 , n22556 , n22557 , n22558 , n22559 , n22560 , n22561 , n22562 ,
     n22563 , n22564 , n22565 , n22566 , n22567 , n22568 , n22569 , n22570 , n22571 , n22572 ,
     n22573 , n22574 , n22575 , n22576 , n22577 , n22578 , n22579 , n22580 , n22581 , n22582 ,
     n22583 , n22584 , n22585 , n22586 , n22587 , n22588 , n22589 , n22590 , n22591 , n22592 ,
     n22593 , n22594 , n22595 , n22596 , n22597 , n22598 , n22599 , n22600 , n22601 , n22602 ,
     n22603 , n22604 , n22605 , n22606 , n22607 , n22608 , n22609 , n22610 , n22611 , n22612 ,
     n22613 , n22614 , n22615 , n22616 , n22617 , n22618 , n22619 , n22620 , n22621 , n22622 ,
     n22623 , n22624 , n22625 , n22626 , n22627 , n22628 , n22629 , n22630 , n22631 , n22632 ,
     n22633 , n22634 , n22635 , n22636 , n22637 , n22638 , n22639 , n22640 , n22641 , n22642 ,
     n22643 , n22644 , n22645 , n22646 , n22647 , n22648 , n22649 , n22650 , n22651 , n22652 ,
     n22653 , n22654 , n22655 , n22656 , n22657 , n22658 , n22659 , n22660 , n22661 , n22662 ,
     n22663 , n22664 , n22665 , n22666 , n22667 , n22668 , n22669 , n22670 , n22671 , n22672 ,
     n22673 , n22674 , n22675 , n22676 , n22677 , n22678 , n22679 , n22680 , n22681 , n22682 ,
     n22683 , n22684 , n22685 , n22686 , n22687 , n22688 , n22689 , n22690 , n22691 , n22692 ,
     n22693 , n22694 , n22695 , n22696 , n22697 , n22698 , n22699 , n22700 , n22701 , n22702 ,
     n22703 , n22704 , n22705 , n22706 , n22707 , n22708 , n22709 , n22710 , n22711 , n22712 ,
     n22713 , n22714 , n22715 , n22716 , n22717 , n22718 , n22719 , n22720 , n22721 , n22722 ,
     n22723 , n22724 , n22725 , n22726 , n22727 , n22728 , n22729 , n22730 , n22731 , n22732 ,
     n22733 , n22734 , n22735 , n22736 , n22737 , n22738 , n22739 , n22740 , n22741 , n22742 ,
     n22743 , n22744 , n22745 , n22746 , n22747 , n22748 , n22749 , n22750 , n22751 , n22752 ,
     n22753 , n22754 , n22755 , n22756 , n22757 , n22758 , n22759 , n22760 , n22761 , n22762 ,
     n22763 , n22764 , n22765 , n22766 , n22767 , n22768 , n22769 , n22770 , n22771 , n22772 ,
     n22773 , n22774 , n22775 , n22776 , n22777 , n22778 , n22779 , n22780 , n22781 , n22782 ,
     n22783 , n22784 , n22785 , n22786 , n22787 , n22788 , n22789 , n22790 , n22791 , n22792 ,
     n22793 , n22794 , n22795 , n22796 , n22797 , n22798 , n22799 , n22800 , n22801 , n22802 ,
     n22803 , n22804 , n22805 , n22806 , n22807 , n22808 , n22809 , n22810 , n22811 , n22812 ,
     n22813 , n22814 , n22815 , n22816 , n22817 , n22818 , n22819 , n22820 , n22821 , n22822 ,
     n22823 , n22824 , n22825 , n22826 , n22827 , n22828 , n22829 , n22830 , n22831 , n22832 ,
     n22833 , n22834 , n22835 , n22836 , n22837 , n22838 , n22839 , n22840 , n22841 , n22842 ,
     n22843 , n22844 , n22845 , n22846 , n22847 , n22848 , n22849 , n22850 , n22851 , n22852 ,
     n22853 , n22854 , n22855 , n22856 , n22857 , n22858 , n22859 , n22860 , n22861 , n22862 ,
     n22863 , n22864 , n22865 , n22866 , n22867 , n22868 , n22869 , n22870 , n22871 , n22872 ,
     n22873 , n22874 , n22875 , n22876 , n22877 , n22878 , n22879 , n22880 , n22881 , n22882 ,
     n22883 , n22884 , n22885 , n22886 , n22887 , n22888 , n22889 , n22890 , n22891 , n22892 ,
     n22893 , n22894 , n22895 , n22896 , n22897 , n22898 , n22899 , n22900 , n22901 , n22902 ,
     n22903 , n22904 , n22905 , n22906 , n22907 , n22908 , n22909 , n22910 , n22911 , n22912 ,
     n22913 , n22914 , n22915 , n22916 , n22917 , n22918 , n22919 , n22920 , n22921 , n22922 ,
     n22923 , n22924 , n22925 , n22926 , n22927 , n22928 , n22929 , n22930 , n22931 , n22932 ,
     n22933 , n22934 , n22935 , n22936 , n22937 , n22938 , n22939 , n22940 , n22941 , n22942 ,
     n22943 , n22944 , n22945 , n22946 , n22947 , n22948 , n22949 , n22950 , n22951 , n22952 ,
     n22953 , n22954 , n22955 , n22956 , n22957 , n22958 , n22959 , n22960 , n22961 , n22962 ,
     n22963 , n22964 , n22965 , n22966 , n22967 , n22968 , n22969 , n22970 , n22971 , n22972 ,
     n22973 , n22974 , n22975 , n22976 , n22977 , n22978 , n22979 , n22980 , n22981 , n22982 ,
     n22983 , n22984 , n22985 , n22986 , n22987 , n22988 , n22989 , n22990 , n22991 , n22992 ,
     n22993 , n22994 , n22995 , n22996 , n22997 , n22998 , n22999 , n23000 , n23001 , n23002 ,
     n23003 , n23004 , n23005 , n23006 , n23007 , n23008 , n23009 , n23010 , n23011 , n23012 ,
     n23013 , n23014 , n23015 , n23016 , n23017 , n23018 , n23019 , n23020 , n23021 , n23022 ,
     n23023 , n23024 , n23025 , n23026 , n23027 , n23028 , n23029 , n23030 , n23031 , n23032 ,
     n23033 , n23034 , n23035 , n23036 , n23037 , n23038 , n23039 , n23040 , n23041 , n23042 ,
     n23043 , n23044 , n23045 , n23046 , n23047 , n23048 , n23049 , n23050 , n23051 , n23052 ,
     n23053 , n23054 , n23055 , n23056 , n23057 , n23058 , n23059 , n23060 , n23061 , n23062 ,
     n23063 , n23064 , n23065 , n23066 , n23067 , n23068 , n23069 , n23070 , n23071 , n23072 ,
     n23073 , n23074 , n23075 , n23076 , n23077 , n23078 , n23079 , n23080 , n23081 , n23082 ,
     n23083 , n23084 , n23085 , n23086 , n23087 , n23088 , n23089 , n23090 , n23091 , n23092 ,
     n23093 , n23094 , n23095 , n23096 , n23097 , n23098 , n23099 , n23100 , n23101 , n23102 ,
     n23103 , n23104 , n23105 , n23106 , n23107 , n23108 , n23109 , n23110 , n23111 , n23112 ,
     n23113 , n23114 , n23115 , n23116 , n23117 , n23118 , n23119 , n23120 , n23121 , n23122 ,
     n23123 , n23124 , n23125 , n23126 , n23127 , n23128 , n23129 , n23130 , n23131 , n23132 ,
     n23133 , n23134 , n23135 , n23136 , n23137 , n23138 , n23139 , n23140 , n23141 , n23142 ,
     n23143 , n23144 , n23145 , n23146 , n23147 , n23148 , n23149 , n23150 , n23151 , n23152 ,
     n23153 , n23154 , n23155 , n23156 , n23157 , n23158 , n23159 , n23160 , n23161 , n23162 ,
     n23163 , n23164 , n23165 , n23166 , n23167 , n23168 , n23169 , n23170 , n23171 , n23172 ,
     n23173 , n23174 , n23175 , n23176 , n23177 , n23178 , n23179 , n23180 , n23181 , n23182 ,
     n23183 , n23184 , n23185 , n23186 , n23187 , n23188 , n23189 , n23190 , n23191 , n23192 ,
     n23193 , n23194 , n23195 , n23196 , n23197 , n23198 , n23199 , n23200 , n23201 , n23202 ,
     n23203 , n23204 , n23205 , n23206 , n23207 , n23208 , n23209 , n23210 , n23211 , n23212 ,
     n23213 , n23214 , n23215 , n23216 , n23217 , n23218 , n23219 , n23220 , n23221 , n23222 ,
     n23223 , n23224 , n23225 , n23226 , n23227 , n23228 , n23229 , n23230 , n23231 , n23232 ,
     n23233 , n23234 , n23235 , n23236 , n23237 , n23238 , n23239 , n23240 , n23241 , n23242 ,
     n23243 , n23244 , n23245 , n23246 , n23247 , n23248 , n23249 , n23250 , n23251 , n23252 ,
     n23253 , n23254 , n23255 , n23256 , n23257 , n23258 , n23259 , n23260 , n23261 , n23262 ,
     n23263 , n23264 , n23265 , n23266 , n23267 , n23268 , n23269 , n23270 , n23271 , n23272 ,
     n23273 , n23274 , n23275 , n23276 , n23277 , n23278 , n23279 , n23280 , n23281 , n23282 ,
     n23283 , n23284 , n23285 , n23286 , n23287 , n23288 , n23289 , n23290 , n23291 , n23292 ,
     n23293 , n23294 , n23295 , n23296 , n23297 , n23298 , n23299 , n23300 , n23301 , n23302 ,
     n23303 , n23304 , n23305 , n23306 , n23307 , n23308 , n23309 , n23310 , n23311 , n23312 ,
     n23313 , n23314 , n23315 , n23316 , n23317 , n23318 , n23319 , n23320 , n23321 , n23322 ,
     n23323 , n23324 , n23325 , n23326 , n23327 , n23328 , n23329 , n23330 , n23331 , n23332 ,
     n23333 , n23334 , n23335 , n23336 , n23337 , n23338 , n23339 , n23340 , n23341 , n23342 ,
     n23343 , n23344 , n23345 , n23346 , n23347 , n23348 , n23349 , n23350 , n23351 , n23352 ,
     n23353 , n23354 , n23355 , n23356 , n23357 , n23358 , n23359 , n23360 , n23361 , n23362 ,
     n23363 , n23364 , n23365 , n23366 , n23367 , n23368 , n23369 , n23370 , n23371 , n23372 ,
     n23373 , n23374 , n23375 , n23376 , n23377 , n23378 , n23379 , n23380 , n23381 , n23382 ,
     n23383 , n23384 , n23385 , n23386 , n23387 , n23388 , n23389 , n23390 , n23391 , n23392 ,
     n23393 , n23394 , n23395 , n23396 , n23397 , n23398 , n23399 , n23400 , n23401 , n23402 ,
     n23403 , n23404 , n23405 , n23406 , n23407 , n23408 , n23409 , n23410 , n23411 , n23412 ,
     n23413 , n23414 , n23415 , n23416 , n23417 , n23418 , n23419 , n23420 , n23421 , n23422 ,
     n23423 , n23424 , n23425 , n23426 , n23427 , n23428 , n23429 , n23430 , n23431 , n23432 ,
     n23433 , n23434 , n23435 , n23436 , n23437 , n23438 , n23439 , n23440 , n23441 , n23442 ,
     n23443 , n23444 , n23445 , n23446 , n23447 , n23448 , n23449 , n23450 , n23451 , n23452 ,
     n23453 , n23454 , n23455 , n23456 , n23457 , n23458 , n23459 , n23460 , n23461 , n23462 ,
     n23463 , n23464 , n23465 , n23466 , n23467 , n23468 , n23469 , n23470 , n23471 , n23472 ,
     n23473 , n23474 , n23475 , n23476 , n23477 , n23478 , n23479 , n23480 , n23481 , n23482 ,
     n23483 , n23484 , n23485 , n23486 , n23487 , n23488 , n23489 , n23490 , n23491 , n23492 ,
     n23493 , n23494 , n23495 , n23496 , n23497 , n23498 , n23499 , n23500 , n23501 , n23502 ,
     n23503 , n23504 , n23505 , n23506 , n23507 , n23508 , n23509 , n23510 , n23511 , n23512 ,
     n23513 , n23514 , n23515 , n23516 , n23517 , n23518 , n23519 , n23520 , n23521 , n23522 ,
     n23523 , n23524 , n23525 , n23526 , n23527 , n23528 , n23529 , n23530 , n23531 , n23532 ,
     n23533 , n23534 , n23535 , n23536 , n23537 , n23538 , n23539 , n23540 , n23541 , n23542 ,
     n23543 , n23544 , n23545 , n23546 , n23547 , n23548 , n23549 , n23550 , n23551 , n23552 ,
     n23553 , n23554 , n23555 , n23556 , n23557 , n23558 , n23559 , n23560 , n23561 , n23562 ,
     n23563 , n23564 , n23565 , n23566 , n23567 , n23568 , n23569 , n23570 , n23571 , n23572 ,
     n23573 , n23574 , n23575 , n23576 , n23577 , n23578 , n23579 , n23580 , n23581 , n23582 ,
     n23583 , n23584 , n23585 , n23586 , n23587 , n23588 , n23589 , n23590 , n23591 , n23592 ,
     n23593 , n23594 , n23595 , n23596 , n23597 , n23598 , n23599 , n23600 , n23601 , n23602 ,
     n23603 , n23604 , n23605 , n23606 , n23607 , n23608 , n23609 , n23610 , n23611 , n23612 ,
     n23613 , n23614 , n23615 , n23616 , n23617 , n23618 , n23619 , n23620 , n23621 , n23622 ,
     n23623 , n23624 , n23625 , n23626 , n23627 , n23628 , n23629 , n23630 , n23631 , n23632 ,
     n23633 , n23634 , n23635 , n23636 , n23637 , n23638 , n23639 , n23640 , n23641 , n23642 ,
     n23643 , n23644 , n23645 , n23646 , n23647 , n23648 , n23649 , n23650 , n23651 , n23652 ,
     n23653 , n23654 , n23655 , n23656 , n23657 , n23658 , n23659 , n23660 , n23661 , n23662 ,
     n23663 , n23664 , n23665 , n23666 , n23667 , n23668 , n23669 , n23670 , n23671 , n23672 ,
     n23673 , n23674 , n23675 , n23676 , n23677 , n23678 , n23679 , n23680 , n23681 , n23682 ,
     n23683 , n23684 , n23685 , n23686 , n23687 , n23688 , n23689 , n23690 , n23691 , n23692 ,
     n23693 , n23694 , n23695 , n23696 , n23697 , n23698 , n23699 , n23700 , n23701 , n23702 ,
     n23703 , n23704 , n23705 , n23706 , n23707 , n23708 , n23709 , n23710 , n23711 , n23712 ,
     n23713 , n23714 , n23715 , n23716 , n23717 , n23718 , n23719 , n23720 , n23721 , n23722 ,
     n23723 , n23724 , n23725 , n23726 , n23727 , n23728 , n23729 , n23730 , n23731 , n23732 ,
     n23733 , n23734 , n23735 , n23736 , n23737 , n23738 , n23739 , n23740 , n23741 , n23742 ,
     n23743 , n23744 , n23745 , n23746 , n23747 , n23748 , n23749 , n23750 , n23751 , n23752 ,
     n23753 , n23754 , n23755 , n23756 , n23757 , n23758 , n23759 , n23760 , n23761 , n23762 ,
     n23763 , n23764 , n23765 , n23766 , n23767 , n23768 , n23769 , n23770 , n23771 , n23772 ,
     n23773 , n23774 , n23775 , n23776 , n23777 , n23778 , n23779 , n23780 , n23781 , n23782 ,
     n23783 , n23784 , n23785 , n23786 , n23787 , n23788 , n23789 , n23790 , n23791 , n23792 ,
     n23793 , n23794 , n23795 , n23796 , n23797 , n23798 , n23799 , n23800 , n23801 , n23802 ,
     n23803 , n23804 , n23805 , n23806 , n23807 , n23808 , n23809 , n23810 , n23811 , n23812 ,
     n23813 , n23814 , n23815 , n23816 , n23817 , n23818 , n23819 , n23820 , n23821 , n23822 ,
     n23823 , n23824 , n23825 , n23826 , n23827 , n23828 , n23829 , n23830 , n23831 , n23832 ,
     n23833 , n23834 , n23835 , n23836 , n23837 , n23838 , n23839 , n23840 , n23841 , n23842 ,
     n23843 , n23844 , n23845 , n23846 , n23847 , n23848 , n23849 , n23850 , n23851 , n23852 ,
     n23853 , n23854 , n23855 , n23856 , n23857 , n23858 , n23859 , n23860 , n23861 , n23862 ,
     n23863 , n23864 , n23865 , n23866 , n23867 , n23868 , n23869 , n23870 , n23871 , n23872 ,
     n23873 , n23874 , n23875 , n23876 , n23877 , n23878 , n23879 , n23880 , n23881 , n23882 ,
     n23883 , n23884 , n23885 , n23886 , n23887 , n23888 , n23889 , n23890 , n23891 , n23892 ,
     n23893 , n23894 , n23895 , n23896 , n23897 , n23898 , n23899 , n23900 , n23901 , n23902 ,
     n23903 , n23904 , n23905 , n23906 , n23907 , n23908 , n23909 , n23910 , n23911 , n23912 ,
     n23913 , n23914 , n23915 , n23916 , n23917 , n23918 , n23919 , n23920 , n23921 , n23922 ,
     n23923 , n23924 , n23925 , n23926 , n23927 , n23928 , n23929 , n23930 , n23931 , n23932 ,
     n23933 , n23934 , n23935 , n23936 , n23937 , n23938 , n23939 , n23940 , n23941 , n23942 ,
     n23943 , n23944 , n23945 , n23946 , n23947 , n23948 , n23949 , n23950 , n23951 , n23952 ,
     n23953 , n23954 , n23955 , n23956 , n23957 , n23958 , n23959 , n23960 , n23961 , n23962 ,
     n23963 , n23964 , n23965 , n23966 , n23967 , n23968 , n23969 , n23970 , n23971 , n23972 ,
     n23973 , n23974 , n23975 , n23976 , n23977 , n23978 , n23979 , n23980 , n23981 , n23982 ,
     n23983 , n23984 , n23985 , n23986 , n23987 , n23988 , n23989 , n23990 , n23991 , n23992 ,
     n23993 , n23994 , n23995 , n23996 , n23997 , n23998 , n23999 , n24000 , n24001 , n24002 ,
     n24003 , n24004 , n24005 , n24006 , n24007 , n24008 , n24009 , n24010 , n24011 , n24012 ,
     n24013 , n24014 , n24015 , n24016 , n24017 , n24018 , n24019 , n24020 , n24021 , n24022 ,
     n24023 , n24024 , n24025 , n24026 , n24027 , n24028 , n24029 , n24030 , n24031 , n24032 ,
     n24033 , n24034 , n24035 , n24036 , n24037 , n24038 , n24039 , n24040 , n24041 , n24042 ,
     n24043 , n24044 , n24045 , n24046 , n24047 , n24048 , n24049 , n24050 , n24051 , n24052 ,
     n24053 , n24054 , n24055 , n24056 , n24057 , n24058 , n24059 , n24060 , n24061 , n24062 ,
     n24063 , n24064 , n24065 , n24066 , n24067 , n24068 , n24069 , n24070 , n24071 , n24072 ,
     n24073 , n24074 , n24075 , n24076 , n24077 , n24078 , n24079 , n24080 , n24081 , n24082 ,
     n24083 , n24084 , n24085 , n24086 , n24087 , n24088 , n24089 , n24090 , n24091 , n24092 ,
     n24093 , n24094 , n24095 , n24096 , n24097 , n24098 , n24099 , n24100 , n24101 , n24102 ,
     n24103 , n24104 , n24105 , n24106 , n24107 , n24108 , n24109 , n24110 , n24111 , n24112 ,
     n24113 , n24114 , n24115 , n24116 , n24117 , n24118 , n24119 , n24120 , n24121 , n24122 ,
     n24123 , n24124 , n24125 , n24126 , n24127 , n24128 , n24129 , n24130 , n24131 , n24132 ,
     n24133 , n24134 , n24135 , n24136 , n24137 , n24138 , n24139 , n24140 , n24141 , n24142 ,
     n24143 , n24144 , n24145 , n24146 , n24147 , n24148 , n24149 , n24150 , n24151 , n24152 ,
     n24153 , n24154 , n24155 , n24156 , n24157 , n24158 , n24159 , n24160 , n24161 , n24162 ,
     n24163 , n24164 , n24165 , n24166 , n24167 , n24168 , n24169 , n24170 , n24171 , n24172 ,
     n24173 , n24174 , n24175 , n24176 , n24177 , n24178 , n24179 , n24180 , n24181 , n24182 ,
     n24183 , n24184 , n24185 , n24186 , n24187 , n24188 , n24189 , n24190 , n24191 , n24192 ,
     n24193 , n24194 , n24195 , n24196 , n24197 , n24198 , n24199 , n24200 , n24201 , n24202 ,
     n24203 , n24204 , n24205 , n24206 , n24207 , n24208 , n24209 , n24210 , n24211 , n24212 ,
     n24213 , n24214 , n24215 , n24216 , n24217 , n24218 , n24219 , n24220 , n24221 , n24222 ,
     n24223 , n24224 , n24225 , n24226 , n24227 , n24228 , n24229 , n24230 , n24231 , n24232 ,
     n24233 , n24234 , n24235 , n24236 , n24237 , n24238 , n24239 , n24240 , n24241 , n24242 ,
     n24243 , n24244 , n24245 , n24246 , n24247 , n24248 , n24249 , n24250 , n24251 , n24252 ,
     n24253 , n24254 , n24255 , n24256 , n24257 , n24258 , n24259 , n24260 , n24261 , n24262 ,
     n24263 , n24264 , n24265 , n24266 , n24267 , n24268 , n24269 , n24270 , n24271 , n24272 ,
     n24273 , n24274 , n24275 , n24276 , n24277 , n24278 , n24279 , n24280 , n24281 , n24282 ,
     n24283 , n24284 , n24285 , n24286 , n24287 , n24288 , n24289 , n24290 , n24291 , n24292 ,
     n24293 , n24294 , n24295 , n24296 , n24297 , n24298 , n24299 , n24300 , n24301 , n24302 ,
     n24303 , n24304 , n24305 , n24306 , n24307 , n24308 , n24309 , n24310 , n24311 , n24312 ,
     n24313 , n24314 , n24315 , n24316 , n24317 , n24318 , n24319 , n24320 , n24321 , n24322 ,
     n24323 , n24324 , n24325 , n24326 , n24327 , n24328 , n24329 , n24330 , n24331 , n24332 ,
     n24333 , n24334 , n24335 , n24336 , n24337 , n24338 , n24339 , n24340 , n24341 , n24342 ,
     n24343 , n24344 , n24345 , n24346 , n24347 , n24348 , n24349 , n24350 , n24351 , n24352 ,
     n24353 , n24354 , n24355 , n24356 , n24357 , n24358 , n24359 , n24360 , n24361 , n24362 ,
     n24363 , n24364 , n24365 , n24366 , n24367 , n24368 , n24369 , n24370 , n24371 , n24372 ,
     n24373 , n24374 , n24375 , n24376 , n24377 , n24378 , n24379 , n24380 , n24381 , n24382 ,
     n24383 , n24384 , n24385 , n24386 , n24387 , n24388 , n24389 , n24390 , n24391 , n24392 ,
     n24393 , n24394 , n24395 , n24396 , n24397 , n24398 , n24399 , n24400 , n24401 , n24402 ,
     n24403 , n24404 , n24405 , n24406 , n24407 , n24408 , n24409 , n24410 , n24411 , n24412 ,
     n24413 , n24414 , n24415 , n24416 , n24417 , n24418 , n24419 , n24420 , n24421 , n24422 ,
     n24423 , n24424 , n24425 , n24426 , n24427 , n24428 , n24429 , n24430 , n24431 , n24432 ,
     n24433 , n24434 , n24435 , n24436 , n24437 , n24438 , n24439 , n24440 , n24441 , n24442 ,
     n24443 , n24444 , n24445 , n24446 , n24447 , n24448 , n24449 , n24450 , n24451 , n24452 ,
     n24453 , n24454 , n24455 , n24456 , n24457 , n24458 , n24459 , n24460 , n24461 , n24462 ,
     n24463 , n24464 , n24465 , n24466 , n24467 , n24468 , n24469 , n24470 , n24471 , n24472 ,
     n24473 , n24474 , n24475 , n24476 , n24477 , n24478 , n24479 , n24480 , n24481 , n24482 ,
     n24483 , n24484 , n24485 , n24486 , n24487 , n24488 , n24489 , n24490 , n24491 , n24492 ,
     n24493 , n24494 , n24495 , n24496 , n24497 , n24498 , n24499 , n24500 , n24501 , n24502 ,
     n24503 , n24504 , n24505 , n24506 , n24507 , n24508 , n24509 , n24510 , n24511 , n24512 ,
     n24513 , n24514 , n24515 , n24516 , n24517 , n24518 , n24519 , n24520 , n24521 , n24522 ,
     n24523 , n24524 , n24525 , n24526 , n24527 , n24528 , n24529 , n24530 , n24531 , n24532 ,
     n24533 , n24534 , n24535 , n24536 , n24537 , n24538 , n24539 , n24540 , n24541 , n24542 ,
     n24543 , n24544 , n24545 , n24546 , n24547 , n24548 , n24549 , n24550 , n24551 , n24552 ,
     n24553 , n24554 , n24555 , n24556 , n24557 , n24558 , n24559 , n24560 , n24561 , n24562 ,
     n24563 , n24564 , n24565 , n24566 , n24567 , n24568 , n24569 , n24570 , n24571 , n24572 ,
     n24573 , n24574 , n24575 , n24576 , n24577 , n24578 , n24579 , n24580 , n24581 , n24582 ,
     n24583 , n24584 , n24585 , n24586 , n24587 , n24588 , n24589 , n24590 , n24591 , n24592 ,
     n24593 , n24594 , n24595 , n24596 , n24597 , n24598 , n24599 , n24600 , n24601 , n24602 ,
     n24603 , n24604 , n24605 , n24606 , n24607 , n24608 , n24609 , n24610 , n24611 , n24612 ,
     n24613 , n24614 , n24615 , n24616 , n24617 , n24618 , n24619 , n24620 , n24621 , n24622 ,
     n24623 , n24624 , n24625 , n24626 , n24627 , n24628 , n24629 , n24630 , n24631 , n24632 ,
     n24633 , n24634 , n24635 , n24636 , n24637 , n24638 , n24639 , n24640 , n24641 , n24642 ,
     n24643 , n24644 , n24645 , n24646 , n24647 , n24648 , n24649 , n24650 , n24651 , n24652 ,
     n24653 , n24654 , n24655 , n24656 , n24657 , n24658 , n24659 , n24660 , n24661 , n24662 ,
     n24663 , n24664 , n24665 , n24666 , n24667 , n24668 , n24669 , n24670 , n24671 , n24672 ,
     n24673 , n24674 , n24675 , n24676 , n24677 , n24678 , n24679 , n24680 , n24681 , n24682 ,
     n24683 , n24684 , n24685 , n24686 , n24687 , n24688 , n24689 , n24690 , n24691 , n24692 ,
     n24693 , n24694 , n24695 , n24696 , n24697 , n24698 , n24699 , n24700 , n24701 , n24702 ,
     n24703 , n24704 , n24705 , n24706 , n24707 , n24708 , n24709 , n24710 , n24711 , n24712 ,
     n24713 , n24714 , n24715 , n24716 , n24717 , n24718 , n24719 , n24720 , n24721 , n24722 ,
     n24723 , n24724 , n24725 , n24726 , n24727 , n24728 , n24729 , n24730 , n24731 , n24732 ,
     n24733 , n24734 , n24735 , n24736 , n24737 , n24738 , n24739 , n24740 , n24741 , n24742 ,
     n24743 , n24744 , n24745 , n24746 , n24747 , n24748 , n24749 , n24750 , n24751 , n24752 ,
     n24753 , n24754 , n24755 , n24756 , n24757 , n24758 , n24759 , n24760 , n24761 , n24762 ,
     n24763 , n24764 , n24765 , n24766 , n24767 , n24768 , n24769 , n24770 , n24771 , n24772 ,
     n24773 , n24774 , n24775 , n24776 , n24777 , n24778 , n24779 , n24780 , n24781 , n24782 ,
     n24783 , n24784 , n24785 , n24786 , n24787 , n24788 , n24789 , n24790 , n24791 , n24792 ,
     n24793 , n24794 , n24795 , n24796 , n24797 , n24798 , n24799 , n24800 , n24801 , n24802 ,
     n24803 , n24804 , n24805 , n24806 , n24807 , n24808 , n24809 , n24810 , n24811 , n24812 ,
     n24813 , n24814 , n24815 , n24816 , n24817 , n24818 , n24819 , n24820 , n24821 , n24822 ,
     n24823 , n24824 , n24825 , n24826 , n24827 , n24828 , n24829 , n24830 , n24831 , n24832 ,
     n24833 , n24834 , n24835 , n24836 , n24837 , n24838 , n24839 , n24840 , n24841 , n24842 ,
     n24843 , n24844 , n24845 , n24846 , n24847 , n24848 , n24849 , n24850 , n24851 , n24852 ,
     n24853 , n24854 , n24855 , n24856 , n24857 , n24858 , n24859 , n24860 , n24861 , n24862 ,
     n24863 , n24864 , n24865 , n24866 , n24867 , n24868 , n24869 , n24870 , n24871 , n24872 ,
     n24873 , n24874 , n24875 , n24876 , n24877 , n24878 , n24879 , n24880 , n24881 , n24882 ,
     n24883 , n24884 , n24885 , n24886 , n24887 , n24888 , n24889 , n24890 , n24891 , n24892 ,
     n24893 , n24894 , n24895 , n24896 , n24897 , n24898 , n24899 , n24900 , n24901 , n24902 ,
     n24903 , n24904 , n24905 , n24906 , n24907 , n24908 , n24909 , n24910 , n24911 , n24912 ,
     n24913 , n24914 , n24915 , n24916 , n24917 , n24918 , n24919 , n24920 , n24921 , n24922 ,
     n24923 , n24924 , n24925 , n24926 , n24927 , n24928 , n24929 , n24930 , n24931 , n24932 ,
     n24933 , n24934 , n24935 , n24936 , n24937 , n24938 , n24939 , n24940 , n24941 , n24942 ,
     n24943 , n24944 , n24945 , n24946 , n24947 , n24948 , n24949 , n24950 , n24951 , n24952 ,
     n24953 , n24954 , n24955 , n24956 , n24957 , n24958 , n24959 , n24960 , n24961 , n24962 ,
     n24963 , n24964 , n24965 , n24966 , n24967 , n24968 , n24969 , n24970 , n24971 , n24972 ,
     n24973 , n24974 , n24975 , n24976 , n24977 , n24978 , n24979 , n24980 , n24981 , n24982 ,
     n24983 , n24984 , n24985 , n24986 , n24987 , n24988 , n24989 , n24990 , n24991 , n24992 ,
     n24993 , n24994 , n24995 , n24996 , n24997 , n24998 , n24999 , n25000 , n25001 , n25002 ,
     n25003 , n25004 , n25005 , n25006 , n25007 , n25008 , n25009 , n25010 , n25011 , n25012 ,
     n25013 , n25014 , n25015 , n25016 , n25017 , n25018 , n25019 , n25020 , n25021 , n25022 ,
     n25023 , n25024 , n25025 , n25026 , n25027 , n25028 , n25029 , n25030 , n25031 , n25032 ,
     n25033 , n25034 , n25035 , n25036 , n25037 , n25038 , n25039 , n25040 , n25041 , n25042 ,
     n25043 , n25044 , n25045 , n25046 , n25047 , n25048 , n25049 , n25050 , n25051 , n25052 ,
     n25053 , n25054 , n25055 , n25056 , n25057 , n25058 , n25059 , n25060 , n25061 , n25062 ,
     n25063 , n25064 , n25065 , n25066 , n25067 , n25068 , n25069 , n25070 , n25071 , n25072 ,
     n25073 , n25074 , n25075 , n25076 , n25077 , n25078 , n25079 , n25080 , n25081 , n25082 ,
     n25083 , n25084 , n25085 , n25086 , n25087 , n25088 , n25089 , n25090 , n25091 , n25092 ,
     n25093 , n25094 , n25095 , n25096 , n25097 , n25098 , n25099 , n25100 , n25101 , n25102 ,
     n25103 , n25104 , n25105 , n25106 , n25107 , n25108 , n25109 , n25110 , n25111 , n25112 ,
     n25113 , n25114 , n25115 , n25116 , n25117 , n25118 , n25119 , n25120 , n25121 , n25122 ,
     n25123 , n25124 , n25125 , n25126 , n25127 , n25128 , n25129 , n25130 , n25131 , n25132 ,
     n25133 , n25134 , n25135 , n25136 , n25137 , n25138 , n25139 , n25140 , n25141 , n25142 ,
     n25143 , n25144 , n25145 , n25146 , n25147 , n25148 , n25149 , n25150 , n25151 , n25152 ,
     n25153 , n25154 , n25155 , n25156 , n25157 , n25158 , n25159 , n25160 , n25161 , n25162 ,
     n25163 , n25164 , n25165 , n25166 , n25167 , n25168 , n25169 , n25170 , n25171 , n25172 ,
     n25173 , n25174 , n25175 , n25176 , n25177 , n25178 , n25179 , n25180 , n25181 , n25182 ,
     n25183 , n25184 , n25185 , n25186 , n25187 , n25188 , n25189 , n25190 , n25191 , n25192 ,
     n25193 , n25194 , n25195 , n25196 , n25197 , n25198 , n25199 , n25200 , n25201 , n25202 ,
     n25203 , n25204 , n25205 , n25206 , n25207 , n25208 , n25209 , n25210 , n25211 , n25212 ,
     n25213 , n25214 , n25215 , n25216 , n25217 , n25218 , n25219 , n25220 , n25221 , n25222 ,
     n25223 , n25224 , n25225 , n25226 , n25227 , n25228 , n25229 , n25230 , n25231 , n25232 ,
     n25233 , n25234 , n25235 , n25236 , n25237 , n25238 , n25239 , n25240 , n25241 , n25242 ,
     n25243 , n25244 , n25245 , n25246 , n25247 , n25248 , n25249 , n25250 , n25251 , n25252 ,
     n25253 , n25254 , n25255 , n25256 , n25257 , n25258 , n25259 , n25260 , n25261 , n25262 ,
     n25263 , n25264 , n25265 , n25266 , n25267 , n25268 , n25269 , n25270 , n25271 , n25272 ,
     n25273 , n25274 , n25275 , n25276 , n25277 , n25278 , n25279 , n25280 , n25281 , n25282 ,
     n25283 , n25284 , n25285 , n25286 , n25287 , n25288 , n25289 , n25290 , n25291 , n25292 ,
     n25293 , n25294 , n25295 , n25296 , n25297 , n25298 , n25299 , n25300 , n25301 , n25302 ,
     n25303 , n25304 , n25305 , n25306 , n25307 , n25308 , n25309 , n25310 , n25311 , n25312 ,
     n25313 , n25314 , n25315 , n25316 , n25317 , n25318 , n25319 , n25320 , n25321 , n25322 ,
     n25323 , n25324 , n25325 , n25326 , n25327 , n25328 , n25329 , n25330 , n25331 , n25332 ,
     n25333 , n25334 , n25335 , n25336 , n25337 , n25338 , n25339 , n25340 , n25341 , n25342 ,
     n25343 , n25344 , n25345 , n25346 , n25347 , n25348 , n25349 , n25350 , n25351 , n25352 ,
     n25353 , n25354 , n25355 , n25356 , n25357 , n25358 , n25359 , n25360 , n25361 , n25362 ,
     n25363 , n25364 , n25365 , n25366 , n25367 , n25368 , n25369 , n25370 , n25371 , n25372 ,
     n25373 , n25374 , n25375 , n25376 , n25377 , n25378 , n25379 , n25380 , n25381 , n25382 ,
     n25383 , n25384 , n25385 , n25386 , n25387 , n25388 , n25389 , n25390 , n25391 , n25392 ,
     n25393 , n25394 , n25395 , n25396 , n25397 , n25398 , n25399 , n25400 , n25401 , n25402 ,
     n25403 , n25404 , n25405 , n25406 , n25407 , n25408 , n25409 , n25410 , n25411 , n25412 ,
     n25413 , n25414 , n25415 , n25416 , n25417 , n25418 , n25419 , n25420 , n25421 , n25422 ,
     n25423 , n25424 , n25425 , n25426 , n25427 , n25428 , n25429 , n25430 , n25431 , n25432 ,
     n25433 , n25434 , n25435 , n25436 , n25437 , n25438 , n25439 , n25440 , n25441 , n25442 ,
     n25443 , n25444 , n25445 , n25446 , n25447 , n25448 , n25449 , n25450 , n25451 , n25452 ,
     n25453 , n25454 , n25455 , n25456 , n25457 , n25458 , n25459 , n25460 , n25461 , n25462 ,
     n25463 , n25464 , n25465 , n25466 , n25467 , n25468 , n25469 , n25470 , n25471 , n25472 ,
     n25473 , n25474 , n25475 , n25476 , n25477 , n25478 , n25479 , n25480 , n25481 , n25482 ,
     n25483 , n25484 , n25485 , n25486 , n25487 , n25488 , n25489 , n25490 , n25491 , n25492 ,
     n25493 , n25494 , n25495 , n25496 , n25497 , n25498 , n25499 , n25500 , n25501 , n25502 ,
     n25503 , n25504 , n25505 , n25506 , n25507 , n25508 , n25509 , n25510 , n25511 , n25512 ,
     n25513 , n25514 , n25515 , n25516 , n25517 , n25518 , n25519 , n25520 , n25521 , n25522 ,
     n25523 , n25524 , n25525 , n25526 , n25527 , n25528 , n25529 , n25530 , n25531 , n25532 ,
     n25533 , n25534 , n25535 , n25536 , n25537 , n25538 , n25539 , n25540 , n25541 , n25542 ,
     n25543 , n25544 , n25545 , n25546 , n25547 , n25548 , n25549 , n25550 , n25551 , n25552 ,
     n25553 , n25554 , n25555 , n25556 , n25557 , n25558 , n25559 , n25560 , n25561 , n25562 ,
     n25563 , n25564 , n25565 , n25566 , n25567 , n25568 , n25569 , n25570 , n25571 , n25572 ,
     n25573 , n25574 , n25575 , n25576 , n25577 , n25578 , n25579 , n25580 , n25581 , n25582 ,
     n25583 , n25584 , n25585 , n25586 , n25587 , n25588 , n25589 , n25590 , n25591 , n25592 ,
     n25593 , n25594 , n25595 , n25596 , n25597 , n25598 , n25599 , n25600 , n25601 , n25602 ,
     n25603 , n25604 , n25605 , n25606 , n25607 , n25608 , n25609 , n25610 , n25611 , n25612 ,
     n25613 , n25614 , n25615 , n25616 , n25617 , n25618 , n25619 , n25620 , n25621 , n25622 ,
     n25623 , n25624 , n25625 , n25626 , n25627 , n25628 , n25629 , n25630 , n25631 , n25632 ,
     n25633 , n25634 , n25635 , n25636 , n25637 , n25638 , n25639 , n25640 , n25641 , n25642 ,
     n25643 , n25644 , n25645 , n25646 , n25647 , n25648 , n25649 , n25650 , n25651 , n25652 ,
     n25653 , n25654 , n25655 , n25656 , n25657 , n25658 , n25659 , n25660 , n25661 , n25662 ,
     n25663 , n25664 , n25665 , n25666 , n25667 , n25668 , n25669 , n25670 , n25671 , n25672 ,
     n25673 , n25674 , n25675 , n25676 , n25677 , n25678 , n25679 , n25680 , n25681 , n25682 ,
     n25683 , n25684 , n25685 , n25686 , n25687 , n25688 , n25689 , n25690 , n25691 , n25692 ,
     n25693 , n25694 , n25695 , n25696 , n25697 , n25698 , n25699 , n25700 , n25701 , n25702 ,
     n25703 , n25704 , n25705 , n25706 , n25707 , n25708 , n25709 , n25710 , n25711 , n25712 ,
     n25713 , n25714 , n25715 , n25716 , n25717 , n25718 , n25719 , n25720 , n25721 , n25722 ,
     n25723 , n25724 , n25725 , n25726 , n25727 , n25728 , n25729 , n25730 , n25731 , n25732 ,
     n25733 , n25734 , n25735 , n25736 , n25737 , n25738 , n25739 , n25740 , n25741 , n25742 ,
     n25743 , n25744 , n25745 , n25746 , n25747 , n25748 , n25749 , n25750 , n25751 , n25752 ,
     n25753 , n25754 , n25755 , n25756 , n25757 , n25758 , n25759 , n25760 , n25761 , n25762 ,
     n25763 , n25764 , n25765 , n25766 , n25767 , n25768 , n25769 , n25770 , n25771 , n25772 ,
     n25773 , n25774 , n25775 , n25776 , n25777 , n25778 , n25779 , n25780 , n25781 , n25782 ,
     n25783 , n25784 , n25785 , n25786 , n25787 , n25788 , n25789 , n25790 , n25791 , n25792 ,
     n25793 , n25794 , n25795 , n25796 , n25797 , n25798 , n25799 , n25800 , n25801 , n25802 ,
     n25803 , n25804 , n25805 , n25806 , n25807 , n25808 , n25809 , n25810 , n25811 , n25812 ,
     n25813 , n25814 , n25815 , n25816 , n25817 , n25818 , n25819 , n25820 , n25821 , n25822 ,
     n25823 , n25824 , n25825 , n25826 , n25827 , n25828 , n25829 , n25830 , n25831 , n25832 ,
     n25833 , n25834 , n25835 , n25836 , n25837 , n25838 , n25839 , n25840 , n25841 , n25842 ,
     n25843 , n25844 , n25845 , n25846 , n25847 , n25848 , n25849 , n25850 , n25851 , n25852 ,
     n25853 , n25854 , n25855 , n25856 , n25857 , n25858 , n25859 , n25860 , n25861 , n25862 ,
     n25863 , n25864 , n25865 , n25866 , n25867 , n25868 , n25869 , n25870 , n25871 , n25872 ,
     n25873 , n25874 , n25875 , n25876 , n25877 , n25878 , n25879 , n25880 , n25881 , n25882 ,
     n25883 , n25884 , n25885 , n25886 , n25887 , n25888 , n25889 , n25890 , n25891 , n25892 ,
     n25893 , n25894 , n25895 , n25896 , n25897 , n25898 , n25899 , n25900 , n25901 , n25902 ,
     n25903 , n25904 , n25905 , n25906 , n25907 , n25908 , n25909 , n25910 , n25911 , n25912 ,
     n25913 , n25914 , n25915 , n25916 , n25917 , n25918 , n25919 , n25920 , n25921 , n25922 ,
     n25923 , n25924 , n25925 , n25926 , n25927 , n25928 , n25929 , n25930 , n25931 , n25932 ,
     n25933 , n25934 , n25935 , n25936 , n25937 , n25938 , n25939 , n25940 , n25941 , n25942 ,
     n25943 , n25944 , n25945 , n25946 , n25947 , n25948 , n25949 , n25950 , n25951 , n25952 ,
     n25953 , n25954 , n25955 , n25956 , n25957 , n25958 , n25959 , n25960 , n25961 , n25962 ,
     n25963 , n25964 , n25965 , n25966 , n25967 , n25968 , n25969 , n25970 , n25971 , n25972 ,
     n25973 , n25974 , n25975 , n25976 , n25977 , n25978 , n25979 , n25980 , n25981 , n25982 ,
     n25983 , n25984 , n25985 , n25986 , n25987 , n25988 , n25989 , n25990 , n25991 , n25992 ,
     n25993 , n25994 , n25995 , n25996 , n25997 , n25998 , n25999 , n26000 , n26001 , n26002 ,
     n26003 , n26004 , n26005 , n26006 , n26007 , n26008 , n26009 , n26010 , n26011 , n26012 ,
     n26013 , n26014 , n26015 , n26016 , n26017 , n26018 , n26019 , n26020 , n26021 , n26022 ,
     n26023 , n26024 , n26025 , n26026 , n26027 , n26028 , n26029 , n26030 , n26031 , n26032 ,
     n26033 , n26034 , n26035 , n26036 , n26037 , n26038 , n26039 , n26040 , n26041 , n26042 ,
     n26043 , n26044 , n26045 , n26046 , n26047 , n26048 , n26049 , n26050 , n26051 , n26052 ,
     n26053 , n26054 , n26055 , n26056 , n26057 , n26058 , n26059 , n26060 , n26061 , n26062 ,
     n26063 , n26064 , n26065 , n26066 , n26067 , n26068 , n26069 , n26070 , n26071 , n26072 ,
     n26073 , n26074 , n26075 , n26076 , n26077 , n26078 , n26079 , n26080 , n26081 , n26082 ,
     n26083 , n26084 , n26085 , n26086 , n26087 , n26088 , n26089 , n26090 , n26091 , n26092 ,
     n26093 , n26094 , n26095 , n26096 , n26097 , n26098 , n26099 , n26100 , n26101 , n26102 ,
     n26103 , n26104 , n26105 , n26106 , n26107 , n26108 , n26109 , n26110 , n26111 , n26112 ,
     n26113 , n26114 , n26115 , n26116 , n26117 , n26118 , n26119 , n26120 , n26121 , n26122 ,
     n26123 , n26124 , n26125 , n26126 , n26127 , n26128 , n26129 , n26130 , n26131 , n26132 ,
     n26133 , n26134 , n26135 , n26136 , n26137 , n26138 , n26139 , n26140 , n26141 , n26142 ,
     n26143 , n26144 , n26145 , n26146 , n26147 , n26148 , n26149 , n26150 , n26151 , n26152 ,
     n26153 , n26154 , n26155 , n26156 , n26157 , n26158 , n26159 , n26160 , n26161 , n26162 ,
     n26163 , n26164 , n26165 , n26166 , n26167 , n26168 , n26169 , n26170 , n26171 , n26172 ,
     n26173 , n26174 , n26175 , n26176 , n26177 , n26178 , n26179 , n26180 , n26181 , n26182 ,
     n26183 , n26184 , n26185 , n26186 , n26187 , n26188 , n26189 , n26190 , n26191 , n26192 ,
     n26193 , n26194 , n26195 , n26196 , n26197 , n26198 , n26199 , n26200 , n26201 , n26202 ,
     n26203 , n26204 , n26205 , n26206 , n26207 , n26208 , n26209 , n26210 , n26211 , n26212 ,
     n26213 , n26214 , n26215 , n26216 , n26217 , n26218 , n26219 , n26220 , n26221 , n26222 ,
     n26223 , n26224 , n26225 , n26226 , n26227 , n26228 , n26229 , n26230 , n26231 , n26232 ,
     n26233 , n26234 , n26235 , n26236 , n26237 , n26238 , n26239 , n26240 , n26241 , n26242 ,
     n26243 , n26244 , n26245 , n26246 , n26247 , n26248 , n26249 , n26250 , n26251 , n26252 ,
     n26253 , n26254 , n26255 , n26256 , n26257 , n26258 , n26259 , n26260 , n26261 , n26262 ,
     n26263 , n26264 , n26265 , n26266 , n26267 , n26268 , n26269 , n26270 , n26271 , n26272 ,
     n26273 , n26274 , n26275 , n26276 , n26277 , n26278 , n26279 , n26280 , n26281 , n26282 ,
     n26283 , n26284 , n26285 , n26286 , n26287 , n26288 , n26289 , n26290 , n26291 , n26292 ,
     n26293 , n26294 , n26295 , n26296 , n26297 , n26298 , n26299 , n26300 , n26301 , n26302 ,
     n26303 , n26304 , n26305 , n26306 , n26307 , n26308 , n26309 , n26310 , n26311 , n26312 ,
     n26313 , n26314 , n26315 , n26316 , n26317 , n26318 , n26319 , n26320 , n26321 , n26322 ,
     n26323 , n26324 , n26325 , n26326 , n26327 , n26328 , n26329 , n26330 , n26331 , n26332 ,
     n26333 , n26334 , n26335 , n26336 , n26337 , n26338 , n26339 , n26340 , n26341 , n26342 ,
     n26343 , n26344 , n26345 , n26346 , n26347 , n26348 , n26349 , n26350 , n26351 , n26352 ,
     n26353 , n26354 , n26355 , n26356 , n26357 , n26358 , n26359 , n26360 , n26361 , n26362 ,
     n26363 , n26364 , n26365 , n26366 , n26367 , n26368 , n26369 , n26370 , n26371 , n26372 ,
     n26373 , n26374 , n26375 , n26376 , n26377 , n26378 , n26379 , n26380 , n26381 , n26382 ,
     n26383 , n26384 , n26385 , n26386 , n26387 , n26388 , n26389 , n26390 , n26391 , n26392 ,
     n26393 , n26394 , n26395 , n26396 , n26397 , n26398 , n26399 , n26400 , n26401 , n26402 ,
     n26403 , n26404 , n26405 , n26406 , n26407 , n26408 , n26409 , n26410 , n26411 , n26412 ,
     n26413 , n26414 , n26415 , n26416 , n26417 , n26418 , n26419 , n26420 , n26421 , n26422 ,
     n26423 , n26424 , n26425 , n26426 , n26427 , n26428 , n26429 , n26430 , n26431 , n26432 ,
     n26433 , n26434 , n26435 , n26436 , n26437 , n26438 , n26439 , n26440 , n26441 , n26442 ,
     n26443 , n26444 , n26445 , n26446 , n26447 , n26448 , n26449 , n26450 , n26451 , n26452 ,
     n26453 , n26454 , n26455 , n26456 , n26457 , n26458 , n26459 , n26460 , n26461 , n26462 ,
     n26463 , n26464 , n26465 , n26466 , n26467 , n26468 , n26469 , n26470 , n26471 , n26472 ,
     n26473 , n26474 , n26475 , n26476 , n26477 , n26478 , n26479 , n26480 , n26481 , n26482 ,
     n26483 , n26484 , n26485 , n26486 , n26487 , n26488 , n26489 , n26490 , n26491 , n26492 ,
     n26493 , n26494 , n26495 , n26496 , n26497 , n26498 , n26499 , n26500 , n26501 , n26502 ,
     n26503 , n26504 , n26505 , n26506 , n26507 , n26508 , n26509 , n26510 , n26511 , n26512 ,
     n26513 , n26514 , n26515 , n26516 , n26517 , n26518 , n26519 , n26520 , n26521 , n26522 ,
     n26523 , n26524 , n26525 , n26526 , n26527 , n26528 , n26529 , n26530 , n26531 , n26532 ,
     n26533 , n26534 , n26535 , n26536 , n26537 , n26538 , n26539 , n26540 , n26541 , n26542 ,
     n26543 , n26544 , n26545 , n26546 , n26547 , n26548 , n26549 , n26550 , n26551 , n26552 ,
     n26553 , n26554 , n26555 , n26556 , n26557 , n26558 , n26559 , n26560 , n26561 , n26562 ,
     n26563 , n26564 , n26565 , n26566 , n26567 , n26568 , n26569 , n26570 , n26571 , n26572 ,
     n26573 , n26574 , n26575 , n26576 , n26577 , n26578 , n26579 , n26580 , n26581 , n26582 ,
     n26583 , n26584 , n26585 , n26586 , n26587 , n26588 , n26589 , n26590 , n26591 , n26592 ,
     n26593 , n26594 , n26595 , n26596 , n26597 , n26598 , n26599 , n26600 , n26601 , n26602 ,
     n26603 , n26604 , n26605 , n26606 , n26607 , n26608 , n26609 , n26610 , n26611 , n26612 ,
     n26613 , n26614 , n26615 , n26616 , n26617 , n26618 , n26619 , n26620 , n26621 , n26622 ,
     n26623 , n26624 , n26625 , n26626 , n26627 , n26628 , n26629 , n26630 , n26631 , n26632 ,
     n26633 , n26634 , n26635 , n26636 , n26637 , n26638 , n26639 , n26640 , n26641 , n26642 ,
     n26643 , n26644 , n26645 , n26646 , n26647 , n26648 , n26649 , n26650 , n26651 , n26652 ,
     n26653 , n26654 , n26655 , n26656 , n26657 , n26658 , n26659 , n26660 , n26661 , n26662 ,
     n26663 , n26664 , n26665 , n26666 , n26667 , n26668 , n26669 , n26670 , n26671 , n26672 ,
     n26673 , n26674 , n26675 , n26676 , n26677 , n26678 , n26679 , n26680 , n26681 , n26682 ,
     n26683 , n26684 , n26685 , n26686 , n26687 , n26688 , n26689 , n26690 , n26691 , n26692 ,
     n26693 , n26694 , n26695 , n26696 , n26697 , n26698 , n26699 , n26700 , n26701 , n26702 ,
     n26703 , n26704 , n26705 , n26706 , n26707 , n26708 , n26709 , n26710 , n26711 , n26712 ,
     n26713 , n26714 , n26715 , n26716 , n26717 , n26718 , n26719 , n26720 , n26721 , n26722 ,
     n26723 , n26724 , n26725 , n26726 , n26727 , n26728 , n26729 , n26730 , n26731 , n26732 ,
     n26733 , n26734 , n26735 , n26736 , n26737 , n26738 , n26739 , n26740 , n26741 , n26742 ,
     n26743 , n26744 , n26745 , n26746 , n26747 , n26748 , n26749 , n26750 , n26751 , n26752 ,
     n26753 , n26754 , n26755 , n26756 , n26757 , n26758 , n26759 , n26760 , n26761 , n26762 ,
     n26763 , n26764 , n26765 , n26766 , n26767 , n26768 , n26769 , n26770 , n26771 , n26772 ,
     n26773 , n26774 , n26775 , n26776 , n26777 , n26778 , n26779 , n26780 , n26781 , n26782 ,
     n26783 , n26784 , n26785 , n26786 , n26787 , n26788 , n26789 , n26790 , n26791 , n26792 ,
     n26793 , n26794 , n26795 , n26796 , n26797 , n26798 , n26799 , n26800 , n26801 , n26802 ,
     n26803 , n26804 , n26805 , n26806 , n26807 , n26808 , n26809 , n26810 , n26811 , n26812 ,
     n26813 , n26814 , n26815 , n26816 , n26817 , n26818 , n26819 , n26820 , n26821 , n26822 ,
     n26823 , n26824 , n26825 , n26826 , n26827 , n26828 , n26829 , n26830 , n26831 , n26832 ,
     n26833 , n26834 , n26835 , n26836 , n26837 , n26838 , n26839 , n26840 , n26841 , n26842 ,
     n26843 , n26844 , n26845 , n26846 , n26847 , n26848 , n26849 , n26850 , n26851 , n26852 ,
     n26853 , n26854 , n26855 , n26856 , n26857 , n26858 , n26859 , n26860 , n26861 , n26862 ,
     n26863 , n26864 , n26865 , n26866 , n26867 , n26868 , n26869 , n26870 , n26871 , n26872 ,
     n26873 , n26874 , n26875 , n26876 , n26877 , n26878 , n26879 , n26880 , n26881 , n26882 ,
     n26883 , n26884 , n26885 , n26886 , n26887 , n26888 , n26889 , n26890 , n26891 , n26892 ,
     n26893 , n26894 , n26895 , n26896 , n26897 , n26898 , n26899 , n26900 , n26901 , n26902 ,
     n26903 , n26904 , n26905 , n26906 , n26907 , n26908 , n26909 , n26910 , n26911 , n26912 ,
     n26913 , n26914 , n26915 , n26916 , n26917 , n26918 , n26919 , n26920 , n26921 , n26922 ,
     n26923 , n26924 , n26925 , n26926 , n26927 , n26928 , n26929 , n26930 , n26931 , n26932 ,
     n26933 , n26934 , n26935 , n26936 , n26937 , n26938 , n26939 , n26940 , n26941 , n26942 ,
     n26943 , n26944 , n26945 , n26946 , n26947 , n26948 , n26949 , n26950 , n26951 , n26952 ,
     n26953 , n26954 , n26955 , n26956 , n26957 , n26958 , n26959 , n26960 , n26961 , n26962 ,
     n26963 , n26964 , n26965 , n26966 , n26967 , n26968 , n26969 , n26970 , n26971 , n26972 ,
     n26973 , n26974 , n26975 , n26976 , n26977 , n26978 , n26979 , n26980 , n26981 , n26982 ,
     n26983 , n26984 , n26985 , n26986 , n26987 , n26988 , n26989 , n26990 , n26991 , n26992 ,
     n26993 , n26994 , n26995 , n26996 , n26997 , n26998 , n26999 , n27000 , n27001 , n27002 ,
     n27003 , n27004 , n27005 , n27006 , n27007 , n27008 , n27009 , n27010 , n27011 , n27012 ,
     n27013 , n27014 , n27015 , n27016 , n27017 , n27018 , n27019 , n27020 , n27021 , n27022 ,
     n27023 , n27024 , n27025 , n27026 , n27027 , n27028 , n27029 , n27030 , n27031 , n27032 ,
     n27033 , n27034 , n27035 , n27036 , n27037 , n27038 , n27039 , n27040 , n27041 , n27042 ,
     n27043 , n27044 , n27045 , n27046 , n27047 , n27048 , n27049 , n27050 , n27051 , n27052 ,
     n27053 , n27054 , n27055 , n27056 , n27057 , n27058 , n27059 , n27060 , n27061 , n27062 ,
     n27063 , n27064 , n27065 , n27066 , n27067 , n27068 , n27069 , n27070 , n27071 , n27072 ,
     n27073 , n27074 , n27075 , n27076 , n27077 , n27078 , n27079 , n27080 , n27081 , n27082 ,
     n27083 , n27084 , n27085 , n27086 , n27087 , n27088 , n27089 , n27090 , n27091 , n27092 ,
     n27093 , n27094 , n27095 , n27096 , n27097 , n27098 , n27099 , n27100 , n27101 , n27102 ,
     n27103 , n27104 , n27105 , n27106 , n27107 , n27108 , n27109 , n27110 , n27111 , n27112 ,
     n27113 , n27114 , n27115 , n27116 , n27117 , n27118 , n27119 , n27120 , n27121 , n27122 ,
     n27123 , n27124 , n27125 , n27126 , n27127 , n27128 , n27129 , n27130 , n27131 , n27132 ,
     n27133 , n27134 , n27135 , n27136 , n27137 , n27138 , n27139 , n27140 , n27141 , n27142 ,
     n27143 , n27144 , n27145 , n27146 , n27147 , n27148 , n27149 , n27150 , n27151 , n27152 ,
     n27153 , n27154 , n27155 , n27156 , n27157 , n27158 , n27159 , n27160 , n27161 , n27162 ,
     n27163 , n27164 , n27165 , n27166 , n27167 , n27168 , n27169 , n27170 , n27171 , n27172 ,
     n27173 , n27174 , n27175 , n27176 , n27177 , n27178 , n27179 , n27180 , n27181 , n27182 ,
     n27183 , n27184 , n27185 , n27186 , n27187 , n27188 , n27189 , n27190 , n27191 , n27192 ,
     n27193 , n27194 , n27195 , n27196 , n27197 , n27198 , n27199 , n27200 , n27201 , n27202 ,
     n27203 , n27204 , n27205 , n27206 , n27207 , n27208 , n27209 , n27210 , n27211 , n27212 ,
     n27213 , n27214 , n27215 , n27216 , n27217 , n27218 , n27219 , n27220 , n27221 , n27222 ,
     n27223 , n27224 , n27225 , n27226 , n27227 , n27228 , n27229 , n27230 , n27231 , n27232 ,
     n27233 , n27234 , n27235 , n27236 , n27237 , n27238 , n27239 , n27240 , n27241 , n27242 ,
     n27243 , n27244 , n27245 , n27246 , n27247 , n27248 , n27249 , n27250 , n27251 , n27252 ,
     n27253 , n27254 , n27255 , n27256 , n27257 , n27258 , n27259 , n27260 , n27261 , n27262 ,
     n27263 , n27264 , n27265 , n27266 , n27267 , n27268 , n27269 , n27270 , n27271 , n27272 ,
     n27273 , n27274 , n27275 , n27276 , n27277 , n27278 , n27279 , n27280 , n27281 , n27282 ,
     n27283 , n27284 , n27285 , n27286 , n27287 , n27288 , n27289 , n27290 , n27291 , n27292 ,
     n27293 , n27294 , n27295 , n27296 , n27297 , n27298 , n27299 , n27300 , n27301 , n27302 ,
     n27303 , n27304 , n27305 , n27306 , n27307 , n27308 , n27309 , n27310 , n27311 , n27312 ,
     n27313 , n27314 , n27315 , n27316 , n27317 , n27318 , n27319 , n27320 , n27321 , n27322 ,
     n27323 , n27324 , n27325 , n27326 , n27327 , n27328 , n27329 , n27330 , n27331 , n27332 ,
     n27333 , n27334 , n27335 , n27336 , n27337 , n27338 , n27339 , n27340 , n27341 , n27342 ,
     n27343 , n27344 , n27345 , n27346 , n27347 , n27348 , n27349 , n27350 , n27351 , n27352 ,
     n27353 , n27354 , n27355 , n27356 , n27357 , n27358 , n27359 , n27360 , n27361 , n27362 ,
     n27363 , n27364 , n27365 , n27366 , n27367 , n27368 , n27369 , n27370 , n27371 , n27372 ,
     n27373 , n27374 , n27375 , n27376 , n27377 , n27378 , n27379 , n27380 , n27381 , n27382 ,
     n27383 , n27384 , n27385 , n27386 , n27387 , n27388 , n27389 , n27390 , n27391 , n27392 ,
     n27393 , n27394 , n27395 , n27396 , n27397 , n27398 , n27399 , n27400 , n27401 , n27402 ,
     n27403 , n27404 , n27405 , n27406 , n27407 , n27408 , n27409 , n27410 , n27411 , n27412 ,
     n27413 , n27414 , n27415 , n27416 , n27417 , n27418 , n27419 , n27420 , n27421 , n27422 ,
     n27423 , n27424 , n27425 , n27426 , n27427 , n27428 , n27429 , n27430 , n27431 , n27432 ,
     n27433 , n27434 , n27435 , n27436 , n27437 , n27438 , n27439 , n27440 , n27441 , n27442 ,
     n27443 , n27444 , n27445 , n27446 , n27447 , n27448 , n27449 , n27450 , n27451 , n27452 ,
     n27453 , n27454 , n27455 , n27456 , n27457 , n27458 , n27459 , n27460 , n27461 , n27462 ,
     n27463 , n27464 , n27465 , n27466 , n27467 , n27468 , n27469 , n27470 , n27471 , n27472 ,
     n27473 , n27474 , n27475 , n27476 , n27477 , n27478 , n27479 , n27480 , n27481 , n27482 ,
     n27483 , n27484 , n27485 , n27486 , n27487 , n27488 , n27489 , n27490 , n27491 , n27492 ,
     n27493 , n27494 , n27495 , n27496 , n27497 , n27498 , n27499 , n27500 , n27501 , n27502 ,
     n27503 , n27504 , n27505 , n27506 , n27507 , n27508 , n27509 , n27510 , n27511 , n27512 ,
     n27513 , n27514 , n27515 , n27516 , n27517 , n27518 , n27519 , n27520 , n27521 , n27522 ,
     n27523 , n27524 , n27525 , n27526 , n27527 , n27528 , n27529 , n27530 , n27531 , n27532 ,
     n27533 , n27534 , n27535 , n27536 , n27537 , n27538 , n27539 , n27540 , n27541 , n27542 ,
     n27543 , n27544 , n27545 , n27546 , n27547 , n27548 , n27549 , n27550 , n27551 , n27552 ,
     n27553 , n27554 , n27555 , n27556 , n27557 , n27558 , n27559 , n27560 , n27561 , n27562 ,
     n27563 , n27564 , n27565 , n27566 , n27567 , n27568 , n27569 , n27570 , n27571 , n27572 ,
     n27573 , n27574 , n27575 , n27576 , n27577 , n27578 , n27579 , n27580 , n27581 , n27582 ,
     n27583 , n27584 , n27585 , n27586 , n27587 , n27588 , n27589 , n27590 , n27591 , n27592 ,
     n27593 , n27594 , n27595 , n27596 , n27597 , n27598 , n27599 , n27600 , n27601 , n27602 ,
     n27603 , n27604 , n27605 , n27606 , n27607 , n27608 , n27609 , n27610 , n27611 , n27612 ,
     n27613 , n27614 , n27615 , n27616 , n27617 , n27618 , n27619 , n27620 , n27621 , n27622 ,
     n27623 , n27624 , n27625 , n27626 , n27627 , n27628 , n27629 , n27630 , n27631 , n27632 ,
     n27633 , n27634 , n27635 , n27636 , n27637 , n27638 , n27639 , n27640 , n27641 , n27642 ,
     n27643 , n27644 , n27645 , n27646 , n27647 , n27648 , n27649 , n27650 , n27651 , n27652 ,
     n27653 , n27654 , n27655 , n27656 , n27657 , n27658 , n27659 , n27660 , n27661 , n27662 ,
     n27663 , n27664 , n27665 , n27666 , n27667 , n27668 , n27669 , n27670 , n27671 , n27672 ,
     n27673 , n27674 , n27675 , n27676 , n27677 , n27678 , n27679 , n27680 , n27681 , n27682 ,
     n27683 , n27684 , n27685 , n27686 , n27687 , n27688 , n27689 , n27690 , n27691 , n27692 ,
     n27693 , n27694 , n27695 , n27696 , n27697 , n27698 , n27699 , n27700 , n27701 , n27702 ,
     n27703 , n27704 , n27705 , n27706 , n27707 , n27708 , n27709 , n27710 , n27711 , n27712 ,
     n27713 , n27714 , n27715 , n27716 , n27717 , n27718 , n27719 , n27720 , n27721 , n27722 ,
     n27723 , n27724 , n27725 , n27726 , n27727 , n27728 , n27729 , n27730 , n27731 , n27732 ,
     n27733 , n27734 , n27735 , n27736 , n27737 , n27738 , n27739 , n27740 , n27741 , n27742 ,
     n27743 , n27744 , n27745 , n27746 , n27747 , n27748 , n27749 , n27750 , n27751 , n27752 ,
     n27753 , n27754 , n27755 , n27756 , n27757 , n27758 , n27759 , n27760 , n27761 , n27762 ,
     n27763 , n27764 , n27765 , n27766 , n27767 , n27768 , n27769 , n27770 , n27771 , n27772 ,
     n27773 , n27774 , n27775 , n27776 , n27777 , n27778 , n27779 , n27780 , n27781 , n27782 ,
     n27783 , n27784 , n27785 , n27786 , n27787 , n27788 , n27789 , n27790 , n27791 , n27792 ,
     n27793 , n27794 , n27795 , n27796 , n27797 , n27798 , n27799 , n27800 , n27801 , n27802 ,
     n27803 , n27804 , n27805 , n27806 , n27807 , n27808 , n27809 , n27810 , n27811 , n27812 ,
     n27813 , n27814 , n27815 , n27816 , n27817 , n27818 , n27819 , n27820 , n27821 , n27822 ,
     n27823 , n27824 , n27825 , n27826 , n27827 , n27828 , n27829 , n27830 , n27831 , n27832 ,
     n27833 , n27834 , n27835 , n27836 , n27837 , n27838 , n27839 , n27840 , n27841 , n27842 ,
     n27843 , n27844 , n27845 , n27846 , n27847 , n27848 , n27849 , n27850 , n27851 , n27852 ,
     n27853 , n27854 , n27855 , n27856 , n27857 , n27858 , n27859 , n27860 , n27861 , n27862 ,
     n27863 , n27864 , n27865 , n27866 , n27867 , n27868 , n27869 , n27870 , n27871 , n27872 ,
     n27873 , n27874 , n27875 , n27876 , n27877 , n27878 , n27879 , n27880 , n27881 , n27882 ,
     n27883 , n27884 , n27885 , n27886 , n27887 , n27888 , n27889 , n27890 , n27891 , n27892 ,
     n27893 , n27894 , n27895 , n27896 , n27897 , n27898 , n27899 , n27900 , n27901 , n27902 ,
     n27903 , n27904 , n27905 , n27906 , n27907 , n27908 , n27909 , n27910 , n27911 , n27912 ,
     n27913 , n27914 , n27915 , n27916 , n27917 , n27918 , n27919 , n27920 , n27921 , n27922 ,
     n27923 , n27924 , n27925 , n27926 , n27927 , n27928 , n27929 , n27930 , n27931 , n27932 ,
     n27933 , n27934 , n27935 , n27936 , n27937 , n27938 , n27939 , n27940 , n27941 , n27942 ,
     n27943 , n27944 , n27945 , n27946 , n27947 , n27948 , n27949 , n27950 , n27951 , n27952 ,
     n27953 , n27954 , n27955 , n27956 , n27957 , n27958 , n27959 , n27960 , n27961 , n27962 ,
     n27963 , n27964 , n27965 , n27966 , n27967 , n27968 , n27969 , n27970 , n27971 , n27972 ,
     n27973 , n27974 , n27975 , n27976 , n27977 , n27978 , n27979 , n27980 , n27981 , n27982 ,
     n27983 , n27984 , n27985 , n27986 , n27987 , n27988 , n27989 , n27990 , n27991 , n27992 ,
     n27993 , n27994 , n27995 , n27996 , n27997 , n27998 , n27999 , n28000 , n28001 , n28002 ,
     n28003 , n28004 , n28005 , n28006 , n28007 , n28008 , n28009 , n28010 , n28011 , n28012 ,
     n28013 , n28014 , n28015 , n28016 , n28017 , n28018 , n28019 , n28020 , n28021 , n28022 ,
     n28023 , n28024 , n28025 , n28026 , n28027 , n28028 , n28029 , n28030 , n28031 , n28032 ,
     n28033 , n28034 , n28035 , n28036 , n28037 , n28038 , n28039 , n28040 , n28041 , n28042 ,
     n28043 , n28044 , n28045 , n28046 , n28047 , n28048 , n28049 , n28050 , n28051 , n28052 ,
     n28053 , n28054 , n28055 , n28056 , n28057 , n28058 , n28059 , n28060 , n28061 , n28062 ,
     n28063 , n28064 , n28065 , n28066 , n28067 , n28068 , n28069 , n28070 , n28071 , n28072 ,
     n28073 , n28074 , n28075 , n28076 , n28077 , n28078 , n28079 , n28080 , n28081 , n28082 ,
     n28083 , n28084 , n28085 , n28086 , n28087 , n28088 , n28089 , n28090 , n28091 , n28092 ,
     n28093 , n28094 , n28095 , n28096 , n28097 , n28098 , n28099 , n28100 , n28101 , n28102 ,
     n28103 , n28104 , n28105 , n28106 , n28107 , n28108 , n28109 , n28110 , n28111 , n28112 ,
     n28113 , n28114 , n28115 , n28116 , n28117 , n28118 , n28119 , n28120 , n28121 , n28122 ,
     n28123 , n28124 , n28125 , n28126 , n28127 , n28128 , n28129 , n28130 , n28131 , n28132 ,
     n28133 , n28134 , n28135 , n28136 , n28137 , n28138 , n28139 , n28140 , n28141 , n28142 ,
     n28143 , n28144 , n28145 , n28146 , n28147 , n28148 , n28149 , n28150 , n28151 , n28152 ,
     n28153 , n28154 , n28155 , n28156 , n28157 , n28158 , n28159 , n28160 , n28161 , n28162 ,
     n28163 , n28164 , n28165 , n28166 , n28167 , n28168 , n28169 , n28170 , n28171 , n28172 ,
     n28173 , n28174 , n28175 , n28176 , n28177 , n28178 , n28179 , n28180 , n28181 , n28182 ,
     n28183 , n28184 , n28185 , n28186 , n28187 , n28188 , n28189 , n28190 , n28191 , n28192 ,
     n28193 , n28194 , n28195 , n28196 , n28197 , n28198 , n28199 , n28200 , n28201 , n28202 ,
     n28203 , n28204 , n28205 , n28206 , n28207 , n28208 , n28209 , n28210 , n28211 , n28212 ,
     n28213 , n28214 , n28215 , n28216 , n28217 , n28218 , n28219 , n28220 , n28221 , n28222 ,
     n28223 , n28224 , n28225 , n28226 , n28227 , n28228 , n28229 , n28230 , n28231 , n28232 ,
     n28233 , n28234 , n28235 , n28236 , n28237 , n28238 , n28239 , n28240 , n28241 , n28242 ,
     n28243 , n28244 , n28245 , n28246 , n28247 , n28248 , n28249 , n28250 , n28251 , n28252 ,
     n28253 , n28254 , n28255 , n28256 , n28257 , n28258 , n28259 , n28260 , n28261 , n28262 ,
     n28263 , n28264 , n28265 , n28266 , n28267 , n28268 , n28269 , n28270 , n28271 , n28272 ,
     n28273 , n28274 , n28275 , n28276 , n28277 , n28278 , n28279 , n28280 , n28281 , n28282 ,
     n28283 , n28284 , n28285 , n28286 , n28287 , n28288 , n28289 , n28290 , n28291 , n28292 ,
     n28293 , n28294 , n28295 , n28296 , n28297 , n28298 , n28299 , n28300 , n28301 , n28302 ,
     n28303 , n28304 , n28305 , n28306 , n28307 , n28308 , n28309 , n28310 , n28311 , n28312 ,
     n28313 , n28314 , n28315 , n28316 , n28317 , n28318 , n28319 , n28320 , n28321 , n28322 ,
     n28323 , n28324 , n28325 , n28326 , n28327 , n28328 , n28329 , n28330 , n28331 , n28332 ,
     n28333 , n28334 , n28335 , n28336 , n28337 , n28338 , n28339 , n28340 , n28341 , n28342 ,
     n28343 , n28344 , n28345 , n28346 , n28347 , n28348 , n28349 , n28350 , n28351 , n28352 ,
     n28353 , n28354 , n28355 , n28356 , n28357 , n28358 , n28359 , n28360 , n28361 , n28362 ,
     n28363 , n28364 , n28365 , n28366 , n28367 , n28368 , n28369 , n28370 , n28371 , n28372 ,
     n28373 , n28374 , n28375 , n28376 , n28377 , n28378 , n28379 , n28380 , n28381 , n28382 ,
     n28383 , n28384 , n28385 , n28386 , n28387 , n28388 , n28389 , n28390 , n28391 , n28392 ,
     n28393 , n28394 , n28395 , n28396 , n28397 , n28398 , n28399 , n28400 , n28401 , n28402 ,
     n28403 , n28404 , n28405 , n28406 , n28407 , n28408 , n28409 , n28410 , n28411 , n28412 ,
     n28413 , n28414 , n28415 , n28416 , n28417 , n28418 , n28419 , n28420 , n28421 , n28422 ,
     n28423 , n28424 , n28425 , n28426 , n28427 , n28428 , n28429 , n28430 , n28431 , n28432 ,
     n28433 , n28434 , n28435 , n28436 , n28437 , n28438 , n28439 , n28440 , n28441 , n28442 ,
     n28443 , n28444 , n28445 , n28446 , n28447 , n28448 , n28449 , n28450 , n28451 , n28452 ,
     n28453 , n28454 , n28455 , n28456 , n28457 , n28458 , n28459 , n28460 , n28461 , n28462 ,
     n28463 , n28464 , n28465 , n28466 , n28467 , n28468 , n28469 , n28470 , n28471 , n28472 ,
     n28473 , n28474 , n28475 , n28476 , n28477 , n28478 , n28479 , n28480 , n28481 , n28482 ,
     n28483 , n28484 , n28485 , n28486 , n28487 , n28488 , n28489 , n28490 , n28491 , n28492 ,
     n28493 , n28494 , n28495 , n28496 , n28497 , n28498 , n28499 , n28500 , n28501 , n28502 ,
     n28503 , n28504 , n28505 , n28506 , n28507 , n28508 , n28509 , n28510 , n28511 , n28512 ,
     n28513 , n28514 , n28515 , n28516 , n28517 , n28518 , n28519 , n28520 , n28521 , n28522 ,
     n28523 , n28524 , n28525 , n28526 , n28527 , n28528 , n28529 , n28530 , n28531 , n28532 ,
     n28533 , n28534 , n28535 , n28536 , n28537 , n28538 , n28539 , n28540 , n28541 , n28542 ,
     n28543 , n28544 , n28545 , n28546 , n28547 , n28548 , n28549 , n28550 , n28551 , n28552 ,
     n28553 , n28554 , n28555 , n28556 , n28557 , n28558 , n28559 , n28560 , n28561 , n28562 ,
     n28563 , n28564 , n28565 , n28566 , n28567 , n28568 , n28569 , n28570 , n28571 , n28572 ,
     n28573 , n28574 , n28575 , n28576 , n28577 , n28578 , n28579 , n28580 , n28581 , n28582 ,
     n28583 , n28584 , n28585 , n28586 , n28587 , n28588 , n28589 , n28590 , n28591 , n28592 ,
     n28593 , n28594 , n28595 , n28596 , n28597 , n28598 , n28599 , n28600 , n28601 , n28602 ,
     n28603 , n28604 , n28605 , n28606 , n28607 , n28608 , n28609 , n28610 , n28611 , n28612 ,
     n28613 , n28614 , n28615 , n28616 , n28617 , n28618 , n28619 , n28620 , n28621 , n28622 ,
     n28623 , n28624 , n28625 , n28626 , n28627 , n28628 , n28629 , n28630 , n28631 , n28632 ,
     n28633 , n28634 , n28635 , n28636 , n28637 , n28638 , n28639 , n28640 , n28641 , n28642 ,
     n28643 , n28644 , n28645 , n28646 , n28647 , n28648 , n28649 , n28650 , n28651 , n28652 ,
     n28653 , n28654 , n28655 , n28656 , n28657 , n28658 , n28659 , n28660 , n28661 , n28662 ,
     n28663 , n28664 , n28665 , n28666 , n28667 , n28668 , n28669 , n28670 , n28671 , n28672 ,
     n28673 , n28674 , n28675 , n28676 , n28677 , n28678 , n28679 , n28680 , n28681 , n28682 ,
     n28683 , n28684 , n28685 , n28686 , n28687 , n28688 , n28689 , n28690 , n28691 , n28692 ,
     n28693 , n28694 , n28695 , n28696 , n28697 , n28698 , n28699 , n28700 , n28701 , n28702 ,
     n28703 , n28704 , n28705 , n28706 , n28707 , n28708 , n28709 , n28710 , n28711 , n28712 ,
     n28713 , n28714 , n28715 , n28716 , n28717 , n28718 , n28719 , n28720 , n28721 , n28722 ,
     n28723 , n28724 , n28725 , n28726 , n28727 , n28728 , n28729 , n28730 , n28731 , n28732 ,
     n28733 , n28734 , n28735 , n28736 , n28737 , n28738 , n28739 , n28740 , n28741 , n28742 ,
     n28743 , n28744 , n28745 , n28746 , n28747 , n28748 , n28749 , n28750 , n28751 , n28752 ,
     n28753 , n28754 , n28755 , n28756 , n28757 , n28758 , n28759 , n28760 , n28761 , n28762 ,
     n28763 , n28764 , n28765 , n28766 , n28767 , n28768 , n28769 , n28770 , n28771 , n28772 ,
     n28773 , n28774 , n28775 , n28776 , n28777 , n28778 , n28779 , n28780 , n28781 , n28782 ,
     n28783 , n28784 , n28785 , n28786 , n28787 , n28788 , n28789 , n28790 , n28791 , n28792 ,
     n28793 , n28794 , n28795 , n28796 , n28797 , n28798 , n28799 , n28800 , n28801 , n28802 ,
     n28803 , n28804 , n28805 , n28806 , n28807 , n28808 , n28809 , n28810 , n28811 , n28812 ,
     n28813 , n28814 , n28815 , n28816 , n28817 , n28818 , n28819 , n28820 , n28821 , n28822 ,
     n28823 , n28824 , n28825 , n28826 , n28827 , n28828 , n28829 , n28830 , n28831 , n28832 ,
     n28833 , n28834 , n28835 , n28836 , n28837 , n28838 , n28839 , n28840 , n28841 , n28842 ,
     n28843 , n28844 , n28845 , n28846 , n28847 , n28848 , n28849 , n28850 , n28851 , n28852 ,
     n28853 , n28854 , n28855 , n28856 , n28857 , n28858 , n28859 , n28860 , n28861 , n28862 ,
     n28863 , n28864 , n28865 , n28866 , n28867 , n28868 , n28869 , n28870 , n28871 , n28872 ,
     n28873 , n28874 , n28875 , n28876 , n28877 , n28878 , n28879 , n28880 , n28881 , n28882 ,
     n28883 , n28884 , n28885 , n28886 , n28887 , n28888 , n28889 , n28890 , n28891 , n28892 ,
     n28893 , n28894 , n28895 , n28896 , n28897 , n28898 , n28899 , n28900 , n28901 , n28902 ,
     n28903 , n28904 , n28905 , n28906 , n28907 , n28908 , n28909 , n28910 , n28911 , n28912 ,
     n28913 , n28914 , n28915 , n28916 , n28917 , n28918 , n28919 , n28920 , n28921 , n28922 ,
     n28923 , n28924 , n28925 , n28926 , n28927 , n28928 , n28929 , n28930 , n28931 , n28932 ,
     n28933 , n28934 , n28935 , n28936 , n28937 , n28938 , n28939 , n28940 , n28941 , n28942 ,
     n28943 , n28944 , n28945 , n28946 , n28947 , n28948 , n28949 , n28950 , n28951 , n28952 ,
     n28953 , n28954 , n28955 , n28956 , n28957 , n28958 , n28959 , n28960 , n28961 , n28962 ,
     n28963 , n28964 , n28965 , n28966 , n28967 , n28968 , n28969 , n28970 , n28971 , n28972 ,
     n28973 , n28974 , n28975 , n28976 , n28977 , n28978 , n28979 , n28980 , n28981 , n28982 ,
     n28983 , n28984 , n28985 , n28986 , n28987 , n28988 , n28989 , n28990 , n28991 , n28992 ,
     n28993 , n28994 , n28995 , n28996 , n28997 , n28998 , n28999 , n29000 , n29001 , n29002 ,
     n29003 , n29004 , n29005 , n29006 , n29007 , n29008 , n29009 , n29010 , n29011 , n29012 ,
     n29013 , n29014 , n29015 , n29016 , n29017 , n29018 , n29019 , n29020 , n29021 , n29022 ,
     n29023 , n29024 , n29025 , n29026 , n29027 , n29028 , n29029 , n29030 , n29031 , n29032 ,
     n29033 , n29034 , n29035 , n29036 , n29037 , n29038 , n29039 , n29040 , n29041 , n29042 ,
     n29043 , n29044 , n29045 , n29046 , n29047 , n29048 , n29049 , n29050 , n29051 , n29052 ,
     n29053 , n29054 , n29055 , n29056 , n29057 , n29058 , n29059 , n29060 , n29061 , n29062 ,
     n29063 , n29064 , n29065 , n29066 , n29067 , n29068 , n29069 , n29070 , n29071 , n29072 ,
     n29073 , n29074 , n29075 , n29076 , n29077 , n29078 , n29079 , n29080 , n29081 , n29082 ,
     n29083 , n29084 , n29085 , n29086 , n29087 , n29088 , n29089 , n29090 , n29091 , n29092 ,
     n29093 , n29094 , n29095 , n29096 , n29097 , n29098 , n29099 , n29100 , n29101 , n29102 ,
     n29103 , n29104 , n29105 , n29106 , n29107 , n29108 , n29109 , n29110 , n29111 , n29112 ,
     n29113 , n29114 , n29115 , n29116 , n29117 , n29118 , n29119 , n29120 , n29121 , n29122 ,
     n29123 , n29124 , n29125 , n29126 , n29127 , n29128 , n29129 , n29130 , n29131 , n29132 ,
     n29133 , n29134 , n29135 , n29136 , n29137 , n29138 , n29139 , n29140 , n29141 , n29142 ,
     n29143 , n29144 , n29145 , n29146 , n29147 , n29148 , n29149 , n29150 , n29151 , n29152 ,
     n29153 , n29154 , n29155 , n29156 , n29157 , n29158 , n29159 , n29160 , n29161 , n29162 ,
     n29163 , n29164 , n29165 , n29166 , n29167 , n29168 , n29169 , n29170 , n29171 , n29172 ,
     n29173 , n29174 , n29175 , n29176 , n29177 , n29178 , n29179 , n29180 , n29181 , n29182 ,
     n29183 , n29184 , n29185 , n29186 , n29187 , n29188 , n29189 , n29190 , n29191 , n29192 ,
     n29193 , n29194 , n29195 , n29196 , n29197 , n29198 , n29199 , n29200 , n29201 , n29202 ,
     n29203 , n29204 , n29205 , n29206 , n29207 , n29208 , n29209 , n29210 , n29211 , n29212 ,
     n29213 , n29214 , n29215 , n29216 , n29217 , n29218 , n29219 , n29220 , n29221 , n29222 ,
     n29223 , n29224 , n29225 , n29226 , n29227 , n29228 , n29229 , n29230 , n29231 , n29232 ,
     n29233 , n29234 , n29235 , n29236 , n29237 , n29238 , n29239 , n29240 , n29241 , n29242 ,
     n29243 , n29244 , n29245 , n29246 , n29247 , n29248 , n29249 , n29250 , n29251 , n29252 ,
     n29253 , n29254 , n29255 , n29256 , n29257 , n29258 , n29259 , n29260 , n29261 , n29262 ,
     n29263 , n29264 , n29265 , n29266 , n29267 , n29268 , n29269 , n29270 , n29271 , n29272 ,
     n29273 , n29274 , n29275 , n29276 , n29277 , n29278 , n29279 , n29280 , n29281 , n29282 ,
     n29283 , n29284 , n29285 , n29286 , n29287 , n29288 , n29289 , n29290 , n29291 , n29292 ,
     n29293 , n29294 , n29295 , n29296 , n29297 , n29298 , n29299 , n29300 , n29301 , n29302 ,
     n29303 , n29304 , n29305 , n29306 , n29307 , n29308 , n29309 , n29310 , n29311 , n29312 ,
     n29313 , n29314 , n29315 , n29316 , n29317 , n29318 , n29319 , n29320 , n29321 , n29322 ,
     n29323 , n29324 , n29325 , n29326 , n29327 , n29328 , n29329 , n29330 , n29331 , n29332 ,
     n29333 , n29334 , n29335 , n29336 , n29337 , n29338 , n29339 , n29340 , n29341 , n29342 ,
     n29343 , n29344 , n29345 , n29346 , n29347 , n29348 , n29349 , n29350 , n29351 , n29352 ,
     n29353 , n29354 , n29355 , n29356 , n29357 , n29358 , n29359 , n29360 , n29361 , n29362 ,
     n29363 , n29364 , n29365 , n29366 , n29367 , n29368 , n29369 , n29370 , n29371 , n29372 ,
     n29373 , n29374 , n29375 , n29376 , n29377 , n29378 , n29379 , n29380 , n29381 , n29382 ,
     n29383 , n29384 , n29385 , n29386 , n29387 , n29388 , n29389 , n29390 , n29391 , n29392 ,
     n29393 , n29394 , n29395 , n29396 , n29397 , n29398 , n29399 , n29400 , n29401 , n29402 ,
     n29403 , n29404 , n29405 , n29406 , n29407 , n29408 , n29409 , n29410 , n29411 , n29412 ,
     n29413 , n29414 , n29415 , n29416 , n29417 , n29418 , n29419 , n29420 , n29421 , n29422 ,
     n29423 , n29424 , n29425 , n29426 , n29427 , n29428 , n29429 , n29430 , n29431 , n29432 ,
     n29433 , n29434 , n29435 , n29436 , n29437 , n29438 , n29439 , n29440 , n29441 , n29442 ,
     n29443 , n29444 , n29445 , n29446 , n29447 , n29448 , n29449 , n29450 , n29451 , n29452 ,
     n29453 , n29454 , n29455 , n29456 , n29457 , n29458 , n29459 , n29460 , n29461 , n29462 ,
     n29463 , n29464 , n29465 , n29466 , n29467 , n29468 , n29469 , n29470 , n29471 , n29472 ,
     n29473 , n29474 , n29475 , n29476 , n29477 , n29478 , n29479 , n29480 , n29481 , n29482 ,
     n29483 , n29484 , n29485 , n29486 , n29487 , n29488 , n29489 , n29490 , n29491 , n29492 ,
     n29493 , n29494 , n29495 , n29496 , n29497 , n29498 , n29499 , n29500 , n29501 , n29502 ,
     n29503 , n29504 , n29505 , n29506 , n29507 , n29508 , n29509 , n29510 , n29511 , n29512 ,
     n29513 , n29514 , n29515 , n29516 , n29517 , n29518 , n29519 , n29520 , n29521 , n29522 ,
     n29523 , n29524 , n29525 , n29526 , n29527 , n29528 , n29529 , n29530 , n29531 , n29532 ,
     n29533 , n29534 , n29535 , n29536 , n29537 , n29538 , n29539 , n29540 , n29541 , n29542 ,
     n29543 , n29544 , n29545 , n29546 , n29547 , n29548 , n29549 , n29550 , n29551 , n29552 ,
     n29553 , n29554 , n29555 , n29556 , n29557 , n29558 , n29559 , n29560 , n29561 , n29562 ,
     n29563 , n29564 , n29565 , n29566 , n29567 , n29568 , n29569 , n29570 , n29571 , n29572 ,
     n29573 , n29574 , n29575 , n29576 , n29577 , n29578 , n29579 , n29580 , n29581 , n29582 ,
     n29583 , n29584 , n29585 , n29586 , n29587 , n29588 , n29589 , n29590 , n29591 , n29592 ,
     n29593 , n29594 , n29595 , n29596 , n29597 , n29598 , n29599 , n29600 , n29601 , n29602 ,
     n29603 , n29604 , n29605 , n29606 , n29607 , n29608 , n29609 , n29610 , n29611 , n29612 ,
     n29613 , n29614 , n29615 , n29616 , n29617 , n29618 , n29619 , n29620 , n29621 , n29622 ,
     n29623 , n29624 , n29625 , n29626 , n29627 , n29628 , n29629 , n29630 , n29631 , n29632 ,
     n29633 , n29634 , n29635 , n29636 , n29637 , n29638 , n29639 , n29640 , n29641 , n29642 ,
     n29643 , n29644 , n29645 , n29646 , n29647 , n29648 , n29649 , n29650 , n29651 , n29652 ,
     n29653 , n29654 , n29655 , n29656 , n29657 , n29658 , n29659 , n29660 , n29661 , n29662 ,
     n29663 , n29664 , n29665 , n29666 , n29667 , n29668 , n29669 , n29670 , n29671 , n29672 ,
     n29673 , n29674 , n29675 , n29676 , n29677 , n29678 , n29679 , n29680 , n29681 , n29682 ,
     n29683 , n29684 , n29685 , n29686 , n29687 , n29688 , n29689 , n29690 , n29691 , n29692 ,
     n29693 , n29694 , n29695 , n29696 , n29697 , n29698 , n29699 , n29700 , n29701 , n29702 ,
     n29703 , n29704 , n29705 , n29706 , n29707 , n29708 , n29709 , n29710 , n29711 , n29712 ,
     n29713 , n29714 , n29715 , n29716 , n29717 , n29718 , n29719 , n29720 , n29721 , n29722 ,
     n29723 , n29724 , n29725 , n29726 , n29727 , n29728 , n29729 , n29730 , n29731 , n29732 ,
     n29733 , n29734 , n29735 , n29736 , n29737 , n29738 , n29739 , n29740 , n29741 , n29742 ,
     n29743 , n29744 , n29745 , n29746 , n29747 , n29748 , n29749 , n29750 , n29751 , n29752 ,
     n29753 , n29754 , n29755 , n29756 , n29757 , n29758 , n29759 , n29760 , n29761 , n29762 ,
     n29763 , n29764 , n29765 , n29766 , n29767 , n29768 , n29769 , n29770 , n29771 , n29772 ,
     n29773 , n29774 , n29775 , n29776 , n29777 , n29778 , n29779 , n29780 , n29781 , n29782 ,
     n29783 , n29784 , n29785 , n29786 , n29787 , n29788 , n29789 , n29790 , n29791 , n29792 ,
     n29793 , n29794 , n29795 , n29796 , n29797 , n29798 , n29799 , n29800 , n29801 , n29802 ,
     n29803 , n29804 , n29805 , n29806 , n29807 , n29808 , n29809 , n29810 , n29811 , n29812 ,
     n29813 , n29814 , n29815 , n29816 , n29817 , n29818 , n29819 , n29820 , n29821 , n29822 ,
     n29823 , n29824 , n29825 , n29826 , n29827 , n29828 , n29829 , n29830 , n29831 , n29832 ,
     n29833 , n29834 , n29835 , n29836 , n29837 , n29838 , n29839 , n29840 , n29841 , n29842 ,
     n29843 , n29844 , n29845 , n29846 , n29847 , n29848 , n29849 , n29850 , n29851 , n29852 ,
     n29853 , n29854 , n29855 , n29856 , n29857 , n29858 , n29859 , n29860 , n29861 , n29862 ,
     n29863 , n29864 , n29865 , n29866 , n29867 , n29868 , n29869 , n29870 , n29871 , n29872 ,
     n29873 , n29874 , n29875 , n29876 , n29877 , n29878 , n29879 , n29880 , n29881 , n29882 ,
     n29883 , n29884 , n29885 , n29886 , n29887 , n29888 , n29889 , n29890 , n29891 , n29892 ,
     n29893 , n29894 , n29895 , n29896 , n29897 , n29898 , n29899 , n29900 , n29901 , n29902 ,
     n29903 , n29904 , n29905 , n29906 , n29907 , n29908 , n29909 , n29910 , n29911 , n29912 ,
     n29913 , n29914 , n29915 , n29916 , n29917 , n29918 , n29919 , n29920 , n29921 , n29922 ,
     n29923 , n29924 , n29925 , n29926 , n29927 , n29928 , n29929 , n29930 , n29931 , n29932 ,
     n29933 , n29934 , n29935 , n29936 , n29937 , n29938 , n29939 , n29940 , n29941 , n29942 ,
     n29943 , n29944 , n29945 , n29946 , n29947 , n29948 , n29949 , n29950 , n29951 , n29952 ,
     n29953 , n29954 , n29955 , n29956 , n29957 , n29958 , n29959 , n29960 , n29961 , n29962 ,
     n29963 , n29964 , n29965 , n29966 , n29967 , n29968 , n29969 , n29970 , n29971 , n29972 ,
     n29973 , n29974 , n29975 , n29976 , n29977 , n29978 , n29979 , n29980 , n29981 , n29982 ,
     n29983 , n29984 , n29985 , n29986 , n29987 , n29988 , n29989 , n29990 , n29991 , n29992 ,
     n29993 , n29994 , n29995 , n29996 , n29997 , n29998 , n29999 , n30000 , n30001 , n30002 ,
     n30003 , n30004 , n30005 , n30006 , n30007 , n30008 , n30009 , n30010 , n30011 , n30012 ,
     n30013 , n30014 , n30015 , n30016 , n30017 , n30018 , n30019 , n30020 , n30021 , n30022 ,
     n30023 , n30024 , n30025 , n30026 , n30027 , n30028 , n30029 , n30030 , n30031 , n30032 ,
     n30033 , n30034 , n30035 , n30036 , n30037 , n30038 , n30039 , n30040 , n30041 , n30042 ,
     n30043 , n30044 , n30045 , n30046 , n30047 , n30048 , n30049 , n30050 , n30051 , n30052 ,
     n30053 , n30054 , n30055 , n30056 , n30057 , n30058 , n30059 , n30060 , n30061 , n30062 ,
     n30063 , n30064 , n30065 , n30066 , n30067 , n30068 , n30069 , n30070 , n30071 , n30072 ,
     n30073 , n30074 , n30075 , n30076 , n30077 , n30078 , n30079 , n30080 , n30081 , n30082 ,
     n30083 , n30084 , n30085 , n30086 , n30087 , n30088 , n30089 , n30090 , n30091 , n30092 ,
     n30093 , n30094 , n30095 , n30096 , n30097 , n30098 , n30099 , n30100 , n30101 , n30102 ,
     n30103 , n30104 , n30105 , n30106 , n30107 , n30108 , n30109 , n30110 , n30111 , n30112 ,
     n30113 , n30114 , n30115 , n30116 , n30117 , n30118 , n30119 , n30120 , n30121 , n30122 ,
     n30123 , n30124 , n30125 , n30126 , n30127 , n30128 , n30129 , n30130 , n30131 , n30132 ,
     n30133 , n30134 , n30135 , n30136 , n30137 , n30138 , n30139 , n30140 , n30141 , n30142 ,
     n30143 , n30144 , n30145 , n30146 , n30147 , n30148 , n30149 , n30150 , n30151 , n30152 ,
     n30153 , n30154 , n30155 , n30156 , n30157 , n30158 , n30159 , n30160 , n30161 , n30162 ,
     n30163 , n30164 , n30165 , n30166 , n30167 , n30168 , n30169 , n30170 , n30171 , n30172 ,
     n30173 , n30174 , n30175 , n30176 , n30177 , n30178 , n30179 , n30180 , n30181 , n30182 ,
     n30183 , n30184 , n30185 , n30186 , n30187 , n30188 , n30189 , n30190 , n30191 , n30192 ,
     n30193 , n30194 , n30195 , n30196 , n30197 , n30198 , n30199 , n30200 , n30201 , n30202 ,
     n30203 , n30204 , n30205 , n30206 , n30207 , n30208 , n30209 , n30210 , n30211 , n30212 ,
     n30213 , n30214 , n30215 , n30216 , n30217 , n30218 , n30219 , n30220 , n30221 , n30222 ,
     n30223 , n30224 , n30225 , n30226 , n30227 , n30228 , n30229 , n30230 , n30231 , n30232 ,
     n30233 , n30234 , n30235 , n30236 , n30237 , n30238 , n30239 , n30240 , n30241 , n30242 ,
     n30243 , n30244 , n30245 , n30246 , n30247 , n30248 , n30249 , n30250 , n30251 , n30252 ,
     n30253 , n30254 , n30255 , n30256 , n30257 , n30258 , n30259 , n30260 , n30261 , n30262 ,
     n30263 , n30264 , n30265 , n30266 , n30267 , n30268 , n30269 , n30270 , n30271 , n30272 ,
     n30273 , n30274 , n30275 , n30276 , n30277 , n30278 , n30279 , n30280 , n30281 , n30282 ,
     n30283 , n30284 , n30285 , n30286 , n30287 , n30288 , n30289 , n30290 , n30291 , n30292 ,
     n30293 , n30294 , n30295 , n30296 , n30297 , n30298 , n30299 , n30300 , n30301 , n30302 ,
     n30303 , n30304 , n30305 , n30306 , n30307 , n30308 , n30309 , n30310 , n30311 , n30312 ,
     n30313 , n30314 , n30315 , n30316 , n30317 , n30318 , n30319 , n30320 , n30321 , n30322 ,
     n30323 , n30324 , n30325 , n30326 , n30327 , n30328 , n30329 , n30330 , n30331 , n30332 ,
     n30333 , n30334 , n30335 , n30336 , n30337 , n30338 , n30339 , n30340 , n30341 , n30342 ,
     n30343 , n30344 , n30345 , n30346 , n30347 , n30348 , n30349 , n30350 , n30351 , n30352 ,
     n30353 , n30354 , n30355 , n30356 , n30357 , n30358 , n30359 , n30360 , n30361 , n30362 ,
     n30363 , n30364 , n30365 , n30366 , n30367 , n30368 , n30369 , n30370 , n30371 , n30372 ,
     n30373 , n30374 , n30375 , n30376 , n30377 , n30378 , n30379 , n30380 , n30381 , n30382 ,
     n30383 , n30384 , n30385 , n30386 , n30387 , n30388 , n30389 , n30390 , n30391 , n30392 ,
     n30393 , n30394 , n30395 , n30396 , n30397 , n30398 , n30399 , n30400 , n30401 , n30402 ,
     n30403 , n30404 , n30405 , n30406 , n30407 , n30408 , n30409 , n30410 , n30411 , n30412 ,
     n30413 , n30414 , n30415 , n30416 , n30417 , n30418 , n30419 , n30420 , n30421 , n30422 ,
     n30423 , n30424 , n30425 , n30426 , n30427 , n30428 , n30429 , n30430 , n30431 , n30432 ,
     n30433 , n30434 , n30435 , n30436 , n30437 , n30438 , n30439 , n30440 , n30441 , n30442 ,
     n30443 , n30444 , n30445 , n30446 , n30447 , n30448 , n30449 , n30450 , n30451 , n30452 ,
     n30453 , n30454 , n30455 , n30456 , n30457 , n30458 , n30459 , n30460 , n30461 , n30462 ,
     n30463 , n30464 , n30465 , n30466 , n30467 , n30468 , n30469 , n30470 , n30471 , n30472 ,
     n30473 , n30474 , n30475 , n30476 , n30477 , n30478 , n30479 , n30480 , n30481 , n30482 ,
     n30483 , n30484 , n30485 , n30486 , n30487 , n30488 , n30489 , n30490 , n30491 , n30492 ,
     n30493 , n30494 , n30495 , n30496 , n30497 , n30498 , n30499 , n30500 , n30501 , n30502 ,
     n30503 , n30504 , n30505 , n30506 , n30507 , n30508 , n30509 , n30510 , n30511 , n30512 ,
     n30513 , n30514 , n30515 , n30516 , n30517 , n30518 , n30519 , n30520 , n30521 , n30522 ,
     n30523 , n30524 , n30525 , n30526 , n30527 , n30528 , n30529 , n30530 , n30531 , n30532 ,
     n30533 , n30534 , n30535 , n30536 , n30537 , n30538 , n30539 , n30540 , n30541 , n30542 ,
     n30543 , n30544 , n30545 , n30546 , n30547 , n30548 , n30549 , n30550 , n30551 , n30552 ,
     n30553 , n30554 , n30555 , n30556 , n30557 , n30558 , n30559 , n30560 , n30561 , n30562 ,
     n30563 , n30564 , n30565 , n30566 , n30567 , n30568 , n30569 , n30570 , n30571 , n30572 ,
     n30573 , n30574 , n30575 , n30576 , n30577 , n30578 , n30579 , n30580 , n30581 , n30582 ,
     n30583 , n30584 , n30585 , n30586 , n30587 , n30588 , n30589 , n30590 , n30591 , n30592 ,
     n30593 , n30594 , n30595 , n30596 , n30597 , n30598 , n30599 , n30600 , n30601 , n30602 ,
     n30603 , n30604 , n30605 , n30606 , n30607 , n30608 , n30609 , n30610 , n30611 , n30612 ,
     n30613 , n30614 , n30615 , n30616 , n30617 , n30618 , n30619 , n30620 , n30621 , n30622 ,
     n30623 , n30624 , n30625 , n30626 , n30627 , n30628 , n30629 , n30630 , n30631 , n30632 ,
     n30633 , n30634 , n30635 , n30636 , n30637 , n30638 , n30639 , n30640 , n30641 , n30642 ,
     n30643 , n30644 , n30645 , n30646 , n30647 , n30648 , n30649 , n30650 , n30651 , n30652 ,
     n30653 , n30654 , n30655 , n30656 , n30657 , n30658 , n30659 , n30660 , n30661 , n30662 ,
     n30663 , n30664 , n30665 , n30666 , n30667 , n30668 , n30669 , n30670 , n30671 , n30672 ,
     n30673 , n30674 , n30675 , n30676 , n30677 , n30678 , n30679 , n30680 , n30681 , n30682 ,
     n30683 , n30684 , n30685 , n30686 , n30687 , n30688 , n30689 , n30690 , n30691 , n30692 ,
     n30693 , n30694 , n30695 , n30696 , n30697 , n30698 , n30699 , n30700 , n30701 , n30702 ,
     n30703 , n30704 , n30705 , n30706 , n30707 , n30708 , n30709 , n30710 , n30711 , n30712 ,
     n30713 , n30714 , n30715 , n30716 , n30717 , n30718 , n30719 , n30720 , n30721 , n30722 ,
     n30723 , n30724 , n30725 , n30726 , n30727 , n30728 , n30729 , n30730 , n30731 , n30732 ,
     n30733 , n30734 , n30735 , n30736 , n30737 , n30738 , n30739 , n30740 , n30741 , n30742 ,
     n30743 , n30744 , n30745 , n30746 , n30747 , n30748 , n30749 , n30750 , n30751 , n30752 ,
     n30753 , n30754 , n30755 , n30756 , n30757 , n30758 , n30759 , n30760 , n30761 , n30762 ,
     n30763 , n30764 , n30765 , n30766 , n30767 , n30768 , n30769 , n30770 , n30771 , n30772 ,
     n30773 , n30774 , n30775 , n30776 , n30777 , n30778 , n30779 , n30780 , n30781 , n30782 ,
     n30783 , n30784 , n30785 , n30786 , n30787 , n30788 , n30789 , n30790 , n30791 , n30792 ,
     n30793 , n30794 , n30795 , n30796 , n30797 , n30798 , n30799 , n30800 , n30801 , n30802 ,
     n30803 , n30804 , n30805 , n30806 , n30807 , n30808 , n30809 , n30810 , n30811 , n30812 ,
     n30813 , n30814 , n30815 , n30816 , n30817 , n30818 , n30819 , n30820 , n30821 , n30822 ,
     n30823 , n30824 , n30825 , n30826 , n30827 , n30828 , n30829 , n30830 , n30831 , n30832 ,
     n30833 , n30834 , n30835 , n30836 , n30837 , n30838 , n30839 , n30840 , n30841 , n30842 ,
     n30843 , n30844 , n30845 , n30846 , n30847 , n30848 , n30849 , n30850 , n30851 , n30852 ,
     n30853 , n30854 , n30855 , n30856 , n30857 , n30858 , n30859 , n30860 , n30861 , n30862 ,
     n30863 , n30864 , n30865 , n30866 , n30867 , n30868 , n30869 , n30870 , n30871 , n30872 ,
     n30873 , n30874 , n30875 , n30876 , n30877 , n30878 , n30879 , n30880 , n30881 , n30882 ,
     n30883 , n30884 , n30885 , n30886 , n30887 , n30888 , n30889 , n30890 , n30891 , n30892 ,
     n30893 , n30894 , n30895 , n30896 , n30897 , n30898 , n30899 , n30900 , n30901 , n30902 ,
     n30903 , n30904 , n30905 , n30906 , n30907 , n30908 , n30909 , n30910 , n30911 , n30912 ,
     n30913 , n30914 , n30915 , n30916 , n30917 , n30918 , n30919 , n30920 , n30921 , n30922 ,
     n30923 , n30924 , n30925 , n30926 , n30927 , n30928 , n30929 , n30930 , n30931 , n30932 ,
     n30933 , n30934 , n30935 , n30936 , n30937 , n30938 , n30939 , n30940 , n30941 , n30942 ,
     n30943 , n30944 , n30945 , n30946 , n30947 , n30948 , n30949 , n30950 , n30951 , n30952 ,
     n30953 , n30954 , n30955 , n30956 , n30957 , n30958 , n30959 , n30960 , n30961 , n30962 ,
     n30963 , n30964 , n30965 , n30966 , n30967 , n30968 , n30969 , n30970 , n30971 , n30972 ,
     n30973 , n30974 , n30975 , n30976 , n30977 , n30978 , n30979 , n30980 , n30981 , n30982 ,
     n30983 , n30984 , n30985 , n30986 , n30987 , n30988 , n30989 , n30990 , n30991 , n30992 ,
     n30993 , n30994 , n30995 , n30996 , n30997 , n30998 , n30999 , n31000 , n31001 , n31002 ,
     n31003 , n31004 , n31005 , n31006 , n31007 , n31008 , n31009 , n31010 , n31011 , n31012 ,
     n31013 , n31014 , n31015 , n31016 , n31017 , n31018 , n31019 , n31020 , n31021 , n31022 ,
     n31023 , n31024 , n31025 , n31026 , n31027 , n31028 , n31029 , n31030 , n31031 , n31032 ,
     n31033 , n31034 , n31035 , n31036 , n31037 , n31038 , n31039 , n31040 , n31041 , n31042 ,
     n31043 , n31044 , n31045 , n31046 , n31047 , n31048 , n31049 , n31050 , n31051 , n31052 ,
     n31053 , n31054 , n31055 , n31056 , n31057 , n31058 , n31059 , n31060 , n31061 , n31062 ,
     n31063 , n31064 , n31065 , n31066 , n31067 , n31068 , n31069 , n31070 , n31071 , n31072 ,
     n31073 , n31074 , n31075 , n31076 , n31077 , n31078 , n31079 , n31080 , n31081 , n31082 ,
     n31083 , n31084 , n31085 , n31086 , n31087 , n31088 , n31089 , n31090 , n31091 , n31092 ,
     n31093 , n31094 , n31095 , n31096 , n31097 , n31098 , n31099 , n31100 , n31101 , n31102 ,
     n31103 , n31104 , n31105 , n31106 , n31107 , n31108 , n31109 , n31110 , n31111 , n31112 ,
     n31113 , n31114 , n31115 , n31116 , n31117 , n31118 , n31119 , n31120 , n31121 , n31122 ,
     n31123 , n31124 , n31125 , n31126 , n31127 , n31128 , n31129 , n31130 , n31131 , n31132 ,
     n31133 , n31134 , n31135 , n31136 , n31137 , n31138 , n31139 , n31140 , n31141 , n31142 ,
     n31143 , n31144 , n31145 , n31146 , n31147 , n31148 , n31149 , n31150 , n31151 , n31152 ,
     n31153 , n31154 , n31155 , n31156 , n31157 , n31158 , n31159 , n31160 , n31161 , n31162 ,
     n31163 , n31164 , n31165 , n31166 , n31167 , n31168 , n31169 , n31170 , n31171 , n31172 ,
     n31173 , n31174 , n31175 , n31176 , n31177 , n31178 , n31179 , n31180 , n31181 , n31182 ,
     n31183 , n31184 , n31185 , n31186 , n31187 , n31188 , n31189 , n31190 , n31191 , n31192 ,
     n31193 , n31194 , n31195 , n31196 , n31197 , n31198 , n31199 , n31200 , n31201 , n31202 ,
     n31203 , n31204 , n31205 , n31206 , n31207 , n31208 , n31209 , n31210 , n31211 , n31212 ,
     n31213 , n31214 , n31215 , n31216 , n31217 , n31218 , n31219 , n31220 , n31221 , n31222 ,
     n31223 , n31224 , n31225 , n31226 , n31227 , n31228 , n31229 , n31230 , n31231 , n31232 ,
     n31233 , n31234 , n31235 , n31236 , n31237 , n31238 , n31239 , n31240 , n31241 , n31242 ,
     n31243 , n31244 , n31245 , n31246 , n31247 , n31248 , n31249 , n31250 , n31251 , n31252 ,
     n31253 , n31254 , n31255 , n31256 , n31257 , n31258 , n31259 , n31260 , n31261 , n31262 ,
     n31263 , n31264 , n31265 , n31266 , n31267 , n31268 , n31269 , n31270 , n31271 , n31272 ,
     n31273 , n31274 , n31275 , n31276 , n31277 , n31278 , n31279 , n31280 , n31281 , n31282 ,
     n31283 , n31284 , n31285 , n31286 , n31287 , n31288 , n31289 , n31290 , n31291 , n31292 ,
     n31293 , n31294 , n31295 , n31296 , n31297 , n31298 , n31299 , n31300 , n31301 , n31302 ,
     n31303 , n31304 , n31305 , n31306 , n31307 , n31308 , n31309 , n31310 , n31311 , n31312 ,
     n31313 , n31314 , n31315 , n31316 , n31317 , n31318 , n31319 , n31320 , n31321 , n31322 ,
     n31323 , n31324 , n31325 , n31326 , n31327 , n31328 , n31329 , n31330 , n31331 , n31332 ,
     n31333 , n31334 , n31335 , n31336 , n31337 , n31338 , n31339 , n31340 , n31341 , n31342 ,
     n31343 , n31344 , n31345 , n31346 , n31347 , n31348 , n31349 , n31350 , n31351 , n31352 ,
     n31353 , n31354 , n31355 , n31356 , n31357 , n31358 , n31359 , n31360 , n31361 , n31362 ,
     n31363 , n31364 , n31365 , n31366 , n31367 , n31368 , n31369 , n31370 , n31371 , n31372 ,
     n31373 , n31374 , n31375 , n31376 , n31377 , n31378 , n31379 , n31380 , n31381 , n31382 ,
     n31383 , n31384 , n31385 , n31386 , n31387 , n31388 , n31389 , n31390 , n31391 , n31392 ,
     n31393 , n31394 , n31395 , n31396 , n31397 , n31398 , n31399 , n31400 , n31401 , n31402 ,
     n31403 , n31404 , n31405 , n31406 , n31407 , n31408 , n31409 , n31410 , n31411 , n31412 ,
     n31413 , n31414 , n31415 , n31416 , n31417 , n31418 , n31419 , n31420 , n31421 , n31422 ,
     n31423 , n31424 , n31425 , n31426 , n31427 , n31428 , n31429 , n31430 , n31431 , n31432 ,
     n31433 , n31434 , n31435 , n31436 , n31437 , n31438 , n31439 , n31440 , n31441 , n31442 ,
     n31443 , n31444 , n31445 , n31446 , n31447 , n31448 , n31449 , n31450 , n31451 , n31452 ,
     n31453 , n31454 , n31455 , n31456 , n31457 , n31458 , n31459 , n31460 , n31461 , n31462 ,
     n31463 , n31464 , n31465 , n31466 , n31467 , n31468 , n31469 , n31470 , n31471 , n31472 ,
     n31473 , n31474 , n31475 , n31476 , n31477 , n31478 , n31479 , n31480 , n31481 , n31482 ,
     n31483 , n31484 , n31485 , n31486 , n31487 , n31488 , n31489 , n31490 , n31491 , n31492 ,
     n31493 , n31494 , n31495 , n31496 , n31497 , n31498 , n31499 , n31500 , n31501 , n31502 ,
     n31503 , n31504 , n31505 , n31506 , n31507 , n31508 , n31509 , n31510 , n31511 , n31512 ,
     n31513 , n31514 , n31515 , n31516 , n31517 , n31518 , n31519 , n31520 , n31521 , n31522 ,
     n31523 , n31524 , n31525 , n31526 , n31527 , n31528 , n31529 , n31530 , n31531 , n31532 ,
     n31533 , n31534 , n31535 , n31536 , n31537 , n31538 , n31539 , n31540 , n31541 , n31542 ,
     n31543 , n31544 , n31545 , n31546 , n31547 , n31548 , n31549 , n31550 , n31551 , n31552 ,
     n31553 , n31554 , n31555 , n31556 , n31557 , n31558 , n31559 , n31560 , n31561 , n31562 ,
     n31563 , n31564 , n31565 , n31566 , n31567 , n31568 , n31569 , n31570 , n31571 , n31572 ,
     n31573 , n31574 , n31575 , n31576 , n31577 , n31578 , n31579 , n31580 , n31581 , n31582 ,
     n31583 , n31584 , n31585 , n31586 , n31587 , n31588 , n31589 , n31590 , n31591 , n31592 ,
     n31593 , n31594 , n31595 , n31596 , n31597 , n31598 , n31599 , n31600 , n31601 , n31602 ,
     n31603 , n31604 , n31605 , n31606 , n31607 , n31608 , n31609 , n31610 , n31611 , n31612 ,
     n31613 , n31614 , n31615 , n31616 , n31617 , n31618 , n31619 , n31620 , n31621 , n31622 ,
     n31623 , n31624 , n31625 , n31626 , n31627 , n31628 , n31629 , n31630 , n31631 , n31632 ,
     n31633 , n31634 , n31635 , n31636 , n31637 , n31638 , n31639 , n31640 , n31641 , n31642 ,
     n31643 , n31644 , n31645 , n31646 , n31647 , n31648 , n31649 , n31650 , n31651 , n31652 ,
     n31653 , n31654 , n31655 , n31656 , n31657 , n31658 , n31659 , n31660 , n31661 , n31662 ,
     n31663 , n31664 , n31665 , n31666 , n31667 , n31668 , n31669 , n31670 , n31671 , n31672 ,
     n31673 , n31674 , n31675 , n31676 , n31677 , n31678 , n31679 , n31680 , n31681 , n31682 ,
     n31683 , n31684 , n31685 , n31686 , n31687 , n31688 , n31689 , n31690 , n31691 , n31692 ,
     n31693 , n31694 , n31695 , n31696 , n31697 , n31698 , n31699 , n31700 , n31701 , n31702 ,
     n31703 , n31704 , n31705 , n31706 , n31707 , n31708 , n31709 , n31710 , n31711 , n31712 ,
     n31713 , n31714 , n31715 , n31716 , n31717 , n31718 , n31719 , n31720 , n31721 , n31722 ,
     n31723 , n31724 , n31725 , n31726 , n31727 , n31728 , n31729 , n31730 , n31731 , n31732 ,
     n31733 , n31734 , n31735 , n31736 , n31737 , n31738 , n31739 , n31740 , n31741 , n31742 ,
     n31743 , n31744 , n31745 , n31746 , n31747 , n31748 , n31749 , n31750 , n31751 , n31752 ,
     n31753 , n31754 , n31755 , n31756 , n31757 , n31758 , n31759 , n31760 , n31761 , n31762 ,
     n31763 , n31764 , n31765 , n31766 , n31767 , n31768 , n31769 , n31770 , n31771 , n31772 ,
     n31773 , n31774 , n31775 , n31776 , n31777 , n31778 , n31779 , n31780 , n31781 , n31782 ,
     n31783 , n31784 , n31785 , n31786 , n31787 , n31788 , n31789 , n31790 , n31791 , n31792 ,
     n31793 , n31794 , n31795 , n31796 , n31797 , n31798 , n31799 , n31800 , n31801 , n31802 ,
     n31803 , n31804 , n31805 , n31806 , n31807 , n31808 , n31809 , n31810 , n31811 , n31812 ,
     n31813 , n31814 , n31815 , n31816 , n31817 , n31818 , n31819 , n31820 , n31821 , n31822 ,
     n31823 , n31824 , n31825 , n31826 , n31827 , n31828 , n31829 , n31830 , n31831 , n31832 ,
     n31833 , n31834 , n31835 , n31836 , n31837 , n31838 , n31839 , n31840 , n31841 , n31842 ,
     n31843 , n31844 , n31845 , n31846 , n31847 , n31848 , n31849 , n31850 , n31851 , n31852 ,
     n31853 , n31854 , n31855 , n31856 , n31857 , n31858 , n31859 , n31860 , n31861 , n31862 ,
     n31863 , n31864 , n31865 , n31866 , n31867 , n31868 , n31869 , n31870 , n31871 , n31872 ,
     n31873 , n31874 , n31875 , n31876 , n31877 , n31878 , n31879 , n31880 , n31881 , n31882 ,
     n31883 , n31884 , n31885 , n31886 , n31887 , n31888 , n31889 , n31890 , n31891 , n31892 ,
     n31893 , n31894 , n31895 , n31896 , n31897 , n31898 , n31899 , n31900 , n31901 , n31902 ,
     n31903 , n31904 , n31905 , n31906 , n31907 , n31908 , n31909 , n31910 , n31911 , n31912 ,
     n31913 , n31914 , n31915 , n31916 , n31917 , n31918 , n31919 , n31920 , n31921 , n31922 ,
     n31923 , n31924 , n31925 , n31926 , n31927 , n31928 , n31929 , n31930 , n31931 , n31932 ,
     n31933 , n31934 , n31935 , n31936 , n31937 , n31938 , n31939 , n31940 , n31941 , n31942 ,
     n31943 , n31944 , n31945 , n31946 , n31947 , n31948 , n31949 , n31950 , n31951 , n31952 ,
     n31953 , n31954 , n31955 , n31956 , n31957 , n31958 , n31959 , n31960 , n31961 , n31962 ,
     n31963 , n31964 , n31965 , n31966 , n31967 , n31968 , n31969 , n31970 , n31971 , n31972 ,
     n31973 , n31974 , n31975 , n31976 , n31977 , n31978 , n31979 , n31980 , n31981 , n31982 ,
     n31983 , n31984 , n31985 , n31986 , n31987 , n31988 , n31989 , n31990 , n31991 , n31992 ,
     n31993 , n31994 , n31995 , n31996 , n31997 , n31998 , n31999 , n32000 , n32001 , n32002 ,
     n32003 , n32004 , n32005 , n32006 , n32007 , n32008 , n32009 , n32010 , n32011 , n32012 ,
     n32013 , n32014 , n32015 , n32016 , n32017 , n32018 , n32019 , n32020 , n32021 , n32022 ,
     n32023 , n32024 , n32025 , n32026 , n32027 , n32028 , n32029 , n32030 , n32031 , n32032 ,
     n32033 , n32034 , n32035 , n32036 , n32037 , n32038 , n32039 , n32040 , n32041 , n32042 ,
     n32043 , n32044 , n32045 , n32046 , n32047 , n32048 , n32049 , n32050 , n32051 , n32052 ,
     n32053 , n32054 , n32055 , n32056 , n32057 , n32058 , n32059 , n32060 , n32061 , n32062 ,
     n32063 , n32064 , n32065 , n32066 , n32067 , n32068 , n32069 , n32070 , n32071 , n32072 ,
     n32073 , n32074 , n32075 , n32076 , n32077 , n32078 , n32079 , n32080 , n32081 , n32082 ,
     n32083 , n32084 , n32085 , n32086 , n32087 , n32088 , n32089 , n32090 , n32091 , n32092 ,
     n32093 , n32094 , n32095 , n32096 , n32097 , n32098 , n32099 , n32100 , n32101 , n32102 ,
     n32103 , n32104 , n32105 , n32106 , n32107 , n32108 , n32109 , n32110 , n32111 , n32112 ,
     n32113 , n32114 , n32115 , n32116 , n32117 , n32118 , n32119 , n32120 , n32121 , n32122 ,
     n32123 , n32124 , n32125 , n32126 , n32127 , n32128 , n32129 , n32130 , n32131 , n32132 ,
     n32133 , n32134 , n32135 , n32136 , n32137 , n32138 , n32139 , n32140 , n32141 , n32142 ,
     n32143 , n32144 , n32145 , n32146 , n32147 , n32148 , n32149 , n32150 , n32151 , n32152 ,
     n32153 , n32154 , n32155 , n32156 , n32157 , n32158 , n32159 , n32160 , n32161 , n32162 ,
     n32163 , n32164 , n32165 , n32166 , n32167 , n32168 , n32169 , n32170 , n32171 , n32172 ,
     n32173 , n32174 , n32175 , n32176 , n32177 , n32178 , n32179 , n32180 , n32181 , n32182 ,
     n32183 , n32184 , n32185 , n32186 , n32187 , n32188 , n32189 , n32190 , n32191 , n32192 ,
     n32193 , n32194 , n32195 , n32196 , n32197 , n32198 , n32199 , n32200 , n32201 , n32202 ,
     n32203 , n32204 , n32205 , n32206 , n32207 , n32208 , n32209 , n32210 , n32211 , n32212 ,
     n32213 , n32214 , n32215 , n32216 , n32217 , n32218 , n32219 , n32220 , n32221 , n32222 ,
     n32223 , n32224 , n32225 , n32226 , n32227 , n32228 , n32229 , n32230 , n32231 , n32232 ,
     n32233 , n32234 , n32235 , n32236 , n32237 , n32238 , n32239 , n32240 , n32241 , n32242 ,
     n32243 , n32244 , n32245 , n32246 , n32247 , n32248 , n32249 , n32250 , n32251 , n32252 ,
     n32253 , n32254 , n32255 , n32256 , n32257 , n32258 , n32259 , n32260 , n32261 , n32262 ,
     n32263 , n32264 , n32265 , n32266 , n32267 , n32268 , n32269 , n32270 , n32271 , n32272 ,
     n32273 , n32274 , n32275 , n32276 , n32277 , n32278 , n32279 , n32280 , n32281 , n32282 ,
     n32283 , n32284 , n32285 , n32286 , n32287 , n32288 , n32289 , n32290 , n32291 , n32292 ,
     n32293 , n32294 , n32295 , n32296 , n32297 , n32298 , n32299 , n32300 , n32301 , n32302 ,
     n32303 , n32304 , n32305 , n32306 , n32307 , n32308 , n32309 , n32310 , n32311 , n32312 ,
     n32313 , n32314 , n32315 , n32316 , n32317 , n32318 , n32319 , n32320 , n32321 , n32322 ,
     n32323 , n32324 , n32325 , n32326 , n32327 , n32328 , n32329 , n32330 , n32331 , n32332 ,
     n32333 , n32334 , n32335 , n32336 , n32337 , n32338 , n32339 , n32340 , n32341 , n32342 ,
     n32343 , n32344 , n32345 , n32346 , n32347 , n32348 , n32349 , n32350 , n32351 , n32352 ,
     n32353 , n32354 , n32355 , n32356 , n32357 , n32358 , n32359 , n32360 , n32361 , n32362 ,
     n32363 , n32364 , n32365 , n32366 , n32367 , n32368 , n32369 , n32370 , n32371 , n32372 ,
     n32373 , n32374 , n32375 , n32376 , n32377 , n32378 , n32379 , n32380 , n32381 , n32382 ,
     n32383 , n32384 , n32385 , n32386 , n32387 , n32388 , n32389 , n32390 , n32391 , n32392 ,
     n32393 , n32394 , n32395 , n32396 , n32397 , n32398 , n32399 , n32400 , n32401 , n32402 ,
     n32403 , n32404 , n32405 , n32406 , n32407 , n32408 , n32409 , n32410 , n32411 , n32412 ,
     n32413 , n32414 , n32415 , n32416 , n32417 , n32418 , n32419 , n32420 , n32421 , n32422 ,
     n32423 , n32424 , n32425 , n32426 , n32427 , n32428 , n32429 , n32430 , n32431 , n32432 ,
     n32433 , n32434 , n32435 , n32436 , n32437 , n32438 , n32439 , n32440 , n32441 , n32442 ,
     n32443 , n32444 , n32445 , n32446 , n32447 , n32448 , n32449 , n32450 , n32451 , n32452 ,
     n32453 , n32454 , n32455 , n32456 , n32457 , n32458 , n32459 , n32460 , n32461 , n32462 ,
     n32463 , n32464 , n32465 , n32466 , n32467 , n32468 , n32469 , n32470 , n32471 , n32472 ,
     n32473 , n32474 , n32475 , n32476 , n32477 , n32478 , n32479 , n32480 , n32481 , n32482 ,
     n32483 , n32484 , n32485 , n32486 , n32487 , n32488 , n32489 , n32490 , n32491 , n32492 ,
     n32493 , n32494 , n32495 , n32496 , n32497 , n32498 , n32499 , n32500 , n32501 , n32502 ,
     n32503 , n32504 , n32505 , n32506 , n32507 , n32508 , n32509 , n32510 , n32511 , n32512 ,
     n32513 , n32514 , n32515 , n32516 , n32517 , n32518 , n32519 , n32520 , n32521 , n32522 ,
     n32523 , n32524 , n32525 , n32526 , n32527 , n32528 , n32529 , n32530 , n32531 , n32532 ,
     n32533 , n32534 , n32535 , n32536 , n32537 , n32538 , n32539 , n32540 , n32541 , n32542 ,
     n32543 , n32544 , n32545 , n32546 , n32547 , n32548 , n32549 , n32550 , n32551 , n32552 ,
     n32553 , n32554 , n32555 , n32556 , n32557 , n32558 , n32559 , n32560 , n32561 , n32562 ,
     n32563 , n32564 , n32565 , n32566 , n32567 , n32568 , n32569 , n32570 , n32571 , n32572 ,
     n32573 , n32574 , n32575 , n32576 , n32577 , n32578 , n32579 , n32580 , n32581 , n32582 ,
     n32583 , n32584 , n32585 , n32586 , n32587 , n32588 , n32589 , n32590 , n32591 , n32592 ,
     n32593 , n32594 , n32595 , n32596 , n32597 , n32598 , n32599 , n32600 , n32601 , n32602 ,
     n32603 , n32604 , n32605 , n32606 , n32607 , n32608 , n32609 , n32610 , n32611 , n32612 ,
     n32613 , n32614 , n32615 , n32616 , n32617 , n32618 , n32619 , n32620 , n32621 , n32622 ,
     n32623 , n32624 , n32625 , n32626 , n32627 , n32628 , n32629 , n32630 , n32631 , n32632 ,
     n32633 , n32634 , n32635 , n32636 , n32637 , n32638 , n32639 , n32640 , n32641 , n32642 ,
     n32643 , n32644 , n32645 , n32646 , n32647 , n32648 , n32649 , n32650 , n32651 , n32652 ,
     n32653 , n32654 , n32655 , n32656 , n32657 , n32658 , n32659 , n32660 , n32661 , n32662 ,
     n32663 , n32664 , n32665 , n32666 , n32667 , n32668 , n32669 , n32670 , n32671 , n32672 ,
     n32673 , n32674 , n32675 , n32676 , n32677 , n32678 , n32679 , n32680 , n32681 , n32682 ,
     n32683 , n32684 , n32685 , n32686 , n32687 , n32688 , n32689 , n32690 , n32691 , n32692 ,
     n32693 , n32694 , n32695 , n32696 , n32697 , n32698 , n32699 , n32700 , n32701 , n32702 ,
     n32703 , n32704 , n32705 , n32706 , n32707 , n32708 , n32709 , n32710 , n32711 , n32712 ,
     n32713 , n32714 , n32715 , n32716 , n32717 , n32718 , n32719 , n32720 , n32721 , n32722 ,
     n32723 , n32724 , n32725 , n32726 , n32727 , n32728 , n32729 , n32730 , n32731 , n32732 ,
     n32733 , n32734 , n32735 , n32736 , n32737 , n32738 , n32739 , n32740 , n32741 , n32742 ,
     n32743 , n32744 , n32745 , n32746 , n32747 , n32748 , n32749 , n32750 , n32751 , n32752 ,
     n32753 , n32754 , n32755 , n32756 , n32757 , n32758 , n32759 , n32760 , n32761 , n32762 ,
     n32763 , n32764 , n32765 , n32766 , n32767 , n32768 , n32769 , n32770 , n32771 , n32772 ,
     n32773 , n32774 , n32775 , n32776 , n32777 , n32778 , n32779 , n32780 , n32781 , n32782 ,
     n32783 , n32784 , n32785 , n32786 , n32787 , n32788 , n32789 , n32790 , n32791 , n32792 ,
     n32793 , n32794 , n32795 , n32796 , n32797 , n32798 , n32799 , n32800 , n32801 , n32802 ,
     n32803 , n32804 , n32805 , n32806 , n32807 , n32808 , n32809 , n32810 , n32811 , n32812 ,
     n32813 , n32814 , n32815 , n32816 , n32817 , n32818 , n32819 , n32820 , n32821 , n32822 ,
     n32823 , n32824 , n32825 , n32826 , n32827 , n32828 , n32829 , n32830 , n32831 , n32832 ,
     n32833 , n32834 , n32835 , n32836 , n32837 , n32838 , n32839 , n32840 , n32841 , n32842 ,
     n32843 , n32844 , n32845 , n32846 , n32847 , n32848 , n32849 , n32850 , n32851 , n32852 ,
     n32853 , n32854 , n32855 , n32856 , n32857 , n32858 , n32859 , n32860 , n32861 , n32862 ,
     n32863 , n32864 , n32865 , n32866 , n32867 , n32868 , n32869 , n32870 , n32871 , n32872 ,
     n32873 , n32874 , n32875 , n32876 , n32877 , n32878 , n32879 , n32880 , n32881 , n32882 ,
     n32883 , n32884 , n32885 , n32886 , n32887 , n32888 , n32889 , n32890 , n32891 , n32892 ,
     n32893 , n32894 , n32895 , n32896 , n32897 , n32898 , n32899 , n32900 , n32901 , n32902 ,
     n32903 , n32904 , n32905 , n32906 , n32907 , n32908 , n32909 , n32910 , n32911 , n32912 ,
     n32913 , n32914 , n32915 , n32916 , n32917 , n32918 , n32919 , n32920 , n32921 , n32922 ,
     n32923 , n32924 , n32925 , n32926 , n32927 , n32928 , n32929 , n32930 , n32931 , n32932 ,
     n32933 , n32934 , n32935 , n32936 , n32937 , n32938 , n32939 , n32940 , n32941 , n32942 ,
     n32943 , n32944 , n32945 , n32946 , n32947 , n32948 , n32949 , n32950 , n32951 , n32952 ,
     n32953 , n32954 , n32955 , n32956 , n32957 , n32958 , n32959 , n32960 , n32961 , n32962 ,
     n32963 , n32964 , n32965 , n32966 , n32967 , n32968 , n32969 , n32970 , n32971 , n32972 ,
     n32973 , n32974 , n32975 , n32976 , n32977 , n32978 , n32979 , n32980 , n32981 , n32982 ,
     n32983 , n32984 , n32985 , n32986 , n32987 , n32988 , n32989 , n32990 , n32991 , n32992 ,
     n32993 , n32994 , n32995 , n32996 , n32997 , n32998 , n32999 , n33000 , n33001 , n33002 ,
     n33003 , n33004 , n33005 , n33006 , n33007 , n33008 , n33009 , n33010 , n33011 , n33012 ,
     n33013 , n33014 , n33015 , n33016 , n33017 , n33018 , n33019 , n33020 , n33021 , n33022 ,
     n33023 , n33024 , n33025 , n33026 , n33027 , n33028 , n33029 , n33030 , n33031 , n33032 ,
     n33033 , n33034 , n33035 , n33036 , n33037 , n33038 , n33039 , n33040 , n33041 , n33042 ,
     n33043 , n33044 , n33045 , n33046 , n33047 , n33048 , n33049 , n33050 , n33051 , n33052 ,
     n33053 , n33054 , n33055 , n33056 , n33057 , n33058 , n33059 , n33060 , n33061 , n33062 ,
     n33063 , n33064 , n33065 , n33066 , n33067 , n33068 , n33069 , n33070 , n33071 , n33072 ,
     n33073 , n33074 , n33075 , n33076 , n33077 , n33078 , n33079 , n33080 , n33081 , n33082 ,
     n33083 , n33084 , n33085 , n33086 , n33087 , n33088 , n33089 , n33090 , n33091 , n33092 ,
     n33093 , n33094 , n33095 , n33096 , n33097 , n33098 , n33099 , n33100 , n33101 , n33102 ,
     n33103 , n33104 , n33105 , n33106 , n33107 , n33108 , n33109 , n33110 , n33111 , n33112 ,
     n33113 , n33114 , n33115 , n33116 , n33117 , n33118 , n33119 , n33120 , n33121 , n33122 ,
     n33123 , n33124 , n33125 , n33126 , n33127 , n33128 , n33129 , n33130 , n33131 , n33132 ,
     n33133 , n33134 , n33135 , n33136 , n33137 , n33138 , n33139 , n33140 , n33141 , n33142 ,
     n33143 , n33144 , n33145 , n33146 , n33147 , n33148 , n33149 , n33150 , n33151 , n33152 ,
     n33153 , n33154 , n33155 , n33156 , n33157 , n33158 , n33159 , n33160 , n33161 , n33162 ,
     n33163 , n33164 , n33165 , n33166 , n33167 , n33168 , n33169 , n33170 , n33171 , n33172 ,
     n33173 , n33174 , n33175 , n33176 , n33177 , n33178 , n33179 , n33180 , n33181 , n33182 ,
     n33183 , n33184 , n33185 , n33186 , n33187 , n33188 , n33189 , n33190 , n33191 , n33192 ,
     n33193 , n33194 , n33195 , n33196 , n33197 , n33198 , n33199 , n33200 , n33201 , n33202 ,
     n33203 , n33204 , n33205 , n33206 , n33207 , n33208 , n33209 , n33210 , n33211 , n33212 ,
     n33213 , n33214 , n33215 , n33216 , n33217 , n33218 , n33219 , n33220 , n33221 , n33222 ,
     n33223 , n33224 , n33225 , n33226 , n33227 , n33228 , n33229 , n33230 , n33231 , n33232 ,
     n33233 , n33234 , n33235 , n33236 , n33237 , n33238 , n33239 , n33240 , n33241 , n33242 ,
     n33243 , n33244 , n33245 , n33246 , n33247 , n33248 , n33249 , n33250 , n33251 , n33252 ,
     n33253 , n33254 , n33255 , n33256 , n33257 , n33258 , n33259 , n33260 , n33261 , n33262 ,
     n33263 , n33264 , n33265 , n33266 , n33267 , n33268 , n33269 , n33270 , n33271 , n33272 ,
     n33273 , n33274 , n33275 , n33276 , n33277 , n33278 , n33279 , n33280 , n33281 , n33282 ,
     n33283 , n33284 , n33285 , n33286 , n33287 , n33288 , n33289 , n33290 , n33291 , n33292 ,
     n33293 , n33294 , n33295 , n33296 , n33297 , n33298 , n33299 , n33300 , n33301 , n33302 ,
     n33303 , n33304 , n33305 , n33306 , n33307 , n33308 , n33309 , n33310 , n33311 , n33312 ,
     n33313 , n33314 , n33315 , n33316 , n33317 , n33318 , n33319 , n33320 , n33321 , n33322 ,
     n33323 , n33324 , n33325 , n33326 , n33327 , n33328 , n33329 , n33330 , n33331 , n33332 ,
     n33333 , n33334 , n33335 , n33336 , n33337 , n33338 , n33339 , n33340 , n33341 , n33342 ,
     n33343 , n33344 , n33345 , n33346 , n33347 , n33348 , n33349 , n33350 , n33351 , n33352 ,
     n33353 , n33354 , n33355 , n33356 , n33357 , n33358 , n33359 , n33360 , n33361 , n33362 ,
     n33363 , n33364 , n33365 , n33366 , n33367 , n33368 , n33369 , n33370 , n33371 , n33372 ,
     n33373 , n33374 , n33375 , n33376 , n33377 , n33378 , n33379 , n33380 , n33381 , n33382 ,
     n33383 , n33384 , n33385 , n33386 , n33387 , n33388 , n33389 , n33390 , n33391 , n33392 ,
     n33393 , n33394 , n33395 , n33396 , n33397 , n33398 , n33399 , n33400 , n33401 , n33402 ,
     n33403 , n33404 , n33405 , n33406 , n33407 , n33408 , n33409 , n33410 , n33411 , n33412 ,
     n33413 , n33414 , n33415 , n33416 , n33417 , n33418 , n33419 , n33420 , n33421 , n33422 ,
     n33423 , n33424 , n33425 , n33426 , n33427 , n33428 , n33429 , n33430 , n33431 , n33432 ,
     n33433 , n33434 , n33435 , n33436 , n33437 , n33438 , n33439 , n33440 , n33441 , n33442 ,
     n33443 , n33444 , n33445 , n33446 , n33447 , n33448 , n33449 , n33450 , n33451 , n33452 ,
     n33453 , n33454 , n33455 , n33456 , n33457 , n33458 , n33459 , n33460 , n33461 , n33462 ,
     n33463 , n33464 , n33465 , n33466 , n33467 , n33468 , n33469 , n33470 , n33471 , n33472 ,
     n33473 , n33474 , n33475 , n33476 , n33477 , n33478 , n33479 , n33480 , n33481 , n33482 ,
     n33483 , n33484 , n33485 , n33486 , n33487 , n33488 , n33489 , n33490 , n33491 , n33492 ,
     n33493 , n33494 , n33495 , n33496 , n33497 , n33498 , n33499 , n33500 , n33501 , n33502 ,
     n33503 , n33504 , n33505 , n33506 , n33507 , n33508 , n33509 , n33510 , n33511 , n33512 ,
     n33513 , n33514 , n33515 , n33516 , n33517 , n33518 , n33519 , n33520 , n33521 , n33522 ,
     n33523 , n33524 , n33525 , n33526 , n33527 , n33528 , n33529 , n33530 , n33531 , n33532 ,
     n33533 , n33534 , n33535 , n33536 , n33537 , n33538 , n33539 , n33540 , n33541 , n33542 ,
     n33543 , n33544 , n33545 , n33546 , n33547 , n33548 , n33549 , n33550 , n33551 , n33552 ,
     n33553 , n33554 , n33555 , n33556 , n33557 , n33558 , n33559 , n33560 , n33561 , n33562 ,
     n33563 , n33564 , n33565 , n33566 , n33567 , n33568 , n33569 , n33570 , n33571 , n33572 ,
     n33573 , n33574 , n33575 , n33576 , n33577 , n33578 , n33579 , n33580 , n33581 , n33582 ,
     n33583 , n33584 , n33585 , n33586 , n33587 , n33588 , n33589 , n33590 , n33591 , n33592 ,
     n33593 , n33594 , n33595 , n33596 , n33597 , n33598 , n33599 , n33600 , n33601 , n33602 ,
     n33603 , n33604 , n33605 , n33606 , n33607 , n33608 , n33609 , n33610 , n33611 , n33612 ,
     n33613 , n33614 , n33615 , n33616 , n33617 , n33618 , n33619 , n33620 , n33621 , n33622 ,
     n33623 , n33624 , n33625 , n33626 , n33627 , n33628 , n33629 , n33630 , n33631 , n33632 ,
     n33633 , n33634 , n33635 , n33636 , n33637 , n33638 , n33639 , n33640 , n33641 , n33642 ,
     n33643 , n33644 , n33645 , n33646 , n33647 , n33648 , n33649 , n33650 , n33651 , n33652 ,
     n33653 , n33654 , n33655 , n33656 , n33657 , n33658 , n33659 , n33660 , n33661 , n33662 ,
     n33663 , n33664 , n33665 , n33666 , n33667 , n33668 , n33669 , n33670 , n33671 , n33672 ,
     n33673 , n33674 , n33675 , n33676 , n33677 , n33678 , n33679 , n33680 , n33681 , n33682 ,
     n33683 , n33684 , n33685 , n33686 , n33687 , n33688 , n33689 , n33690 , n33691 , n33692 ,
     n33693 , n33694 , n33695 , n33696 , n33697 , n33698 , n33699 , n33700 , n33701 , n33702 ,
     n33703 , n33704 , n33705 , n33706 , n33707 , n33708 , n33709 , n33710 , n33711 , n33712 ,
     n33713 , n33714 , n33715 , n33716 , n33717 , n33718 , n33719 , n33720 , n33721 , n33722 ,
     n33723 , n33724 , n33725 , n33726 , n33727 , n33728 , n33729 , n33730 , n33731 , n33732 ,
     n33733 , n33734 , n33735 , n33736 , n33737 , n33738 , n33739 , n33740 , n33741 , n33742 ,
     n33743 , n33744 , n33745 , n33746 , n33747 , n33748 , n33749 , n33750 , n33751 , n33752 ,
     n33753 , n33754 , n33755 , n33756 , n33757 , n33758 , n33759 , n33760 , n33761 , n33762 ,
     n33763 , n33764 , n33765 , n33766 , n33767 , n33768 , n33769 , n33770 , n33771 , n33772 ,
     n33773 , n33774 , n33775 , n33776 , n33777 , n33778 , n33779 , n33780 , n33781 , n33782 ,
     n33783 , n33784 , n33785 , n33786 , n33787 , n33788 , n33789 , n33790 , n33791 , n33792 ,
     n33793 , n33794 , n33795 , n33796 , n33797 , n33798 , n33799 , n33800 , n33801 , n33802 ,
     n33803 , n33804 , n33805 , n33806 , n33807 , n33808 , n33809 , n33810 , n33811 , n33812 ,
     n33813 , n33814 , n33815 , n33816 , n33817 , n33818 , n33819 , n33820 , n33821 , n33822 ,
     n33823 , n33824 , n33825 , n33826 , n33827 , n33828 , n33829 , n33830 , n33831 , n33832 ,
     n33833 , n33834 , n33835 , n33836 , n33837 , n33838 , n33839 , n33840 , n33841 , n33842 ,
     n33843 , n33844 , n33845 , n33846 , n33847 , n33848 , n33849 , n33850 , n33851 , n33852 ,
     n33853 , n33854 , n33855 , n33856 , n33857 , n33858 , n33859 , n33860 , n33861 , n33862 ,
     n33863 , n33864 , n33865 , n33866 , n33867 , n33868 , n33869 , n33870 , n33871 , n33872 ,
     n33873 , n33874 , n33875 , n33876 , n33877 , n33878 , n33879 , n33880 , n33881 , n33882 ,
     n33883 , n33884 , n33885 , n33886 , n33887 , n33888 , n33889 , n33890 , n33891 , n33892 ,
     n33893 , n33894 , n33895 , n33896 , n33897 , n33898 , n33899 , n33900 , n33901 , n33902 ,
     n33903 , n33904 , n33905 , n33906 , n33907 , n33908 , n33909 , n33910 , n33911 , n33912 ,
     n33913 , n33914 , n33915 , n33916 , n33917 , n33918 , n33919 , n33920 , n33921 , n33922 ,
     n33923 , n33924 , n33925 , n33926 , n33927 , n33928 , n33929 , n33930 , n33931 , n33932 ,
     n33933 , n33934 , n33935 , n33936 , n33937 , n33938 , n33939 , n33940 , n33941 , n33942 ,
     n33943 , n33944 , n33945 , n33946 , n33947 , n33948 , n33949 , n33950 , n33951 , n33952 ,
     n33953 , n33954 , n33955 , n33956 , n33957 , n33958 , n33959 , n33960 , n33961 , n33962 ,
     n33963 , n33964 , n33965 , n33966 , n33967 , n33968 , n33969 , n33970 , n33971 , n33972 ,
     n33973 , n33974 , n33975 , n33976 , n33977 , n33978 , n33979 , n33980 , n33981 , n33982 ,
     n33983 , n33984 , n33985 , n33986 , n33987 , n33988 , n33989 , n33990 , n33991 , n33992 ,
     n33993 , n33994 , n33995 , n33996 , n33997 , n33998 , n33999 , n34000 , n34001 , n34002 ,
     n34003 , n34004 , n34005 , n34006 , n34007 , n34008 , n34009 , n34010 , n34011 , n34012 ,
     n34013 , n34014 , n34015 , n34016 , n34017 , n34018 , n34019 , n34020 , n34021 , n34022 ,
     n34023 , n34024 , n34025 , n34026 , n34027 , n34028 , n34029 , n34030 , n34031 , n34032 ,
     n34033 , n34034 , n34035 , n34036 , n34037 , n34038 , n34039 , n34040 , n34041 , n34042 ,
     n34043 , n34044 , n34045 , n34046 , n34047 , n34048 , n34049 , n34050 , n34051 , n34052 ,
     n34053 , n34054 , n34055 , n34056 , n34057 , n34058 , n34059 , n34060 , n34061 , n34062 ,
     n34063 , n34064 , n34065 , n34066 , n34067 , n34068 , n34069 , n34070 , n34071 , n34072 ,
     n34073 , n34074 , n34075 , n34076 , n34077 , n34078 , n34079 , n34080 , n34081 , n34082 ,
     n34083 , n34084 , n34085 , n34086 , n34087 , n34088 , n34089 , n34090 , n34091 , n34092 ,
     n34093 , n34094 , n34095 , n34096 , n34097 , n34098 , n34099 , n34100 , n34101 , n34102 ,
     n34103 , n34104 , n34105 , n34106 , n34107 , n34108 , n34109 , n34110 , n34111 , n34112 ,
     n34113 , n34114 , n34115 , n34116 , n34117 , n34118 , n34119 , n34120 , n34121 , n34122 ,
     n34123 , n34124 , n34125 , n34126 , n34127 , n34128 , n34129 , n34130 , n34131 , n34132 ,
     n34133 , n34134 , n34135 , n34136 , n34137 , n34138 , n34139 , n34140 , n34141 , n34142 ,
     n34143 , n34144 , n34145 , n34146 , n34147 , n34148 , n34149 , n34150 , n34151 , n34152 ,
     n34153 , n34154 , n34155 , n34156 , n34157 , n34158 , n34159 , n34160 , n34161 , n34162 ,
     n34163 , n34164 , n34165 , n34166 , n34167 , n34168 , n34169 , n34170 , n34171 , n34172 ,
     n34173 , n34174 , n34175 , n34176 , n34177 , n34178 , n34179 , n34180 , n34181 , n34182 ,
     n34183 , n34184 , n34185 , n34186 , n34187 , n34188 , n34189 , n34190 , n34191 , n34192 ,
     n34193 , n34194 , n34195 , n34196 , n34197 , n34198 , n34199 , n34200 , n34201 , n34202 ,
     n34203 , n34204 , n34205 , n34206 , n34207 , n34208 , n34209 , n34210 , n34211 , n34212 ,
     n34213 , n34214 , n34215 , n34216 , n34217 , n34218 , n34219 , n34220 , n34221 , n34222 ,
     n34223 , n34224 , n34225 , n34226 , n34227 , n34228 , n34229 , n34230 , n34231 , n34232 ,
     n34233 , n34234 , n34235 , n34236 , n34237 , n34238 , n34239 , n34240 , n34241 , n34242 ,
     n34243 , n34244 , n34245 , n34246 , n34247 , n34248 , n34249 , n34250 , n34251 , n34252 ,
     n34253 , n34254 , n34255 , n34256 , n34257 , n34258 , n34259 , n34260 , n34261 , n34262 ,
     n34263 , n34264 , n34265 , n34266 , n34267 , n34268 , n34269 , n34270 , n34271 , n34272 ,
     n34273 , n34274 , n34275 , n34276 , n34277 , n34278 , n34279 , n34280 , n34281 , n34282 ,
     n34283 , n34284 , n34285 , n34286 , n34287 , n34288 , n34289 , n34290 , n34291 , n34292 ,
     n34293 , n34294 , n34295 , n34296 , n34297 , n34298 , n34299 , n34300 , n34301 , n34302 ,
     n34303 , n34304 , n34305 , n34306 , n34307 , n34308 , n34309 , n34310 , n34311 , n34312 ,
     n34313 , n34314 , n34315 , n34316 , n34317 , n34318 , n34319 , n34320 , n34321 , n34322 ,
     n34323 , n34324 , n34325 , n34326 , n34327 , n34328 , n34329 , n34330 , n34331 , n34332 ,
     n34333 , n34334 , n34335 , n34336 , n34337 , n34338 , n34339 , n34340 , n34341 , n34342 ,
     n34343 , n34344 , n34345 , n34346 , n34347 , n34348 , n34349 , n34350 , n34351 , n34352 ,
     n34353 , n34354 , n34355 , n34356 , n34357 , n34358 , n34359 , n34360 , n34361 , n34362 ,
     n34363 , n34364 , n34365 , n34366 , n34367 , n34368 , n34369 , n34370 , n34371 , n34372 ,
     n34373 , n34374 , n34375 , n34376 , n34377 , n34378 , n34379 , n34380 , n34381 , n34382 ,
     n34383 , n34384 , n34385 , n34386 , n34387 , n34388 , n34389 , n34390 , n34391 , n34392 ,
     n34393 , n34394 , n34395 , n34396 , n34397 , n34398 , n34399 , n34400 , n34401 , n34402 ,
     n34403 , n34404 , n34405 , n34406 , n34407 , n34408 , n34409 , n34410 , n34411 , n34412 ,
     n34413 , n34414 , n34415 , n34416 , n34417 , n34418 , n34419 , n34420 , n34421 , n34422 ,
     n34423 , n34424 , n34425 , n34426 , n34427 , n34428 , n34429 , n34430 , n34431 , n34432 ,
     n34433 , n34434 , n34435 , n34436 , n34437 , n34438 , n34439 , n34440 , n34441 , n34442 ,
     n34443 , n34444 , n34445 , n34446 , n34447 , n34448 , n34449 , n34450 , n34451 , n34452 ,
     n34453 , n34454 , n34455 , n34456 , n34457 , n34458 , n34459 , n34460 , n34461 , n34462 ,
     n34463 , n34464 , n34465 , n34466 , n34467 , n34468 , n34469 , n34470 , n34471 , n34472 ,
     n34473 , n34474 , n34475 , n34476 , n34477 , n34478 , n34479 , n34480 , n34481 , n34482 ,
     n34483 , n34484 , n34485 , n34486 , n34487 , n34488 , n34489 , n34490 , n34491 , n34492 ,
     n34493 , n34494 , n34495 , n34496 , n34497 , n34498 , n34499 , n34500 , n34501 , n34502 ,
     n34503 , n34504 , n34505 , n34506 , n34507 , n34508 , n34509 , n34510 , n34511 , n34512 ,
     n34513 , n34514 , n34515 , n34516 , n34517 , n34518 , n34519 , n34520 , n34521 , n34522 ,
     n34523 , n34524 , n34525 , n34526 , n34527 , n34528 , n34529 , n34530 , n34531 , n34532 ,
     n34533 , n34534 , n34535 , n34536 , n34537 , n34538 , n34539 , n34540 , n34541 , n34542 ,
     n34543 , n34544 , n34545 , n34546 , n34547 , n34548 , n34549 , n34550 , n34551 , n34552 ,
     n34553 , n34554 , n34555 , n34556 , n34557 , n34558 , n34559 , n34560 , n34561 , n34562 ,
     n34563 , n34564 , n34565 , n34566 , n34567 , n34568 , n34569 , n34570 , n34571 , n34572 ,
     n34573 , n34574 , n34575 , n34576 , n34577 , n34578 , n34579 , n34580 , n34581 , n34582 ,
     n34583 , n34584 , n34585 , n34586 , n34587 , n34588 , n34589 , n34590 , n34591 , n34592 ,
     n34593 , n34594 , n34595 , n34596 , n34597 , n34598 , n34599 , n34600 , n34601 , n34602 ,
     n34603 , n34604 , n34605 , n34606 , n34607 , n34608 , n34609 , n34610 , n34611 , n34612 ,
     n34613 , n34614 , n34615 , n34616 , n34617 , n34618 , n34619 , n34620 , n34621 , n34622 ,
     n34623 , n34624 , n34625 , n34626 , n34627 , n34628 , n34629 , n34630 , n34631 , n34632 ,
     n34633 , n34634 , n34635 , n34636 , n34637 , n34638 , n34639 , n34640 , n34641 , n34642 ,
     n34643 , n34644 , n34645 , n34646 , n34647 , n34648 , n34649 , n34650 , n34651 , n34652 ,
     n34653 , n34654 , n34655 , n34656 , n34657 , n34658 , n34659 , n34660 , n34661 , n34662 ,
     n34663 , n34664 , n34665 , n34666 , n34667 , n34668 , n34669 , n34670 , n34671 , n34672 ,
     n34673 , n34674 , n34675 , n34676 , n34677 , n34678 , n34679 , n34680 , n34681 , n34682 ,
     n34683 , n34684 , n34685 , n34686 , n34687 , n34688 , n34689 , n34690 , n34691 , n34692 ,
     n34693 , n34694 , n34695 , n34696 , n34697 , n34698 , n34699 , n34700 , n34701 , n34702 ,
     n34703 , n34704 , n34705 , n34706 , n34707 , n34708 , n34709 , n34710 , n34711 , n34712 ,
     n34713 , n34714 , n34715 , n34716 , n34717 , n34718 , n34719 , n34720 , n34721 , n34722 ,
     n34723 , n34724 , n34725 , n34726 , n34727 , n34728 , n34729 , n34730 , n34731 , n34732 ,
     n34733 , n34734 , n34735 , n34736 , n34737 , n34738 , n34739 , n34740 , n34741 , n34742 ,
     n34743 , n34744 , n34745 , n34746 , n34747 , n34748 , n34749 , n34750 , n34751 , n34752 ,
     n34753 , n34754 , n34755 , n34756 , n34757 , n34758 , n34759 , n34760 , n34761 , n34762 ,
     n34763 , n34764 , n34765 , n34766 , n34767 , n34768 , n34769 , n34770 , n34771 , n34772 ,
     n34773 , n34774 , n34775 , n34776 , n34777 , n34778 , n34779 , n34780 , n34781 , n34782 ,
     n34783 , n34784 , n34785 , n34786 , n34787 , n34788 , n34789 , n34790 , n34791 , n34792 ,
     n34793 , n34794 , n34795 , n34796 , n34797 , n34798 , n34799 , n34800 , n34801 , n34802 ,
     n34803 , n34804 , n34805 , n34806 , n34807 , n34808 , n34809 , n34810 , n34811 , n34812 ,
     n34813 , n34814 , n34815 , n34816 , n34817 , n34818 , n34819 , n34820 , n34821 , n34822 ,
     n34823 , n34824 , n34825 , n34826 , n34827 , n34828 , n34829 , n34830 , n34831 , n34832 ,
     n34833 , n34834 , n34835 , n34836 , n34837 , n34838 , n34839 , n34840 , n34841 , n34842 ,
     n34843 , n34844 , n34845 , n34846 , n34847 , n34848 , n34849 , n34850 , n34851 , n34852 ,
     n34853 , n34854 , n34855 , n34856 , n34857 , n34858 , n34859 , n34860 , n34861 , n34862 ,
     n34863 , n34864 , n34865 , n34866 , n34867 , n34868 , n34869 , n34870 , n34871 , n34872 ,
     n34873 , n34874 , n34875 , n34876 , n34877 , n34878 , n34879 , n34880 , n34881 , n34882 ,
     n34883 , n34884 , n34885 , n34886 , n34887 , n34888 , n34889 , n34890 , n34891 , n34892 ,
     n34893 , n34894 , n34895 , n34896 , n34897 , n34898 , n34899 , n34900 , n34901 , n34902 ,
     n34903 , n34904 , n34905 , n34906 , n34907 , n34908 , n34909 , n34910 , n34911 , n34912 ,
     n34913 , n34914 , n34915 , n34916 , n34917 , n34918 , n34919 , n34920 , n34921 , n34922 ,
     n34923 , n34924 , n34925 , n34926 , n34927 , n34928 , n34929 , n34930 , n34931 , n34932 ,
     n34933 , n34934 , n34935 , n34936 , n34937 , n34938 , n34939 , n34940 , n34941 , n34942 ,
     n34943 , n34944 , n34945 , n34946 , n34947 , n34948 , n34949 , n34950 , n34951 , n34952 ,
     n34953 , n34954 , n34955 , n34956 , n34957 , n34958 , n34959 , n34960 , n34961 , n34962 ,
     n34963 , n34964 , n34965 , n34966 , n34967 , n34968 , n34969 , n34970 , n34971 , n34972 ,
     n34973 , n34974 , n34975 , n34976 , n34977 , n34978 , n34979 , n34980 , n34981 , n34982 ,
     n34983 , n34984 , n34985 , n34986 , n34987 , n34988 , n34989 , n34990 , n34991 , n34992 ,
     n34993 , n34994 , n34995 , n34996 , n34997 , n34998 , n34999 , n35000 , n35001 , n35002 ,
     n35003 , n35004 , n35005 , n35006 , n35007 , n35008 , n35009 , n35010 , n35011 , n35012 ,
     n35013 , n35014 , n35015 , n35016 , n35017 , n35018 , n35019 , n35020 , n35021 , n35022 ,
     n35023 , n35024 , n35025 , n35026 , n35027 , n35028 , n35029 , n35030 , n35031 , n35032 ,
     n35033 , n35034 , n35035 , n35036 , n35037 , n35038 , n35039 , n35040 , n35041 , n35042 ,
     n35043 , n35044 , n35045 , n35046 , n35047 , n35048 , n35049 , n35050 , n35051 , n35052 ,
     n35053 , n35054 , n35055 , n35056 , n35057 , n35058 , n35059 , n35060 , n35061 , n35062 ,
     n35063 , n35064 , n35065 , n35066 , n35067 , n35068 , n35069 , n35070 , n35071 , n35072 ,
     n35073 , n35074 , n35075 , n35076 , n35077 , n35078 , n35079 , n35080 , n35081 , n35082 ,
     n35083 , n35084 , n35085 , n35086 , n35087 , n35088 , n35089 , n35090 , n35091 , n35092 ,
     n35093 , n35094 , n35095 , n35096 , n35097 , n35098 , n35099 , n35100 , n35101 , n35102 ,
     n35103 , n35104 , n35105 , n35106 , n35107 , n35108 , n35109 , n35110 , n35111 , n35112 ,
     n35113 , n35114 , n35115 , n35116 , n35117 , n35118 , n35119 , n35120 , n35121 , n35122 ,
     n35123 , n35124 , n35125 , n35126 , n35127 , n35128 , n35129 , n35130 , n35131 , n35132 ,
     n35133 , n35134 , n35135 , n35136 , n35137 , n35138 , n35139 , n35140 , n35141 , n35142 ,
     n35143 , n35144 , n35145 , n35146 , n35147 , n35148 , n35149 , n35150 , n35151 , n35152 ,
     n35153 , n35154 , n35155 , n35156 , n35157 , n35158 , n35159 , n35160 , n35161 , n35162 ,
     n35163 , n35164 , n35165 , n35166 , n35167 , n35168 , n35169 , n35170 , n35171 , n35172 ,
     n35173 , n35174 , n35175 , n35176 , n35177 , n35178 , n35179 , n35180 , n35181 , n35182 ,
     n35183 , n35184 , n35185 , n35186 , n35187 , n35188 , n35189 , n35190 , n35191 , n35192 ,
     n35193 , n35194 , n35195 , n35196 , n35197 , n35198 , n35199 , n35200 , n35201 , n35202 ,
     n35203 , n35204 , n35205 , n35206 , n35207 , n35208 , n35209 , n35210 , n35211 , n35212 ,
     n35213 , n35214 , n35215 , n35216 , n35217 , n35218 , n35219 , n35220 , n35221 , n35222 ,
     n35223 , n35224 , n35225 , n35226 , n35227 , n35228 , n35229 , n35230 , n35231 , n35232 ,
     n35233 , n35234 , n35235 , n35236 , n35237 , n35238 , n35239 , n35240 , n35241 , n35242 ,
     n35243 , n35244 , n35245 , n35246 , n35247 , n35248 , n35249 , n35250 , n35251 , n35252 ,
     n35253 , n35254 , n35255 , n35256 , n35257 , n35258 , n35259 , n35260 , n35261 , n35262 ,
     n35263 , n35264 , n35265 , n35266 , n35267 , n35268 , n35269 , n35270 , n35271 , n35272 ,
     n35273 , n35274 , n35275 , n35276 , n35277 , n35278 , n35279 , n35280 , n35281 , n35282 ,
     n35283 , n35284 , n35285 , n35286 , n35287 , n35288 , n35289 , n35290 , n35291 , n35292 ,
     n35293 , n35294 , n35295 , n35296 , n35297 , n35298 , n35299 , n35300 , n35301 , n35302 ,
     n35303 , n35304 , n35305 , n35306 , n35307 , n35308 , n35309 , n35310 , n35311 , n35312 ,
     n35313 , n35314 , n35315 , n35316 , n35317 , n35318 , n35319 , n35320 , n35321 , n35322 ,
     n35323 , n35324 , n35325 , n35326 , n35327 , n35328 , n35329 , n35330 , n35331 , n35332 ,
     n35333 , n35334 , n35335 , n35336 , n35337 , n35338 , n35339 , n35340 , n35341 , n35342 ,
     n35343 , n35344 , n35345 , n35346 , n35347 , n35348 , n35349 , n35350 , n35351 , n35352 ,
     n35353 , n35354 , n35355 , n35356 , n35357 , n35358 , n35359 , n35360 , n35361 , n35362 ,
     n35363 , n35364 , n35365 , n35366 , n35367 , n35368 , n35369 , n35370 , n35371 , n35372 ,
     n35373 , n35374 , n35375 , n35376 , n35377 , n35378 , n35379 , n35380 , n35381 , n35382 ,
     n35383 , n35384 , n35385 , n35386 , n35387 , n35388 , n35389 , n35390 , n35391 , n35392 ,
     n35393 , n35394 , n35395 , n35396 , n35397 , n35398 , n35399 , n35400 , n35401 , n35402 ,
     n35403 , n35404 , n35405 , n35406 , n35407 , n35408 , n35409 , n35410 , n35411 , n35412 ,
     n35413 , n35414 , n35415 , n35416 , n35417 , n35418 , n35419 , n35420 , n35421 , n35422 ,
     n35423 , n35424 , n35425 , n35426 , n35427 , n35428 , n35429 , n35430 , n35431 , n35432 ,
     n35433 , n35434 , n35435 , n35436 , n35437 , n35438 , n35439 , n35440 , n35441 , n35442 ,
     n35443 , n35444 , n35445 , n35446 , n35447 , n35448 , n35449 , n35450 , n35451 , n35452 ,
     n35453 , n35454 , n35455 , n35456 , n35457 , n35458 , n35459 , n35460 , n35461 , n35462 ,
     n35463 , n35464 , n35465 , n35466 , n35467 , n35468 , n35469 , n35470 , n35471 , n35472 ,
     n35473 , n35474 , n35475 , n35476 , n35477 , n35478 , n35479 , n35480 , n35481 , n35482 ,
     n35483 , n35484 , n35485 , n35486 , n35487 , n35488 , n35489 , n35490 , n35491 , n35492 ,
     n35493 , n35494 , n35495 , n35496 , n35497 , n35498 , n35499 , n35500 , n35501 , n35502 ,
     n35503 , n35504 , n35505 , n35506 , n35507 , n35508 , n35509 , n35510 , n35511 , n35512 ,
     n35513 , n35514 , n35515 , n35516 , n35517 , n35518 , n35519 , n35520 , n35521 , n35522 ,
     n35523 , n35524 , n35525 , n35526 , n35527 , n35528 , n35529 , n35530 , n35531 , n35532 ,
     n35533 , n35534 , n35535 , n35536 , n35537 , n35538 , n35539 , n35540 , n35541 , n35542 ,
     n35543 , n35544 , n35545 , n35546 , n35547 , n35548 , n35549 , n35550 , n35551 , n35552 ,
     n35553 , n35554 , n35555 , n35556 , n35557 , n35558 , n35559 , n35560 , n35561 , n35562 ,
     n35563 , n35564 , n35565 , n35566 , n35567 , n35568 , n35569 , n35570 , n35571 , n35572 ,
     n35573 , n35574 , n35575 , n35576 , n35577 , n35578 , n35579 , n35580 , n35581 , n35582 ,
     n35583 , n35584 , n35585 , n35586 , n35587 , n35588 , n35589 , n35590 , n35591 , n35592 ,
     n35593 , n35594 , n35595 , n35596 , n35597 , n35598 , n35599 , n35600 , n35601 , n35602 ,
     n35603 , n35604 , n35605 , n35606 , n35607 , n35608 , n35609 , n35610 , n35611 , n35612 ,
     n35613 , n35614 , n35615 , n35616 , n35617 , n35618 , n35619 , n35620 , n35621 , n35622 ,
     n35623 , n35624 , n35625 , n35626 , n35627 , n35628 , n35629 , n35630 , n35631 , n35632 ,
     n35633 , n35634 , n35635 , n35636 , n35637 , n35638 , n35639 , n35640 , n35641 , n35642 ,
     n35643 , n35644 , n35645 , n35646 , n35647 , n35648 , n35649 , n35650 , n35651 , n35652 ,
     n35653 , n35654 , n35655 , n35656 , n35657 , n35658 , n35659 , n35660 , n35661 , n35662 ,
     n35663 , n35664 , n35665 , n35666 , n35667 , n35668 , n35669 , n35670 , n35671 , n35672 ,
     n35673 , n35674 , n35675 , n35676 , n35677 , n35678 , n35679 , n35680 , n35681 , n35682 ,
     n35683 , n35684 , n35685 , n35686 , n35687 , n35688 , n35689 , n35690 , n35691 , n35692 ,
     n35693 , n35694 , n35695 , n35696 , n35697 , n35698 , n35699 , n35700 , n35701 , n35702 ,
     n35703 , n35704 , n35705 , n35706 , n35707 , n35708 , n35709 , n35710 , n35711 , n35712 ,
     n35713 , n35714 , n35715 , n35716 , n35717 , n35718 , n35719 , n35720 , n35721 , n35722 ,
     n35723 , n35724 , n35725 , n35726 , n35727 , n35728 , n35729 , n35730 , n35731 , n35732 ,
     n35733 , n35734 , n35735 , n35736 , n35737 , n35738 , n35739 , n35740 , n35741 , n35742 ,
     n35743 , n35744 , n35745 , n35746 , n35747 , n35748 , n35749 , n35750 , n35751 , n35752 ,
     n35753 , n35754 , n35755 , n35756 , n35757 , n35758 , n35759 , n35760 , n35761 , n35762 ,
     n35763 , n35764 , n35765 , n35766 , n35767 , n35768 , n35769 , n35770 , n35771 , n35772 ,
     n35773 , n35774 , n35775 , n35776 , n35777 , n35778 , n35779 , n35780 , n35781 , n35782 ,
     n35783 , n35784 , n35785 , n35786 , n35787 , n35788 , n35789 , n35790 , n35791 , n35792 ,
     n35793 , n35794 , n35795 , n35796 , n35797 , n35798 , n35799 , n35800 , n35801 , n35802 ,
     n35803 , n35804 , n35805 , n35806 , n35807 , n35808 , n35809 , n35810 , n35811 , n35812 ,
     n35813 , n35814 , n35815 , n35816 , n35817 , n35818 , n35819 , n35820 , n35821 , n35822 ,
     n35823 , n35824 , n35825 , n35826 , n35827 , n35828 , n35829 , n35830 , n35831 , n35832 ,
     n35833 , n35834 , n35835 , n35836 , n35837 , n35838 , n35839 , n35840 , n35841 , n35842 ,
     n35843 , n35844 , n35845 , n35846 , n35847 , n35848 , n35849 , n35850 , n35851 , n35852 ,
     n35853 , n35854 , n35855 , n35856 , n35857 , n35858 , n35859 , n35860 , n35861 , n35862 ,
     n35863 , n35864 , n35865 , n35866 , n35867 , n35868 , n35869 , n35870 , n35871 , n35872 ,
     n35873 , n35874 , n35875 , n35876 , n35877 , n35878 , n35879 , n35880 , n35881 , n35882 ,
     n35883 , n35884 , n35885 , n35886 , n35887 , n35888 , n35889 , n35890 , n35891 , n35892 ,
     n35893 , n35894 , n35895 , n35896 , n35897 , n35898 , n35899 , n35900 , n35901 , n35902 ,
     n35903 , n35904 , n35905 , n35906 , n35907 , n35908 , n35909 , n35910 , n35911 , n35912 ,
     n35913 , n35914 , n35915 , n35916 , n35917 , n35918 , n35919 , n35920 , n35921 , n35922 ,
     n35923 , n35924 , n35925 , n35926 , n35927 , n35928 , n35929 , n35930 , n35931 , n35932 ,
     n35933 , n35934 , n35935 , n35936 , n35937 , n35938 , n35939 , n35940 , n35941 , n35942 ,
     n35943 , n35944 , n35945 , n35946 , n35947 , n35948 , n35949 , n35950 , n35951 , n35952 ,
     n35953 , n35954 , n35955 , n35956 , n35957 , n35958 , n35959 , n35960 , n35961 , n35962 ,
     n35963 , n35964 , n35965 , n35966 , n35967 , n35968 , n35969 , n35970 , n35971 , n35972 ,
     n35973 , n35974 , n35975 , n35976 , n35977 , n35978 , n35979 , n35980 , n35981 , n35982 ,
     n35983 , n35984 , n35985 , n35986 , n35987 , n35988 , n35989 , n35990 , n35991 , n35992 ,
     n35993 , n35994 , n35995 , n35996 , n35997 , n35998 , n35999 , n36000 , n36001 , n36002 ,
     n36003 , n36004 , n36005 , n36006 , n36007 , n36008 , n36009 , n36010 , n36011 , n36012 ,
     n36013 , n36014 , n36015 , n36016 , n36017 , n36018 , n36019 , n36020 , n36021 , n36022 ,
     n36023 , n36024 , n36025 , n36026 , n36027 , n36028 , n36029 , n36030 , n36031 , n36032 ,
     n36033 , n36034 , n36035 , n36036 , n36037 , n36038 , n36039 , n36040 , n36041 , n36042 ,
     n36043 , n36044 , n36045 , n36046 , n36047 , n36048 , n36049 , n36050 , n36051 , n36052 ,
     n36053 , n36054 , n36055 , n36056 , n36057 , n36058 , n36059 , n36060 , n36061 , n36062 ,
     n36063 , n36064 , n36065 , n36066 , n36067 , n36068 , n36069 , n36070 , n36071 , n36072 ,
     n36073 , n36074 , n36075 , n36076 , n36077 , n36078 , n36079 , n36080 , n36081 , n36082 ,
     n36083 , n36084 , n36085 , n36086 , n36087 , n36088 , n36089 , n36090 , n36091 , n36092 ,
     n36093 , n36094 , n36095 , n36096 , n36097 , n36098 , n36099 , n36100 , n36101 , n36102 ,
     n36103 , n36104 , n36105 , n36106 , n36107 , n36108 , n36109 , n36110 , n36111 , n36112 ,
     n36113 , n36114 , n36115 , n36116 , n36117 , n36118 , n36119 , n36120 , n36121 , n36122 ,
     n36123 , n36124 , n36125 , n36126 , n36127 , n36128 , n36129 , n36130 , n36131 , n36132 ,
     n36133 , n36134 , n36135 , n36136 , n36137 , n36138 , n36139 , n36140 , n36141 , n36142 ,
     n36143 , n36144 , n36145 , n36146 , n36147 , n36148 , n36149 , n36150 , n36151 , n36152 ,
     n36153 , n36154 , n36155 , n36156 , n36157 , n36158 , n36159 , n36160 , n36161 , n36162 ,
     n36163 , n36164 , n36165 , n36166 , n36167 , n36168 , n36169 , n36170 , n36171 , n36172 ,
     n36173 , n36174 , n36175 , n36176 , n36177 , n36178 , n36179 , n36180 , n36181 , n36182 ,
     n36183 , n36184 , n36185 , n36186 , n36187 , n36188 , n36189 , n36190 , n36191 , n36192 ,
     n36193 , n36194 , n36195 , n36196 , n36197 , n36198 , n36199 , n36200 , n36201 , n36202 ,
     n36203 , n36204 , n36205 , n36206 , n36207 , n36208 , n36209 , n36210 , n36211 , n36212 ,
     n36213 , n36214 , n36215 , n36216 , n36217 , n36218 , n36219 , n36220 , n36221 , n36222 ,
     n36223 , n36224 , n36225 , n36226 , n36227 , n36228 , n36229 , n36230 , n36231 , n36232 ,
     n36233 , n36234 , n36235 , n36236 , n36237 , n36238 , n36239 , n36240 , n36241 , n36242 ,
     n36243 , n36244 , n36245 , n36246 , n36247 , n36248 , n36249 , n36250 , n36251 , n36252 ,
     n36253 , n36254 , n36255 , n36256 , n36257 , n36258 , n36259 , n36260 , n36261 , n36262 ,
     n36263 , n36264 , n36265 , n36266 , n36267 , n36268 , n36269 , n36270 , n36271 , n36272 ,
     n36273 , n36274 , n36275 , n36276 , n36277 , n36278 , n36279 , n36280 , n36281 , n36282 ,
     n36283 , n36284 , n36285 , n36286 , n36287 , n36288 , n36289 , n36290 , n36291 , n36292 ,
     n36293 , n36294 , n36295 , n36296 , n36297 , n36298 , n36299 , n36300 , n36301 , n36302 ,
     n36303 , n36304 , n36305 , n36306 , n36307 , n36308 , n36309 , n36310 , n36311 , n36312 ,
     n36313 , n36314 , n36315 , n36316 , n36317 , n36318 , n36319 , n36320 , n36321 , n36322 ,
     n36323 , n36324 , n36325 , n36326 , n36327 , n36328 , n36329 , n36330 , n36331 , n36332 ,
     n36333 , n36334 , n36335 , n36336 , n36337 , n36338 , n36339 , n36340 , n36341 , n36342 ,
     n36343 , n36344 , n36345 , n36346 , n36347 , n36348 , n36349 , n36350 , n36351 , n36352 ,
     n36353 , n36354 , n36355 , n36356 , n36357 , n36358 , n36359 , n36360 , n36361 , n36362 ,
     n36363 , n36364 , n36365 , n36366 , n36367 , n36368 , n36369 , n36370 , n36371 , n36372 ,
     n36373 , n36374 , n36375 , n36376 , n36377 , n36378 , n36379 , n36380 , n36381 , n36382 ,
     n36383 , n36384 , n36385 , n36386 , n36387 , n36388 , n36389 , n36390 , n36391 , n36392 ,
     n36393 , n36394 , n36395 , n36396 , n36397 , n36398 , n36399 , n36400 , n36401 , n36402 ,
     n36403 , n36404 , n36405 , n36406 , n36407 , n36408 , n36409 , n36410 , n36411 , n36412 ,
     n36413 , n36414 , n36415 , n36416 , n36417 , n36418 , n36419 , n36420 , n36421 , n36422 ,
     n36423 , n36424 , n36425 , n36426 , n36427 , n36428 , n36429 , n36430 , n36431 , n36432 ,
     n36433 , n36434 , n36435 , n36436 , n36437 , n36438 , n36439 , n36440 , n36441 , n36442 ,
     n36443 , n36444 , n36445 , n36446 , n36447 , n36448 , n36449 , n36450 , n36451 , n36452 ,
     n36453 , n36454 , n36455 , n36456 , n36457 , n36458 , n36459 , n36460 , n36461 , n36462 ,
     n36463 , n36464 , n36465 , n36466 , n36467 , n36468 , n36469 , n36470 , n36471 , n36472 ,
     n36473 , n36474 , n36475 , n36476 , n36477 , n36478 , n36479 , n36480 , n36481 , n36482 ,
     n36483 , n36484 , n36485 , n36486 , n36487 , n36488 , n36489 , n36490 , n36491 , n36492 ,
     n36493 , n36494 , n36495 , n36496 , n36497 , n36498 , n36499 , n36500 , n36501 , n36502 ,
     n36503 , n36504 , n36505 , n36506 , n36507 , n36508 , n36509 , n36510 , n36511 , n36512 ,
     n36513 , n36514 , n36515 , n36516 , n36517 , n36518 , n36519 , n36520 , n36521 , n36522 ,
     n36523 , n36524 , n36525 , n36526 , n36527 , n36528 , n36529 , n36530 , n36531 , n36532 ,
     n36533 , n36534 , n36535 , n36536 , n36537 , n36538 , n36539 , n36540 , n36541 , n36542 ,
     n36543 , n36544 , n36545 , n36546 , n36547 , n36548 , n36549 , n36550 , n36551 , n36552 ,
     n36553 , n36554 , n36555 , n36556 , n36557 , n36558 , n36559 , n36560 , n36561 , n36562 ,
     n36563 , n36564 , n36565 , n36566 , n36567 , n36568 , n36569 , n36570 , n36571 , n36572 ,
     n36573 , n36574 , n36575 , n36576 , n36577 , n36578 , n36579 , n36580 , n36581 , n36582 ,
     n36583 , n36584 , n36585 , n36586 , n36587 , n36588 , n36589 , n36590 , n36591 , n36592 ,
     n36593 , n36594 , n36595 , n36596 , n36597 , n36598 , n36599 , n36600 , n36601 , n36602 ,
     n36603 , n36604 , n36605 , n36606 , n36607 , n36608 , n36609 , n36610 , n36611 , n36612 ,
     n36613 , n36614 , n36615 , n36616 , n36617 , n36618 , n36619 , n36620 , n36621 , n36622 ,
     n36623 , n36624 , n36625 , n36626 , n36627 , n36628 , n36629 , n36630 , n36631 , n36632 ,
     n36633 , n36634 , n36635 , n36636 , n36637 , n36638 , n36639 , n36640 , n36641 , n36642 ,
     n36643 , n36644 , n36645 , n36646 , n36647 , n36648 , n36649 , n36650 , n36651 , n36652 ,
     n36653 , n36654 , n36655 , n36656 , n36657 , n36658 , n36659 , n36660 , n36661 , n36662 ,
     n36663 , n36664 , n36665 , n36666 , n36667 , n36668 , n36669 , n36670 , n36671 , n36672 ,
     n36673 , n36674 , n36675 , n36676 , n36677 , n36678 , n36679 , n36680 , n36681 , n36682 ,
     n36683 , n36684 , n36685 , n36686 , n36687 , n36688 , n36689 , n36690 , n36691 , n36692 ,
     n36693 , n36694 , n36695 , n36696 , n36697 , n36698 , n36699 , n36700 , n36701 , n36702 ,
     n36703 , n36704 , n36705 , n36706 , n36707 , n36708 , n36709 , n36710 , n36711 , n36712 ,
     n36713 , n36714 , n36715 , n36716 , n36717 , n36718 , n36719 , n36720 , n36721 , n36722 ,
     n36723 , n36724 , n36725 , n36726 , n36727 , n36728 , n36729 , n36730 , n36731 , n36732 ,
     n36733 , n36734 , n36735 , n36736 , n36737 , n36738 , n36739 , n36740 , n36741 , n36742 ,
     n36743 , n36744 , n36745 , n36746 , n36747 , n36748 , n36749 , n36750 , n36751 , n36752 ,
     n36753 , n36754 , n36755 , n36756 , n36757 , n36758 , n36759 , n36760 , n36761 , n36762 ,
     n36763 , n36764 , n36765 , n36766 , n36767 , n36768 , n36769 , n36770 , n36771 , n36772 ,
     n36773 , n36774 , n36775 , n36776 , n36777 , n36778 , n36779 , n36780 , n36781 , n36782 ,
     n36783 , n36784 , n36785 , n36786 , n36787 , n36788 , n36789 , n36790 , n36791 , n36792 ,
     n36793 , n36794 , n36795 , n36796 , n36797 , n36798 , n36799 , n36800 , n36801 , n36802 ,
     n36803 , n36804 , n36805 , n36806 , n36807 , n36808 , n36809 , n36810 , n36811 , n36812 ,
     n36813 , n36814 , n36815 , n36816 , n36817 , n36818 , n36819 , n36820 , n36821 , n36822 ,
     n36823 , n36824 , n36825 , n36826 , n36827 , n36828 , n36829 , n36830 , n36831 , n36832 ,
     n36833 , n36834 , n36835 , n36836 , n36837 , n36838 , n36839 , n36840 , n36841 , n36842 ,
     n36843 , n36844 , n36845 , n36846 , n36847 , n36848 , n36849 , n36850 , n36851 , n36852 ,
     n36853 , n36854 , n36855 , n36856 , n36857 , n36858 , n36859 , n36860 , n36861 , n36862 ,
     n36863 , n36864 , n36865 , n36866 , n36867 , n36868 , n36869 , n36870 , n36871 , n36872 ,
     n36873 , n36874 , n36875 , n36876 , n36877 , n36878 , n36879 , n36880 , n36881 , n36882 ,
     n36883 , n36884 , n36885 , n36886 , n36887 , n36888 , n36889 , n36890 , n36891 , n36892 ,
     n36893 , n36894 , n36895 , n36896 , n36897 , n36898 , n36899 , n36900 , n36901 , n36902 ,
     n36903 , n36904 , n36905 , n36906 , n36907 , n36908 , n36909 , n36910 , n36911 , n36912 ,
     n36913 , n36914 , n36915 , n36916 , n36917 , n36918 , n36919 , n36920 , n36921 , n36922 ,
     n36923 , n36924 , n36925 , n36926 , n36927 , n36928 , n36929 , n36930 , n36931 , n36932 ,
     n36933 , n36934 , n36935 , n36936 , n36937 , n36938 , n36939 , n36940 , n36941 , n36942 ,
     n36943 , n36944 , n36945 , n36946 , n36947 , n36948 , n36949 , n36950 , n36951 , n36952 ,
     n36953 , n36954 , n36955 , n36956 , n36957 , n36958 , n36959 , n36960 , n36961 , n36962 ,
     n36963 , n36964 , n36965 , n36966 , n36967 , n36968 , n36969 , n36970 , n36971 , n36972 ,
     n36973 , n36974 , n36975 , n36976 , n36977 , n36978 , n36979 , n36980 , n36981 , n36982 ,
     n36983 , n36984 , n36985 , n36986 , n36987 , n36988 , n36989 , n36990 , n36991 , n36992 ,
     n36993 , n36994 , n36995 , n36996 , n36997 , n36998 , n36999 , n37000 , n37001 , n37002 ,
     n37003 , n37004 , n37005 , n37006 , n37007 , n37008 , n37009 , n37010 , n37011 , n37012 ,
     n37013 , n37014 , n37015 , n37016 , n37017 , n37018 , n37019 , n37020 , n37021 , n37022 ,
     n37023 , n37024 , n37025 , n37026 , n37027 , n37028 , n37029 , n37030 , n37031 , n37032 ,
     n37033 , n37034 , n37035 , n37036 , n37037 , n37038 , n37039 , n37040 , n37041 , n37042 ,
     n37043 , n37044 , n37045 , n37046 , n37047 , n37048 , n37049 , n37050 , n37051 , n37052 ,
     n37053 , n37054 , n37055 , n37056 , n37057 , n37058 , n37059 , n37060 , n37061 , n37062 ,
     n37063 , n37064 , n37065 , n37066 , n37067 , n37068 , n37069 , n37070 , n37071 , n37072 ,
     n37073 , n37074 , n37075 , n37076 , n37077 , n37078 , n37079 , n37080 , n37081 , n37082 ,
     n37083 , n37084 , n37085 , n37086 , n37087 , n37088 , n37089 , n37090 , n37091 , n37092 ,
     n37093 , n37094 , n37095 , n37096 , n37097 , n37098 , n37099 , n37100 , n37101 , n37102 ,
     n37103 , n37104 , n37105 , n37106 , n37107 , n37108 , n37109 , n37110 , n37111 , n37112 ,
     n37113 , n37114 , n37115 , n37116 , n37117 , n37118 , n37119 , n37120 , n37121 , n37122 ,
     n37123 , n37124 , n37125 , n37126 , n37127 , n37128 , n37129 , n37130 , n37131 , n37132 ,
     n37133 , n37134 , n37135 , n37136 , n37137 , n37138 , n37139 , n37140 , n37141 , n37142 ,
     n37143 , n37144 , n37145 , n37146 , n37147 , n37148 , n37149 , n37150 , n37151 , n37152 ,
     n37153 , n37154 , n37155 , n37156 , n37157 , n37158 , n37159 , n37160 , n37161 , n37162 ,
     n37163 , n37164 , n37165 , n37166 , n37167 , n37168 , n37169 , n37170 , n37171 , n37172 ,
     n37173 , n37174 , n37175 , n37176 , n37177 , n37178 , n37179 , n37180 , n37181 , n37182 ,
     n37183 , n37184 , n37185 , n37186 , n37187 , n37188 , n37189 , n37190 , n37191 , n37192 ,
     n37193 , n37194 , n37195 , n37196 , n37197 , n37198 , n37199 , n37200 , n37201 , n37202 ,
     n37203 , n37204 , n37205 , n37206 , n37207 , n37208 , n37209 , n37210 , n37211 , n37212 ,
     n37213 , n37214 , n37215 , n37216 , n37217 , n37218 , n37219 , n37220 , n37221 , n37222 ,
     n37223 , n37224 , n37225 , n37226 , n37227 , n37228 , n37229 , n37230 , n37231 , n37232 ,
     n37233 , n37234 , n37235 , n37236 , n37237 , n37238 , n37239 , n37240 , n37241 , n37242 ,
     n37243 , n37244 , n37245 , n37246 , n37247 , n37248 , n37249 , n37250 , n37251 , n37252 ,
     n37253 , n37254 , n37255 , n37256 , n37257 , n37258 , n37259 , n37260 , n37261 , n37262 ,
     n37263 , n37264 , n37265 , n37266 , n37267 , n37268 , n37269 , n37270 , n37271 , n37272 ,
     n37273 , n37274 , n37275 , n37276 , n37277 , n37278 , n37279 , n37280 , n37281 , n37282 ,
     n37283 , n37284 , n37285 , n37286 , n37287 , n37288 , n37289 , n37290 , n37291 , n37292 ,
     n37293 , n37294 , n37295 , n37296 , n37297 , n37298 , n37299 , n37300 , n37301 , n37302 ,
     n37303 , n37304 , n37305 , n37306 , n37307 , n37308 , n37309 , n37310 , n37311 , n37312 ,
     n37313 , n37314 , n37315 , n37316 , n37317 , n37318 , n37319 , n37320 , n37321 , n37322 ,
     n37323 , n37324 , n37325 , n37326 , n37327 , n37328 , n37329 , n37330 , n37331 , n37332 ,
     n37333 , n37334 , n37335 , n37336 , n37337 , n37338 , n37339 , n37340 , n37341 , n37342 ,
     n37343 , n37344 , n37345 , n37346 , n37347 , n37348 , n37349 , n37350 , n37351 , n37352 ,
     n37353 , n37354 , n37355 , n37356 , n37357 , n37358 , n37359 , n37360 , n37361 , n37362 ,
     n37363 , n37364 , n37365 , n37366 , n37367 , n37368 , n37369 , n37370 , n37371 , n37372 ,
     n37373 , n37374 , n37375 , n37376 , n37377 , n37378 , n37379 , n37380 , n37381 , n37382 ,
     n37383 , n37384 , n37385 , n37386 , n37387 , n37388 , n37389 , n37390 , n37391 , n37392 ,
     n37393 , n37394 , n37395 , n37396 , n37397 , n37398 , n37399 , n37400 , n37401 , n37402 ,
     n37403 , n37404 , n37405 , n37406 , n37407 , n37408 , n37409 , n37410 , n37411 , n37412 ,
     n37413 , n37414 , n37415 , n37416 , n37417 , n37418 , n37419 , n37420 , n37421 , n37422 ,
     n37423 , n37424 , n37425 , n37426 , n37427 , n37428 , n37429 , n37430 , n37431 , n37432 ,
     n37433 , n37434 , n37435 , n37436 , n37437 , n37438 , n37439 , n37440 , n37441 , n37442 ,
     n37443 , n37444 , n37445 , n37446 , n37447 , n37448 , n37449 , n37450 , n37451 , n37452 ,
     n37453 , n37454 , n37455 , n37456 , n37457 , n37458 , n37459 , n37460 , n37461 , n37462 ,
     n37463 , n37464 , n37465 , n37466 , n37467 , n37468 , n37469 , n37470 , n37471 , n37472 ,
     n37473 , n37474 , n37475 , n37476 , n37477 , n37478 , n37479 , n37480 , n37481 , n37482 ,
     n37483 , n37484 , n37485 , n37486 , n37487 , n37488 , n37489 , n37490 , n37491 , n37492 ,
     n37493 , n37494 , n37495 , n37496 , n37497 , n37498 , n37499 , n37500 , n37501 , n37502 ,
     n37503 , n37504 , n37505 , n37506 , n37507 , n37508 , n37509 , n37510 , n37511 , n37512 ,
     n37513 , n37514 , n37515 , n37516 , n37517 , n37518 , n37519 , n37520 , n37521 , n37522 ,
     n37523 , n37524 , n37525 , n37526 , n37527 , n37528 , n37529 , n37530 , n37531 , n37532 ,
     n37533 , n37534 , n37535 , n37536 , n37537 , n37538 , n37539 , n37540 , n37541 , n37542 ,
     n37543 , n37544 , n37545 , n37546 , n37547 , n37548 , n37549 , n37550 , n37551 , n37552 ,
     n37553 , n37554 , n37555 , n37556 , n37557 , n37558 , n37559 , n37560 , n37561 , n37562 ,
     n37563 , n37564 , n37565 , n37566 , n37567 , n37568 , n37569 , n37570 , n37571 , n37572 ,
     n37573 , n37574 , n37575 , n37576 , n37577 , n37578 , n37579 , n37580 , n37581 , n37582 ,
     n37583 , n37584 , n37585 , n37586 , n37587 , n37588 , n37589 , n37590 , n37591 , n37592 ,
     n37593 , n37594 , n37595 , n37596 , n37597 , n37598 , n37599 , n37600 , n37601 , n37602 ,
     n37603 , n37604 , n37605 , n37606 , n37607 , n37608 , n37609 , n37610 , n37611 , n37612 ,
     n37613 , n37614 , n37615 , n37616 , n37617 , n37618 , n37619 , n37620 , n37621 , n37622 ,
     n37623 , n37624 , n37625 , n37626 , n37627 , n37628 , n37629 , n37630 , n37631 , n37632 ,
     n37633 , n37634 , n37635 , n37636 , n37637 , n37638 , n37639 , n37640 , n37641 , n37642 ,
     n37643 , n37644 , n37645 , n37646 , n37647 , n37648 , n37649 , n37650 , n37651 , n37652 ,
     n37653 , n37654 , n37655 , n37656 , n37657 , n37658 , n37659 , n37660 , n37661 , n37662 ,
     n37663 , n37664 , n37665 , n37666 , n37667 , n37668 , n37669 , n37670 , n37671 , n37672 ,
     n37673 , n37674 , n37675 , n37676 , n37677 , n37678 , n37679 , n37680 , n37681 , n37682 ,
     n37683 , n37684 , n37685 , n37686 , n37687 , n37688 , n37689 , n37690 , n37691 , n37692 ,
     n37693 , n37694 , n37695 , n37696 , n37697 , n37698 , n37699 , n37700 , n37701 , n37702 ,
     n37703 , n37704 , n37705 , n37706 , n37707 , n37708 , n37709 , n37710 , n37711 , n37712 ,
     n37713 , n37714 , n37715 , n37716 , n37717 , n37718 , n37719 , n37720 , n37721 , n37722 ,
     n37723 , n37724 , n37725 , n37726 , n37727 , n37728 , n37729 , n37730 , n37731 , n37732 ,
     n37733 , n37734 , n37735 , n37736 , n37737 , n37738 , n37739 , n37740 , n37741 , n37742 ,
     n37743 , n37744 , n37745 , n37746 , n37747 , n37748 , n37749 , n37750 , n37751 , n37752 ,
     n37753 , n37754 , n37755 , n37756 , n37757 , n37758 , n37759 , n37760 , n37761 , n37762 ,
     n37763 , n37764 , n37765 , n37766 , n37767 , n37768 , n37769 , n37770 , n37771 , n37772 ,
     n37773 , n37774 , n37775 , n37776 , n37777 , n37778 , n37779 , n37780 , n37781 , n37782 ,
     n37783 , n37784 , n37785 , n37786 , n37787 , n37788 , n37789 , n37790 , n37791 , n37792 ,
     n37793 , n37794 , n37795 , n37796 , n37797 , n37798 , n37799 , n37800 , n37801 , n37802 ,
     n37803 , n37804 , n37805 , n37806 , n37807 , n37808 , n37809 , n37810 , n37811 , n37812 ,
     n37813 , n37814 , n37815 , n37816 , n37817 , n37818 , n37819 , n37820 , n37821 , n37822 ,
     n37823 , n37824 , n37825 , n37826 , n37827 , n37828 , n37829 , n37830 , n37831 , n37832 ,
     n37833 , n37834 , n37835 , n37836 , n37837 , n37838 , n37839 , n37840 , n37841 , n37842 ,
     n37843 , n37844 , n37845 , n37846 , n37847 , n37848 , n37849 , n37850 , n37851 , n37852 ,
     n37853 , n37854 , n37855 , n37856 , n37857 , n37858 , n37859 , n37860 , n37861 , n37862 ,
     n37863 , n37864 , n37865 , n37866 , n37867 , n37868 , n37869 , n37870 , n37871 , n37872 ,
     n37873 , n37874 , n37875 , n37876 , n37877 , n37878 , n37879 , n37880 , n37881 , n37882 ,
     n37883 , n37884 , n37885 , n37886 , n37887 , n37888 , n37889 , n37890 , n37891 , n37892 ,
     n37893 , n37894 , n37895 , n37896 , n37897 , n37898 , n37899 , n37900 , n37901 , n37902 ,
     n37903 , n37904 , n37905 , n37906 , n37907 , n37908 , n37909 , n37910 , n37911 , n37912 ,
     n37913 , n37914 , n37915 , n37916 , n37917 , n37918 , n37919 , n37920 , n37921 , n37922 ,
     n37923 , n37924 , n37925 , n37926 , n37927 , n37928 , n37929 , n37930 , n37931 , n37932 ,
     n37933 , n37934 , n37935 , n37936 , n37937 , n37938 , n37939 , n37940 , n37941 , n37942 ,
     n37943 , n37944 , n37945 , n37946 , n37947 , n37948 , n37949 , n37950 , n37951 , n37952 ,
     n37953 , n37954 , n37955 , n37956 , n37957 , n37958 , n37959 , n37960 , n37961 , n37962 ,
     n37963 , n37964 , n37965 , n37966 , n37967 , n37968 , n37969 , n37970 , n37971 , n37972 ,
     n37973 , n37974 , n37975 , n37976 , n37977 , n37978 , n37979 , n37980 , n37981 , n37982 ,
     n37983 , n37984 , n37985 , n37986 , n37987 , n37988 , n37989 , n37990 , n37991 , n37992 ,
     n37993 , n37994 , n37995 , n37996 , n37997 , n37998 , n37999 , n38000 , n38001 , n38002 ,
     n38003 , n38004 , n38005 , n38006 , n38007 , n38008 , n38009 , n38010 , n38011 , n38012 ,
     n38013 , n38014 , n38015 , n38016 , n38017 , n38018 , n38019 , n38020 , n38021 , n38022 ,
     n38023 , n38024 , n38025 , n38026 , n38027 , n38028 , n38029 , n38030 , n38031 , n38032 ,
     n38033 , n38034 , n38035 , n38036 , n38037 , n38038 , n38039 , n38040 , n38041 , n38042 ,
     n38043 , n38044 , n38045 , n38046 , n38047 , n38048 , n38049 , n38050 , n38051 , n38052 ,
     n38053 , n38054 , n38055 , n38056 , n38057 , n38058 , n38059 , n38060 , n38061 , n38062 ,
     n38063 , n38064 , n38065 , n38066 , n38067 , n38068 , n38069 , n38070 , n38071 , n38072 ,
     n38073 , n38074 , n38075 , n38076 , n38077 , n38078 , n38079 , n38080 , n38081 , n38082 ,
     n38083 , n38084 , n38085 , n38086 , n38087 , n38088 , n38089 , n38090 , n38091 , n38092 ,
     n38093 , n38094 , n38095 , n38096 , n38097 , n38098 , n38099 , n38100 , n38101 , n38102 ,
     n38103 , n38104 , n38105 , n38106 , n38107 , n38108 , n38109 , n38110 , n38111 , n38112 ,
     n38113 , n38114 , n38115 , n38116 , n38117 , n38118 , n38119 , n38120 , n38121 , n38122 ,
     n38123 , n38124 , n38125 , n38126 , n38127 , n38128 , n38129 , n38130 , n38131 , n38132 ,
     n38133 , n38134 , n38135 , n38136 , n38137 , n38138 , n38139 , n38140 , n38141 , n38142 ,
     n38143 , n38144 , n38145 , n38146 , n38147 , n38148 , n38149 , n38150 , n38151 , n38152 ,
     n38153 , n38154 , n38155 , n38156 , n38157 , n38158 , n38159 , n38160 , n38161 , n38162 ,
     n38163 , n38164 , n38165 , n38166 , n38167 , n38168 , n38169 , n38170 , n38171 , n38172 ,
     n38173 , n38174 , n38175 , n38176 , n38177 , n38178 , n38179 , n38180 , n38181 , n38182 ,
     n38183 , n38184 , n38185 , n38186 , n38187 , n38188 , n38189 , n38190 , n38191 , n38192 ,
     n38193 , n38194 , n38195 , n38196 , n38197 , n38198 , n38199 , n38200 , n38201 , n38202 ,
     n38203 , n38204 , n38205 , n38206 , n38207 , n38208 , n38209 , n38210 , n38211 , n38212 ,
     n38213 , n38214 , n38215 , n38216 , n38217 , n38218 , n38219 , n38220 , n38221 , n38222 ,
     n38223 , n38224 , n38225 , n38226 , n38227 , n38228 , n38229 , n38230 , n38231 , n38232 ,
     n38233 , n38234 , n38235 , n38236 , n38237 , n38238 , n38239 , n38240 , n38241 , n38242 ,
     n38243 , n38244 , n38245 , n38246 , n38247 , n38248 , n38249 , n38250 , n38251 , n38252 ,
     n38253 , n38254 , n38255 , n38256 , n38257 , n38258 , n38259 , n38260 , n38261 , n38262 ,
     n38263 , n38264 , n38265 , n38266 , n38267 , n38268 , n38269 , n38270 , n38271 , n38272 ,
     n38273 , n38274 , n38275 , n38276 , n38277 , n38278 , n38279 , n38280 , n38281 , n38282 ,
     n38283 , n38284 , n38285 , n38286 , n38287 , n38288 , n38289 , n38290 , n38291 , n38292 ,
     n38293 , n38294 , n38295 , n38296 , n38297 , n38298 , n38299 , n38300 , n38301 , n38302 ,
     n38303 , n38304 , n38305 , n38306 , n38307 , n38308 , n38309 , n38310 , n38311 , n38312 ,
     n38313 , n38314 , n38315 , n38316 , n38317 , n38318 , n38319 , n38320 , n38321 , n38322 ,
     n38323 , n38324 , n38325 , n38326 , n38327 , n38328 , n38329 , n38330 , n38331 , n38332 ,
     n38333 , n38334 , n38335 , n38336 , n38337 , n38338 , n38339 , n38340 , n38341 , n38342 ,
     n38343 , n38344 , n38345 , n38346 , n38347 , n38348 , n38349 , n38350 , n38351 , n38352 ,
     n38353 , n38354 , n38355 , n38356 , n38357 , n38358 , n38359 , n38360 , n38361 , n38362 ,
     n38363 , n38364 , n38365 , n38366 , n38367 , n38368 , n38369 , n38370 , n38371 , n38372 ,
     n38373 , n38374 , n38375 , n38376 , n38377 , n38378 , n38379 , n38380 , n38381 , n38382 ,
     n38383 , n38384 , n38385 , n38386 , n38387 , n38388 , n38389 , n38390 , n38391 , n38392 ,
     n38393 , n38394 , n38395 , n38396 , n38397 , n38398 , n38399 , n38400 , n38401 , n38402 ,
     n38403 , n38404 , n38405 , n38406 , n38407 , n38408 , n38409 , n38410 , n38411 , n38412 ,
     n38413 , n38414 , n38415 , n38416 , n38417 , n38418 , n38419 , n38420 , n38421 , n38422 ,
     n38423 , n38424 , n38425 , n38426 , n38427 , n38428 , n38429 , n38430 , n38431 , n38432 ,
     n38433 , n38434 , n38435 , n38436 , n38437 , n38438 , n38439 , n38440 , n38441 , n38442 ,
     n38443 , n38444 , n38445 , n38446 , n38447 , n38448 , n38449 , n38450 , n38451 , n38452 ,
     n38453 , n38454 , n38455 , n38456 , n38457 , n38458 , n38459 , n38460 , n38461 , n38462 ,
     n38463 , n38464 , n38465 , n38466 , n38467 , n38468 , n38469 , n38470 , n38471 , n38472 ,
     n38473 , n38474 , n38475 , n38476 , n38477 , n38478 , n38479 , n38480 , n38481 , n38482 ,
     n38483 , n38484 , n38485 , n38486 , n38487 , n38488 , n38489 , n38490 , n38491 , n38492 ,
     n38493 , n38494 , n38495 , n38496 , n38497 , n38498 , n38499 , n38500 , n38501 , n38502 ,
     n38503 , n38504 , n38505 , n38506 , n38507 , n38508 , n38509 , n38510 , n38511 , n38512 ,
     n38513 , n38514 , n38515 , n38516 , n38517 , n38518 , n38519 , n38520 , n38521 , n38522 ,
     n38523 , n38524 , n38525 , n38526 , n38527 , n38528 , n38529 , n38530 , n38531 , n38532 ,
     n38533 , n38534 , n38535 , n38536 , n38537 , n38538 , n38539 , n38540 , n38541 , n38542 ,
     n38543 , n38544 , n38545 , n38546 , n38547 , n38548 , n38549 , n38550 , n38551 , n38552 ,
     n38553 , n38554 , n38555 , n38556 , n38557 , n38558 , n38559 , n38560 , n38561 , n38562 ,
     n38563 , n38564 , n38565 , n38566 , n38567 , n38568 , n38569 , n38570 , n38571 , n38572 ,
     n38573 , n38574 , n38575 , n38576 , n38577 , n38578 , n38579 , n38580 , n38581 , n38582 ,
     n38583 , n38584 , n38585 , n38586 , n38587 , n38588 , n38589 , n38590 , n38591 , n38592 ,
     n38593 , n38594 , n38595 , n38596 , n38597 , n38598 , n38599 , n38600 , n38601 , n38602 ,
     n38603 , n38604 , n38605 , n38606 , n38607 , n38608 , n38609 , n38610 , n38611 , n38612 ,
     n38613 , n38614 , n38615 , n38616 , n38617 , n38618 , n38619 , n38620 , n38621 , n38622 ,
     n38623 , n38624 , n38625 , n38626 , n38627 , n38628 , n38629 , n38630 , n38631 , n38632 ,
     n38633 , n38634 , n38635 , n38636 , n38637 , n38638 , n38639 , n38640 , n38641 , n38642 ,
     n38643 , n38644 , n38645 , n38646 , n38647 , n38648 , n38649 , n38650 , n38651 , n38652 ,
     n38653 , n38654 , n38655 , n38656 , n38657 , n38658 , n38659 , n38660 , n38661 , n38662 ,
     n38663 , n38664 , n38665 , n38666 , n38667 , n38668 , n38669 , n38670 , n38671 , n38672 ,
     n38673 , n38674 , n38675 , n38676 , n38677 , n38678 , n38679 , n38680 , n38681 , n38682 ,
     n38683 , n38684 , n38685 , n38686 , n38687 , n38688 , n38689 , n38690 , n38691 , n38692 ,
     n38693 , n38694 , n38695 , n38696 , n38697 , n38698 , n38699 , n38700 , n38701 , n38702 ,
     n38703 , n38704 , n38705 , n38706 , n38707 , n38708 , n38709 , n38710 , n38711 , n38712 ,
     n38713 , n38714 , n38715 , n38716 , n38717 , n38718 , n38719 , n38720 , n38721 , n38722 ,
     n38723 , n38724 , n38725 , n38726 , n38727 , n38728 , n38729 , n38730 , n38731 , n38732 ,
     n38733 , n38734 , n38735 , n38736 , n38737 , n38738 , n38739 , n38740 , n38741 , n38742 ,
     n38743 , n38744 , n38745 , n38746 , n38747 , n38748 , n38749 , n38750 , n38751 , n38752 ,
     n38753 , n38754 , n38755 , n38756 , n38757 , n38758 , n38759 , n38760 , n38761 , n38762 ,
     n38763 , n38764 , n38765 , n38766 , n38767 , n38768 , n38769 , n38770 , n38771 , n38772 ,
     n38773 , n38774 , n38775 , n38776 , n38777 , n38778 , n38779 , n38780 , n38781 , n38782 ,
     n38783 , n38784 , n38785 , n38786 , n38787 , n38788 , n38789 , n38790 , n38791 , n38792 ,
     n38793 , n38794 , n38795 , n38796 , n38797 , n38798 , n38799 , n38800 , n38801 , n38802 ,
     n38803 , n38804 , n38805 , n38806 , n38807 , n38808 , n38809 , n38810 , n38811 , n38812 ,
     n38813 , n38814 , n38815 , n38816 , n38817 , n38818 , n38819 , n38820 , n38821 , n38822 ,
     n38823 , n38824 , n38825 , n38826 , n38827 , n38828 , n38829 , n38830 , n38831 , n38832 ,
     n38833 , n38834 , n38835 , n38836 , n38837 , n38838 , n38839 , n38840 , n38841 , n38842 ,
     n38843 , n38844 , n38845 , n38846 , n38847 , n38848 , n38849 , n38850 , n38851 , n38852 ,
     n38853 , n38854 , n38855 , n38856 , n38857 , n38858 , n38859 , n38860 , n38861 , n38862 ,
     n38863 , n38864 , n38865 , n38866 , n38867 , n38868 , n38869 , n38870 , n38871 , n38872 ,
     n38873 , n38874 , n38875 , n38876 , n38877 , n38878 , n38879 , n38880 , n38881 , n38882 ,
     n38883 , n38884 , n38885 , n38886 , n38887 , n38888 , n38889 , n38890 , n38891 , n38892 ,
     n38893 , n38894 , n38895 , n38896 , n38897 , n38898 , n38899 , n38900 , n38901 , n38902 ,
     n38903 , n38904 , n38905 , n38906 , n38907 , n38908 , n38909 , n38910 , n38911 , n38912 ,
     n38913 , n38914 , n38915 , n38916 , n38917 , n38918 , n38919 , n38920 , n38921 , n38922 ,
     n38923 , n38924 , n38925 , n38926 , n38927 , n38928 , n38929 , n38930 , n38931 , n38932 ,
     n38933 , n38934 , n38935 , n38936 , n38937 , n38938 , n38939 , n38940 , n38941 , n38942 ,
     n38943 , n38944 , n38945 , n38946 , n38947 , n38948 , n38949 , n38950 , n38951 , n38952 ,
     n38953 , n38954 , n38955 , n38956 , n38957 , n38958 , n38959 , n38960 , n38961 , n38962 ,
     n38963 , n38964 , n38965 , n38966 , n38967 , n38968 , n38969 , n38970 , n38971 , n38972 ,
     n38973 , n38974 , n38975 , n38976 , n38977 , n38978 , n38979 , n38980 , n38981 , n38982 ,
     n38983 , n38984 , n38985 , n38986 , n38987 , n38988 , n38989 , n38990 , n38991 , n38992 ,
     n38993 , n38994 , n38995 , n38996 , n38997 , n38998 , n38999 , n39000 , n39001 , n39002 ,
     n39003 , n39004 , n39005 , n39006 , n39007 , n39008 , n39009 , n39010 , n39011 , n39012 ,
     n39013 , n39014 , n39015 , n39016 , n39017 , n39018 , n39019 , n39020 , n39021 , n39022 ,
     n39023 , n39024 , n39025 , n39026 , n39027 , n39028 , n39029 , n39030 , n39031 , n39032 ,
     n39033 , n39034 , n39035 , n39036 , n39037 , n39038 , n39039 , n39040 , n39041 , n39042 ,
     n39043 , n39044 , n39045 , n39046 , n39047 , n39048 , n39049 , n39050 , n39051 , n39052 ,
     n39053 , n39054 , n39055 , n39056 , n39057 , n39058 , n39059 , n39060 , n39061 , n39062 ,
     n39063 , n39064 , n39065 , n39066 , n39067 , n39068 , n39069 , n39070 , n39071 , n39072 ,
     n39073 , n39074 , n39075 , n39076 , n39077 , n39078 , n39079 , n39080 , n39081 , n39082 ,
     n39083 , n39084 , n39085 , n39086 , n39087 , n39088 , n39089 , n39090 , n39091 , n39092 ,
     n39093 , n39094 , n39095 , n39096 , n39097 , n39098 , n39099 , n39100 , n39101 , n39102 ,
     n39103 , n39104 , n39105 , n39106 , n39107 , n39108 , n39109 , n39110 , n39111 , n39112 ,
     n39113 , n39114 , n39115 , n39116 , n39117 , n39118 , n39119 , n39120 , n39121 , n39122 ,
     n39123 , n39124 , n39125 , n39126 , n39127 , n39128 , n39129 , n39130 , n39131 , n39132 ,
     n39133 , n39134 , n39135 , n39136 , n39137 , n39138 , n39139 , n39140 , n39141 , n39142 ,
     n39143 , n39144 , n39145 , n39146 , n39147 , n39148 , n39149 , n39150 , n39151 , n39152 ,
     n39153 , n39154 , n39155 , n39156 , n39157 , n39158 , n39159 , n39160 , n39161 , n39162 ,
     n39163 , n39164 , n39165 , n39166 , n39167 , n39168 , n39169 , n39170 , n39171 , n39172 ,
     n39173 , n39174 , n39175 , n39176 , n39177 , n39178 , n39179 , n39180 , n39181 , n39182 ,
     n39183 , n39184 , n39185 , n39186 , n39187 , n39188 , n39189 , n39190 , n39191 , n39192 ,
     n39193 , n39194 , n39195 , n39196 , n39197 , n39198 , n39199 , n39200 , n39201 , n39202 ,
     n39203 , n39204 , n39205 , n39206 , n39207 , n39208 , n39209 , n39210 , n39211 , n39212 ,
     n39213 , n39214 , n39215 , n39216 , n39217 , n39218 , n39219 , n39220 , n39221 , n39222 ,
     n39223 , n39224 , n39225 , n39226 , n39227 , n39228 , n39229 , n39230 , n39231 , n39232 ,
     n39233 , n39234 , n39235 , n39236 , n39237 , n39238 , n39239 , n39240 , n39241 , n39242 ,
     n39243 , n39244 , n39245 , n39246 , n39247 , n39248 , n39249 , n39250 , n39251 , n39252 ,
     n39253 , n39254 , n39255 , n39256 , n39257 , n39258 , n39259 , n39260 , n39261 , n39262 ,
     n39263 , n39264 , n39265 , n39266 , n39267 , n39268 , n39269 , n39270 , n39271 , n39272 ,
     n39273 , n39274 , n39275 , n39276 , n39277 , n39278 , n39279 , n39280 , n39281 , n39282 ,
     n39283 , n39284 , n39285 , n39286 , n39287 , n39288 , n39289 , n39290 , n39291 , n39292 ,
     n39293 , n39294 , n39295 , n39296 , n39297 , n39298 , n39299 , n39300 , n39301 , n39302 ,
     n39303 , n39304 , n39305 , n39306 , n39307 , n39308 , n39309 , n39310 , n39311 , n39312 ,
     n39313 , n39314 , n39315 , n39316 , n39317 , n39318 , n39319 , n39320 , n39321 , n39322 ,
     n39323 , n39324 , n39325 , n39326 , n39327 , n39328 , n39329 , n39330 , n39331 , n39332 ,
     n39333 , n39334 , n39335 , n39336 , n39337 , n39338 , n39339 , n39340 , n39341 , n39342 ,
     n39343 , n39344 , n39345 , n39346 , n39347 , n39348 , n39349 , n39350 , n39351 , n39352 ,
     n39353 , n39354 , n39355 , n39356 , n39357 , n39358 , n39359 , n39360 , n39361 , n39362 ,
     n39363 , n39364 , n39365 , n39366 , n39367 , n39368 , n39369 , n39370 , n39371 , n39372 ,
     n39373 , n39374 , n39375 , n39376 , n39377 , n39378 , n39379 , n39380 , n39381 , n39382 ,
     n39383 , n39384 , n39385 , n39386 , n39387 , n39388 , n39389 , n39390 , n39391 , n39392 ,
     n39393 , n39394 , n39395 , n39396 , n39397 , n39398 , n39399 , n39400 , n39401 , n39402 ,
     n39403 , n39404 , n39405 , n39406 , n39407 , n39408 , n39409 , n39410 , n39411 , n39412 ,
     n39413 , n39414 , n39415 , n39416 , n39417 , n39418 , n39419 , n39420 , n39421 , n39422 ,
     n39423 , n39424 , n39425 , n39426 , n39427 , n39428 , n39429 , n39430 , n39431 , n39432 ,
     n39433 , n39434 , n39435 , n39436 , n39437 , n39438 , n39439 , n39440 , n39441 , n39442 ,
     n39443 , n39444 , n39445 , n39446 , n39447 , n39448 , n39449 , n39450 , n39451 , n39452 ,
     n39453 , n39454 , n39455 , n39456 , n39457 , n39458 , n39459 , n39460 , n39461 , n39462 ,
     n39463 , n39464 , n39465 , n39466 , n39467 , n39468 , n39469 , n39470 , n39471 , n39472 ,
     n39473 , n39474 , n39475 , n39476 , n39477 , n39478 , n39479 , n39480 , n39481 , n39482 ,
     n39483 , n39484 , n39485 , n39486 , n39487 , n39488 , n39489 , n39490 , n39491 , n39492 ,
     n39493 , n39494 , n39495 , n39496 , n39497 , n39498 , n39499 , n39500 , n39501 , n39502 ,
     n39503 , n39504 , n39505 , n39506 , n39507 , n39508 , n39509 , n39510 , n39511 , n39512 ,
     n39513 , n39514 , n39515 , n39516 , n39517 , n39518 , n39519 , n39520 , n39521 , n39522 ,
     n39523 , n39524 , n39525 , n39526 , n39527 , n39528 , n39529 , n39530 , n39531 , n39532 ,
     n39533 , n39534 , n39535 , n39536 , n39537 , n39538 , n39539 , n39540 , n39541 , n39542 ,
     n39543 , n39544 , n39545 , n39546 , n39547 , n39548 , n39549 , n39550 , n39551 , n39552 ,
     n39553 , n39554 , n39555 , n39556 , n39557 , n39558 , n39559 , n39560 , n39561 , n39562 ,
     n39563 , n39564 , n39565 , n39566 , n39567 , n39568 , n39569 , n39570 , n39571 , n39572 ,
     n39573 , n39574 , n39575 , n39576 , n39577 , n39578 , n39579 , n39580 , n39581 , n39582 ,
     n39583 , n39584 , n39585 , n39586 , n39587 , n39588 , n39589 , n39590 , n39591 , n39592 ,
     n39593 , n39594 , n39595 , n39596 , n39597 , n39598 , n39599 , n39600 , n39601 , n39602 ,
     n39603 , n39604 , n39605 , n39606 , n39607 , n39608 , n39609 , n39610 , n39611 , n39612 ,
     n39613 , n39614 , n39615 , n39616 , n39617 , n39618 , n39619 , n39620 , n39621 , n39622 ,
     n39623 , n39624 , n39625 , n39626 , n39627 , n39628 , n39629 , n39630 , n39631 , n39632 ,
     n39633 , n39634 , n39635 , n39636 , n39637 , n39638 , n39639 , n39640 , n39641 , n39642 ,
     n39643 , n39644 , n39645 , n39646 , n39647 , n39648 , n39649 , n39650 , n39651 , n39652 ,
     n39653 , n39654 , n39655 , n39656 , n39657 , n39658 , n39659 , n39660 , n39661 , n39662 ,
     n39663 , n39664 , n39665 , n39666 , n39667 , n39668 , n39669 , n39670 , n39671 , n39672 ,
     n39673 , n39674 , n39675 , n39676 , n39677 , n39678 , n39679 , n39680 , n39681 , n39682 ,
     n39683 , n39684 , n39685 , n39686 , n39687 , n39688 , n39689 , n39690 , n39691 , n39692 ,
     n39693 , n39694 , n39695 , n39696 , n39697 , n39698 , n39699 , n39700 , n39701 , n39702 ,
     n39703 , n39704 , n39705 , n39706 , n39707 , n39708 , n39709 , n39710 , n39711 , n39712 ,
     n39713 , n39714 , n39715 , n39716 , n39717 , n39718 , n39719 , n39720 , n39721 , n39722 ,
     n39723 , n39724 , n39725 , n39726 , n39727 , n39728 , n39729 , n39730 , n39731 , n39732 ,
     n39733 , n39734 , n39735 , n39736 , n39737 , n39738 , n39739 , n39740 , n39741 , n39742 ,
     n39743 , n39744 , n39745 , n39746 , n39747 , n39748 , n39749 , n39750 , n39751 , n39752 ,
     n39753 , n39754 , n39755 , n39756 , n39757 , n39758 , n39759 , n39760 , n39761 , n39762 ,
     n39763 , n39764 , n39765 , n39766 , n39767 , n39768 , n39769 , n39770 , n39771 , n39772 ,
     n39773 , n39774 , n39775 , n39776 , n39777 , n39778 , n39779 , n39780 , n39781 , n39782 ,
     n39783 , n39784 , n39785 , n39786 , n39787 , n39788 , n39789 , n39790 , n39791 , n39792 ,
     n39793 , n39794 , n39795 , n39796 , n39797 , n39798 , n39799 , n39800 , n39801 , n39802 ,
     n39803 , n39804 , n39805 , n39806 , n39807 , n39808 , n39809 , n39810 , n39811 , n39812 ,
     n39813 , n39814 , n39815 , n39816 , n39817 , n39818 , n39819 , n39820 , n39821 , n39822 ,
     n39823 , n39824 , n39825 , n39826 , n39827 , n39828 , n39829 , n39830 , n39831 , n39832 ,
     n39833 , n39834 , n39835 , n39836 , n39837 , n39838 , n39839 , n39840 , n39841 , n39842 ,
     n39843 , n39844 , n39845 , n39846 , n39847 , n39848 , n39849 , n39850 , n39851 , n39852 ,
     n39853 , n39854 , n39855 , n39856 , n39857 , n39858 , n39859 , n39860 , n39861 , n39862 ,
     n39863 , n39864 , n39865 , n39866 , n39867 , n39868 , n39869 , n39870 , n39871 , n39872 ,
     n39873 , n39874 , n39875 , n39876 , n39877 , n39878 , n39879 , n39880 , n39881 , n39882 ,
     n39883 , n39884 , n39885 , n39886 , n39887 , n39888 , n39889 , n39890 , n39891 , n39892 ,
     n39893 , n39894 , n39895 , n39896 , n39897 , n39898 , n39899 , n39900 , n39901 , n39902 ,
     n39903 , n39904 , n39905 , n39906 , n39907 , n39908 , n39909 , n39910 , n39911 , n39912 ,
     n39913 , n39914 , n39915 , n39916 , n39917 , n39918 , n39919 , n39920 , n39921 , n39922 ,
     n39923 , n39924 , n39925 , n39926 , n39927 , n39928 , n39929 , n39930 , n39931 , n39932 ,
     n39933 , n39934 , n39935 , n39936 , n39937 , n39938 , n39939 , n39940 , n39941 , n39942 ,
     n39943 , n39944 , n39945 , n39946 , n39947 , n39948 , n39949 , n39950 , n39951 , n39952 ,
     n39953 , n39954 , n39955 , n39956 , n39957 , n39958 , n39959 , n39960 , n39961 , n39962 ,
     n39963 , n39964 , n39965 , n39966 , n39967 , n39968 , n39969 , n39970 , n39971 , n39972 ,
     n39973 , n39974 , n39975 , n39976 , n39977 , n39978 , n39979 , n39980 , n39981 , n39982 ,
     n39983 , n39984 , n39985 , n39986 , n39987 , n39988 , n39989 , n39990 , n39991 , n39992 ,
     n39993 , n39994 , n39995 , n39996 , n39997 , n39998 , n39999 , n40000 , n40001 , n40002 ,
     n40003 , n40004 , n40005 , n40006 , n40007 , n40008 , n40009 , n40010 , n40011 , n40012 ,
     n40013 , n40014 , n40015 , n40016 , n40017 , n40018 , n40019 , n40020 , n40021 , n40022 ,
     n40023 , n40024 , n40025 , n40026 , n40027 , n40028 , n40029 , n40030 , n40031 , n40032 ,
     n40033 , n40034 , n40035 , n40036 , n40037 , n40038 , n40039 , n40040 , n40041 , n40042 ,
     n40043 , n40044 , n40045 , n40046 , n40047 , n40048 , n40049 , n40050 , n40051 , n40052 ,
     n40053 , n40054 , n40055 , n40056 , n40057 , n40058 , n40059 , n40060 , n40061 , n40062 ,
     n40063 , n40064 , n40065 , n40066 , n40067 , n40068 , n40069 , n40070 , n40071 , n40072 ,
     n40073 , n40074 , n40075 , n40076 , n40077 , n40078 , n40079 , n40080 , n40081 , n40082 ,
     n40083 , n40084 , n40085 , n40086 , n40087 , n40088 , n40089 , n40090 , n40091 , n40092 ,
     n40093 , n40094 , n40095 , n40096 , n40097 , n40098 , n40099 , n40100 , n40101 , n40102 ,
     n40103 , n40104 , n40105 , n40106 , n40107 , n40108 , n40109 , n40110 , n40111 , n40112 ,
     n40113 , n40114 , n40115 , n40116 , n40117 , n40118 , n40119 , n40120 , n40121 , n40122 ,
     n40123 , n40124 , n40125 , n40126 , n40127 , n40128 , n40129 , n40130 , n40131 , n40132 ,
     n40133 , n40134 , n40135 , n40136 , n40137 , n40138 , n40139 , n40140 , n40141 , n40142 ,
     n40143 , n40144 , n40145 , n40146 , n40147 , n40148 , n40149 , n40150 , n40151 , n40152 ,
     n40153 , n40154 , n40155 , n40156 , n40157 , n40158 , n40159 , n40160 , n40161 , n40162 ,
     n40163 , n40164 , n40165 , n40166 , n40167 , n40168 , n40169 , n40170 , n40171 , n40172 ,
     n40173 , n40174 , n40175 , n40176 , n40177 , n40178 , n40179 , n40180 , n40181 , n40182 ,
     n40183 , n40184 , n40185 , n40186 , n40187 , n40188 , n40189 , n40190 , n40191 , n40192 ,
     n40193 , n40194 , n40195 , n40196 , n40197 , n40198 , n40199 , n40200 , n40201 , n40202 ,
     n40203 , n40204 , n40205 , n40206 , n40207 , n40208 , n40209 , n40210 , n40211 , n40212 ,
     n40213 , n40214 , n40215 , n40216 , n40217 , n40218 , n40219 , n40220 , n40221 , n40222 ,
     n40223 , n40224 , n40225 , n40226 , n40227 , n40228 , n40229 , n40230 , n40231 , n40232 ,
     n40233 , n40234 , n40235 , n40236 , n40237 , n40238 , n40239 , n40240 , n40241 , n40242 ,
     n40243 , n40244 , n40245 , n40246 , n40247 , n40248 , n40249 , n40250 , n40251 , n40252 ,
     n40253 , n40254 , n40255 , n40256 , n40257 , n40258 , n40259 , n40260 , n40261 , n40262 ,
     n40263 , n40264 , n40265 , n40266 , n40267 , n40268 , n40269 , n40270 , n40271 , n40272 ,
     n40273 , n40274 , n40275 , n40276 , n40277 , n40278 , n40279 , n40280 , n40281 , n40282 ,
     n40283 , n40284 , n40285 , n40286 , n40287 , n40288 , n40289 , n40290 , n40291 , n40292 ,
     n40293 , n40294 , n40295 , n40296 , n40297 , n40298 , n40299 , n40300 , n40301 , n40302 ,
     n40303 , n40304 , n40305 , n40306 , n40307 , n40308 , n40309 , n40310 , n40311 , n40312 ,
     n40313 , n40314 , n40315 , n40316 , n40317 , n40318 , n40319 , n40320 , n40321 , n40322 ,
     n40323 , n40324 , n40325 , n40326 , n40327 , n40328 , n40329 , n40330 , n40331 , n40332 ,
     n40333 , n40334 , n40335 , n40336 , n40337 , n40338 , n40339 , n40340 , n40341 , n40342 ,
     n40343 , n40344 , n40345 , n40346 , n40347 , n40348 , n40349 , n40350 , n40351 , n40352 ,
     n40353 , n40354 , n40355 , n40356 , n40357 , n40358 , n40359 , n40360 , n40361 , n40362 ,
     n40363 , n40364 , n40365 , n40366 , n40367 , n40368 , n40369 , n40370 , n40371 , n40372 ,
     n40373 , n40374 , n40375 , n40376 , n40377 , n40378 , n40379 , n40380 , n40381 , n40382 ,
     n40383 , n40384 , n40385 , n40386 , n40387 , n40388 , n40389 , n40390 , n40391 , n40392 ,
     n40393 , n40394 , n40395 , n40396 , n40397 , n40398 , n40399 , n40400 , n40401 , n40402 ,
     n40403 , n40404 , n40405 , n40406 , n40407 , n40408 , n40409 , n40410 , n40411 , n40412 ,
     n40413 , n40414 , n40415 , n40416 , n40417 , n40418 , n40419 , n40420 , n40421 , n40422 ,
     n40423 , n40424 , n40425 , n40426 , n40427 , n40428 , n40429 , n40430 , n40431 , n40432 ,
     n40433 , n40434 , n40435 , n40436 , n40437 , n40438 , n40439 , n40440 , n40441 , n40442 ,
     n40443 , n40444 , n40445 , n40446 , n40447 , n40448 , n40449 , n40450 , n40451 , n40452 ,
     n40453 , n40454 , n40455 , n40456 , n40457 , n40458 , n40459 , n40460 , n40461 , n40462 ,
     n40463 , n40464 , n40465 , n40466 , n40467 , n40468 , n40469 , n40470 , n40471 , n40472 ,
     n40473 , n40474 , n40475 , n40476 , n40477 , n40478 , n40479 , n40480 , n40481 , n40482 ,
     n40483 , n40484 , n40485 , n40486 , n40487 , n40488 , n40489 , n40490 , n40491 , n40492 ,
     n40493 , n40494 , n40495 , n40496 , n40497 , n40498 , n40499 , n40500 , n40501 , n40502 ,
     n40503 , n40504 , n40505 , n40506 , n40507 , n40508 , n40509 , n40510 , n40511 , n40512 ,
     n40513 , n40514 , n40515 , n40516 , n40517 , n40518 , n40519 , n40520 , n40521 , n40522 ,
     n40523 , n40524 , n40525 , n40526 , n40527 , n40528 , n40529 , n40530 , n40531 , n40532 ,
     n40533 , n40534 , n40535 , n40536 , n40537 , n40538 , n40539 , n40540 , n40541 , n40542 ,
     n40543 , n40544 , n40545 , n40546 , n40547 , n40548 , n40549 , n40550 , n40551 , n40552 ,
     n40553 , n40554 , n40555 , n40556 , n40557 , n40558 , n40559 , n40560 , n40561 , n40562 ,
     n40563 , n40564 , n40565 , n40566 , n40567 , n40568 , n40569 , n40570 , n40571 , n40572 ,
     n40573 , n40574 , n40575 , n40576 , n40577 , n40578 , n40579 , n40580 , n40581 , n40582 ,
     n40583 , n40584 , n40585 , n40586 , n40587 , n40588 , n40589 , n40590 , n40591 , n40592 ,
     n40593 , n40594 , n40595 , n40596 , n40597 , n40598 , n40599 , n40600 , n40601 , n40602 ,
     n40603 , n40604 , n40605 , n40606 , n40607 , n40608 , n40609 , n40610 , n40611 , n40612 ,
     n40613 , n40614 , n40615 , n40616 , n40617 , n40618 , n40619 , n40620 , n40621 , n40622 ,
     n40623 , n40624 , n40625 , n40626 , n40627 , n40628 , n40629 , n40630 , n40631 , n40632 ,
     n40633 , n40634 , n40635 , n40636 , n40637 , n40638 , n40639 , n40640 , n40641 , n40642 ,
     n40643 , n40644 , n40645 , n40646 , n40647 , n40648 , n40649 , n40650 , n40651 , n40652 ,
     n40653 , n40654 , n40655 , n40656 , n40657 , n40658 , n40659 , n40660 , n40661 , n40662 ,
     n40663 , n40664 , n40665 , n40666 , n40667 , n40668 , n40669 , n40670 , n40671 , n40672 ,
     n40673 , n40674 , n40675 , n40676 , n40677 , n40678 , n40679 , n40680 , n40681 , n40682 ,
     n40683 , n40684 , n40685 , n40686 , n40687 , n40688 , n40689 , n40690 , n40691 , n40692 ,
     n40693 , n40694 , n40695 , n40696 , n40697 , n40698 , n40699 , n40700 , n40701 , n40702 ,
     n40703 , n40704 , n40705 , n40706 , n40707 , n40708 , n40709 , n40710 , n40711 , n40712 ,
     n40713 , n40714 , n40715 , n40716 , n40717 , n40718 , n40719 , n40720 , n40721 , n40722 ,
     n40723 , n40724 , n40725 , n40726 , n40727 , n40728 , n40729 , n40730 , n40731 , n40732 ,
     n40733 , n40734 , n40735 , n40736 , n40737 , n40738 , n40739 , n40740 , n40741 , n40742 ,
     n40743 , n40744 , n40745 , n40746 , n40747 , n40748 , n40749 , n40750 , n40751 , n40752 ,
     n40753 , n40754 , n40755 , n40756 , n40757 , n40758 , n40759 , n40760 , n40761 , n40762 ,
     n40763 , n40764 , n40765 , n40766 , n40767 , n40768 , n40769 , n40770 , n40771 , n40772 ,
     n40773 , n40774 , n40775 , n40776 , n40777 , n40778 , n40779 , n40780 , n40781 , n40782 ,
     n40783 , n40784 , n40785 , n40786 , n40787 , n40788 , n40789 , n40790 , n40791 , n40792 ,
     n40793 , n40794 , n40795 , n40796 , n40797 , n40798 , n40799 , n40800 , n40801 , n40802 ,
     n40803 , n40804 , n40805 , n40806 , n40807 , n40808 , n40809 , n40810 , n40811 , n40812 ,
     n40813 , n40814 , n40815 , n40816 , n40817 , n40818 , n40819 , n40820 , n40821 , n40822 ,
     n40823 , n40824 , n40825 , n40826 , n40827 , n40828 , n40829 , n40830 , n40831 , n40832 ,
     n40833 , n40834 , n40835 , n40836 , n40837 , n40838 , n40839 , n40840 , n40841 , n40842 ,
     n40843 , n40844 , n40845 , n40846 , n40847 , n40848 , n40849 , n40850 , n40851 , n40852 ,
     n40853 , n40854 , n40855 , n40856 , n40857 , n40858 , n40859 , n40860 , n40861 , n40862 ,
     n40863 , n40864 , n40865 , n40866 , n40867 , n40868 , n40869 , n40870 , n40871 , n40872 ,
     n40873 , n40874 , n40875 , n40876 , n40877 , n40878 , n40879 , n40880 , n40881 , n40882 ,
     n40883 , n40884 , n40885 , n40886 , n40887 , n40888 , n40889 , n40890 , n40891 , n40892 ,
     n40893 , n40894 , n40895 , n40896 , n40897 , n40898 , n40899 , n40900 , n40901 , n40902 ,
     n40903 , n40904 , n40905 , n40906 , n40907 , n40908 , n40909 , n40910 , n40911 , n40912 ,
     n40913 , n40914 , n40915 , n40916 , n40917 , n40918 , n40919 , n40920 , n40921 , n40922 ,
     n40923 , n40924 , n40925 , n40926 , n40927 , n40928 , n40929 , n40930 , n40931 , n40932 ,
     n40933 , n40934 , n40935 , n40936 , n40937 , n40938 , n40939 , n40940 , n40941 , n40942 ,
     n40943 , n40944 , n40945 , n40946 , n40947 , n40948 , n40949 , n40950 , n40951 , n40952 ,
     n40953 , n40954 , n40955 , n40956 , n40957 , n40958 , n40959 , n40960 , n40961 , n40962 ,
     n40963 , n40964 , n40965 , n40966 , n40967 , n40968 , n40969 , n40970 , n40971 , n40972 ,
     n40973 , n40974 , n40975 , n40976 , n40977 , n40978 , n40979 , n40980 , n40981 , n40982 ,
     n40983 , n40984 , n40985 , n40986 , n40987 , n40988 , n40989 , n40990 , n40991 , n40992 ,
     n40993 , n40994 , n40995 , n40996 , n40997 , n40998 , n40999 , n41000 , n41001 , n41002 ,
     n41003 , n41004 , n41005 , n41006 , n41007 , n41008 , n41009 , n41010 , n41011 , n41012 ,
     n41013 , n41014 , n41015 , n41016 , n41017 , n41018 , n41019 , n41020 , n41021 , n41022 ,
     n41023 , n41024 , n41025 , n41026 , n41027 , n41028 , n41029 , n41030 , n41031 , n41032 ,
     n41033 , n41034 , n41035 , n41036 , n41037 , n41038 , n41039 , n41040 , n41041 , n41042 ,
     n41043 , n41044 , n41045 , n41046 , n41047 , n41048 , n41049 , n41050 , n41051 , n41052 ,
     n41053 , n41054 , n41055 , n41056 , n41057 , n41058 , n41059 , n41060 , n41061 , n41062 ,
     n41063 , n41064 , n41065 , n41066 , n41067 , n41068 , n41069 , n41070 , n41071 , n41072 ,
     n41073 , n41074 , n41075 , n41076 , n41077 , n41078 , n41079 , n41080 , n41081 , n41082 ,
     n41083 , n41084 , n41085 , n41086 , n41087 , n41088 , n41089 , n41090 , n41091 , n41092 ,
     n41093 , n41094 , n41095 , n41096 , n41097 , n41098 , n41099 , n41100 , n41101 , n41102 ,
     n41103 , n41104 , n41105 , n41106 , n41107 , n41108 , n41109 , n41110 , n41111 , n41112 ,
     n41113 , n41114 , n41115 , n41116 , n41117 , n41118 , n41119 , n41120 , n41121 , n41122 ,
     n41123 , n41124 , n41125 , n41126 , n41127 , n41128 , n41129 , n41130 , n41131 , n41132 ,
     n41133 , n41134 , n41135 , n41136 , n41137 , n41138 , n41139 , n41140 , n41141 , n41142 ,
     n41143 , n41144 , n41145 , n41146 , n41147 , n41148 , n41149 , n41150 , n41151 , n41152 ,
     n41153 , n41154 , n41155 , n41156 , n41157 , n41158 , n41159 , n41160 , n41161 , n41162 ,
     n41163 , n41164 , n41165 , n41166 , n41167 , n41168 , n41169 , n41170 , n41171 , n41172 ,
     n41173 , n41174 , n41175 , n41176 , n41177 , n41178 , n41179 , n41180 , n41181 , n41182 ,
     n41183 , n41184 , n41185 , n41186 , n41187 , n41188 , n41189 , n41190 , n41191 , n41192 ,
     n41193 , n41194 , n41195 , n41196 , n41197 , n41198 , n41199 , n41200 , n41201 , n41202 ,
     n41203 , n41204 , n41205 , n41206 , n41207 , n41208 , n41209 , n41210 , n41211 , n41212 ,
     n41213 , n41214 , n41215 , n41216 , n41217 , n41218 , n41219 , n41220 , n41221 , n41222 ,
     n41223 , n41224 , n41225 , n41226 , n41227 , n41228 , n41229 , n41230 , n41231 , n41232 ,
     n41233 , n41234 , n41235 , n41236 , n41237 , n41238 , n41239 , n41240 , n41241 , n41242 ,
     n41243 , n41244 , n41245 , n41246 , n41247 , n41248 , n41249 , n41250 , n41251 , n41252 ,
     n41253 , n41254 , n41255 , n41256 , n41257 , n41258 , n41259 , n41260 , n41261 , n41262 ,
     n41263 , n41264 , n41265 , n41266 , n41267 , n41268 , n41269 , n41270 , n41271 , n41272 ,
     n41273 , n41274 , n41275 , n41276 , n41277 , n41278 , n41279 , n41280 , n41281 , n41282 ,
     n41283 , n41284 , n41285 , n41286 , n41287 , n41288 , n41289 , n41290 , n41291 , n41292 ,
     n41293 , n41294 , n41295 , n41296 , n41297 , n41298 , n41299 , n41300 , n41301 , n41302 ,
     n41303 , n41304 , n41305 , n41306 , n41307 , n41308 , n41309 , n41310 , n41311 , n41312 ,
     n41313 , n41314 , n41315 , n41316 , n41317 , n41318 , n41319 , n41320 , n41321 , n41322 ,
     n41323 , n41324 , n41325 , n41326 , n41327 , n41328 , n41329 , n41330 , n41331 , n41332 ,
     n41333 , n41334 , n41335 , n41336 , n41337 , n41338 , n41339 , n41340 , n41341 , n41342 ,
     n41343 , n41344 , n41345 , n41346 , n41347 , n41348 , n41349 , n41350 , n41351 , n41352 ,
     n41353 , n41354 , n41355 , n41356 , n41357 , n41358 , n41359 , n41360 , n41361 , n41362 ,
     n41363 , n41364 , n41365 , n41366 , n41367 , n41368 , n41369 , n41370 , n41371 , n41372 ,
     n41373 , n41374 , n41375 , n41376 , n41377 , n41378 , n41379 , n41380 , n41381 , n41382 ,
     n41383 , n41384 , n41385 , n41386 , n41387 , n41388 , n41389 , n41390 , n41391 , n41392 ,
     n41393 , n41394 , n41395 , n41396 , n41397 , n41398 , n41399 , n41400 , n41401 , n41402 ,
     n41403 , n41404 , n41405 , n41406 , n41407 , n41408 , n41409 , n41410 , n41411 , n41412 ,
     n41413 , n41414 , n41415 , n41416 , n41417 , n41418 , n41419 , n41420 , n41421 , n41422 ,
     n41423 , n41424 , n41425 , n41426 , n41427 , n41428 , n41429 , n41430 , n41431 , n41432 ,
     n41433 , n41434 , n41435 , n41436 , n41437 , n41438 , n41439 , n41440 , n41441 , n41442 ,
     n41443 , n41444 , n41445 , n41446 , n41447 , n41448 , n41449 , n41450 , n41451 , n41452 ,
     n41453 , n41454 , n41455 , n41456 , n41457 , n41458 , n41459 , n41460 , n41461 , n41462 ,
     n41463 , n41464 , n41465 , n41466 , n41467 , n41468 , n41469 , n41470 , n41471 , n41472 ,
     n41473 , n41474 , n41475 , n41476 , n41477 , n41478 , n41479 , n41480 , n41481 , n41482 ,
     n41483 , n41484 , n41485 , n41486 , n41487 , n41488 , n41489 , n41490 , n41491 , n41492 ,
     n41493 , n41494 , n41495 , n41496 , n41497 , n41498 , n41499 , n41500 , n41501 , n41502 ,
     n41503 , n41504 , n41505 , n41506 , n41507 , n41508 , n41509 , n41510 , n41511 , n41512 ,
     n41513 , n41514 , n41515 , n41516 , n41517 , n41518 , n41519 , n41520 , n41521 , n41522 ,
     n41523 , n41524 , n41525 , n41526 , n41527 , n41528 , n41529 , n41530 , n41531 , n41532 ,
     n41533 , n41534 , n41535 , n41536 , n41537 , n41538 , n41539 , n41540 , n41541 , n41542 ,
     n41543 , n41544 , n41545 , n41546 , n41547 , n41548 , n41549 , n41550 , n41551 , n41552 ,
     n41553 , n41554 , n41555 , n41556 , n41557 , n41558 , n41559 , n41560 , n41561 , n41562 ,
     n41563 , n41564 , n41565 , n41566 , n41567 , n41568 , n41569 , n41570 , n41571 , n41572 ,
     n41573 , n41574 , n41575 , n41576 , n41577 , n41578 , n41579 , n41580 , n41581 , n41582 ,
     n41583 , n41584 , n41585 , n41586 , n41587 , n41588 , n41589 , n41590 , n41591 , n41592 ,
     n41593 , n41594 , n41595 , n41596 , n41597 , n41598 , n41599 , n41600 , n41601 , n41602 ,
     n41603 , n41604 , n41605 , n41606 , n41607 , n41608 , n41609 , n41610 , n41611 , n41612 ,
     n41613 , n41614 , n41615 , n41616 , n41617 , n41618 , n41619 , n41620 , n41621 , n41622 ,
     n41623 , n41624 , n41625 , n41626 , n41627 , n41628 , n41629 , n41630 , n41631 , n41632 ,
     n41633 , n41634 , n41635 , n41636 , n41637 , n41638 , n41639 , n41640 , n41641 , n41642 ,
     n41643 , n41644 , n41645 , n41646 , n41647 , n41648 , n41649 , n41650 , n41651 , n41652 ,
     n41653 , n41654 , n41655 , n41656 , n41657 , n41658 , n41659 , n41660 , n41661 , n41662 ,
     n41663 , n41664 , n41665 , n41666 , n41667 , n41668 , n41669 , n41670 , n41671 , n41672 ,
     n41673 , n41674 , n41675 , n41676 , n41677 , n41678 , n41679 , n41680 , n41681 , n41682 ,
     n41683 , n41684 , n41685 , n41686 , n41687 , n41688 , n41689 , n41690 , n41691 , n41692 ,
     n41693 , n41694 , n41695 , n41696 , n41697 , n41698 , n41699 , n41700 , n41701 , n41702 ,
     n41703 , n41704 , n41705 , n41706 , n41707 , n41708 , n41709 , n41710 , n41711 , n41712 ,
     n41713 , n41714 , n41715 , n41716 , n41717 , n41718 , n41719 , n41720 , n41721 , n41722 ,
     n41723 , n41724 , n41725 , n41726 , n41727 , n41728 , n41729 , n41730 , n41731 , n41732 ,
     n41733 , n41734 , n41735 , n41736 , n41737 , n41738 , n41739 , n41740 , n41741 , n41742 ,
     n41743 , n41744 , n41745 , n41746 , n41747 , n41748 , n41749 , n41750 , n41751 , n41752 ,
     n41753 , n41754 , n41755 , n41756 , n41757 , n41758 , n41759 , n41760 , n41761 , n41762 ,
     n41763 , n41764 , n41765 , n41766 , n41767 , n41768 , n41769 , n41770 , n41771 , n41772 ,
     n41773 , n41774 , n41775 , n41776 , n41777 , n41778 , n41779 , n41780 , n41781 , n41782 ,
     n41783 , n41784 , n41785 , n41786 , n41787 , n41788 , n41789 , n41790 , n41791 , n41792 ,
     n41793 , n41794 , n41795 , n41796 , n41797 , n41798 , n41799 , n41800 , n41801 , n41802 ,
     n41803 , n41804 , n41805 , n41806 , n41807 , n41808 , n41809 , n41810 , n41811 , n41812 ,
     n41813 , n41814 , n41815 , n41816 , n41817 , n41818 , n41819 , n41820 , n41821 , n41822 ,
     n41823 , n41824 , n41825 , n41826 , n41827 , n41828 , n41829 , n41830 , n41831 , n41832 ,
     n41833 , n41834 , n41835 , n41836 , n41837 , n41838 , n41839 , n41840 , n41841 , n41842 ,
     n41843 , n41844 , n41845 , n41846 , n41847 , n41848 , n41849 , n41850 , n41851 , n41852 ,
     n41853 , n41854 , n41855 , n41856 , n41857 , n41858 , n41859 , n41860 , n41861 , n41862 ,
     n41863 , n41864 , n41865 , n41866 , n41867 , n41868 , n41869 , n41870 , n41871 , n41872 ,
     n41873 , n41874 , n41875 , n41876 , n41877 , n41878 , n41879 , n41880 , n41881 , n41882 ,
     n41883 , n41884 , n41885 , n41886 , n41887 , n41888 , n41889 , n41890 , n41891 , n41892 ,
     n41893 , n41894 , n41895 , n41896 , n41897 , n41898 , n41899 , n41900 , n41901 , n41902 ,
     n41903 , n41904 , n41905 , n41906 , n41907 , n41908 , n41909 , n41910 , n41911 , n41912 ,
     n41913 , n41914 , n41915 , n41916 , n41917 , n41918 , n41919 , n41920 , n41921 , n41922 ,
     n41923 , n41924 , n41925 , n41926 , n41927 , n41928 , n41929 , n41930 , n41931 , n41932 ,
     n41933 , n41934 , n41935 , n41936 , n41937 , n41938 , n41939 , n41940 , n41941 , n41942 ,
     n41943 , n41944 , n41945 , n41946 , n41947 , n41948 , n41949 , n41950 , n41951 , n41952 ,
     n41953 , n41954 , n41955 , n41956 , n41957 , n41958 , n41959 , n41960 , n41961 , n41962 ,
     n41963 , n41964 , n41965 , n41966 , n41967 , n41968 , n41969 , n41970 , n41971 , n41972 ,
     n41973 , n41974 , n41975 , n41976 , n41977 , n41978 , n41979 , n41980 , n41981 , n41982 ,
     n41983 , n41984 , n41985 , n41986 , n41987 , n41988 , n41989 , n41990 , n41991 , n41992 ,
     n41993 , n41994 , n41995 , n41996 , n41997 , n41998 , n41999 , n42000 , n42001 , n42002 ,
     n42003 , n42004 , n42005 , n42006 , n42007 , n42008 , n42009 , n42010 , n42011 , n42012 ,
     n42013 , n42014 , n42015 , n42016 , n42017 , n42018 , n42019 , n42020 , n42021 , n42022 ,
     n42023 , n42024 , n42025 , n42026 , n42027 , n42028 , n42029 , n42030 , n42031 , n42032 ,
     n42033 , n42034 , n42035 , n42036 , n42037 , n42038 , n42039 , n42040 , n42041 , n42042 ,
     n42043 , n42044 , n42045 , n42046 , n42047 , n42048 , n42049 , n42050 , n42051 , n42052 ,
     n42053 , n42054 , n42055 , n42056 , n42057 , n42058 , n42059 , n42060 , n42061 , n42062 ,
     n42063 , n42064 , n42065 , n42066 , n42067 , n42068 , n42069 , n42070 , n42071 , n42072 ,
     n42073 , n42074 , n42075 , n42076 , n42077 , n42078 , n42079 , n42080 , n42081 , n42082 ,
     n42083 , n42084 , n42085 , n42086 , n42087 , n42088 , n42089 , n42090 , n42091 , n42092 ,
     n42093 , n42094 , n42095 , n42096 , n42097 , n42098 , n42099 , n42100 , n42101 , n42102 ,
     n42103 , n42104 , n42105 , n42106 , n42107 , n42108 , n42109 , n42110 , n42111 , n42112 ,
     n42113 , n42114 , n42115 , n42116 , n42117 , n42118 , n42119 , n42120 , n42121 , n42122 ,
     n42123 , n42124 , n42125 , n42126 , n42127 , n42128 , n42129 , n42130 , n42131 , n42132 ,
     n42133 , n42134 , n42135 , n42136 , n42137 , n42138 , n42139 , n42140 , n42141 , n42142 ,
     n42143 , n42144 , n42145 , n42146 , n42147 , n42148 , n42149 , n42150 , n42151 , n42152 ,
     n42153 , n42154 , n42155 , n42156 , n42157 , n42158 , n42159 , n42160 , n42161 , n42162 ,
     n42163 , n42164 , n42165 , n42166 , n42167 , n42168 , n42169 , n42170 , n42171 , n42172 ,
     n42173 , n42174 , n42175 , n42176 , n42177 , n42178 , n42179 , n42180 , n42181 , n42182 ,
     n42183 , n42184 , n42185 , n42186 , n42187 , n42188 , n42189 , n42190 , n42191 , n42192 ,
     n42193 , n42194 , n42195 , n42196 , n42197 , n42198 , n42199 , n42200 , n42201 , n42202 ,
     n42203 , n42204 , n42205 , n42206 , n42207 , n42208 , n42209 , n42210 , n42211 , n42212 ,
     n42213 , n42214 , n42215 , n42216 , n42217 , n42218 , n42219 , n42220 , n42221 , n42222 ,
     n42223 , n42224 , n42225 , n42226 , n42227 , n42228 , n42229 , n42230 , n42231 , n42232 ,
     n42233 , n42234 , n42235 , n42236 , n42237 , n42238 , n42239 , n42240 , n42241 , n42242 ,
     n42243 , n42244 , n42245 , n42246 , n42247 , n42248 , n42249 , n42250 , n42251 , n42252 ,
     n42253 , n42254 , n42255 , n42256 , n42257 , n42258 , n42259 , n42260 , n42261 , n42262 ,
     n42263 , n42264 , n42265 , n42266 , n42267 , n42268 , n42269 , n42270 , n42271 , n42272 ,
     n42273 , n42274 , n42275 , n42276 , n42277 , n42278 , n42279 , n42280 , n42281 , n42282 ,
     n42283 , n42284 , n42285 , n42286 , n42287 , n42288 , n42289 , n42290 , n42291 , n42292 ,
     n42293 , n42294 , n42295 , n42296 , n42297 , n42298 , n42299 , n42300 , n42301 , n42302 ,
     n42303 , n42304 , n42305 , n42306 , n42307 , n42308 , n42309 , n42310 , n42311 , n42312 ,
     n42313 , n42314 , n42315 , n42316 , n42317 , n42318 , n42319 , n42320 , n42321 , n42322 ,
     n42323 , n42324 , n42325 , n42326 , n42327 , n42328 , n42329 , n42330 , n42331 , n42332 ,
     n42333 , n42334 , n42335 , n42336 , n42337 , n42338 , n42339 , n42340 , n42341 , n42342 ,
     n42343 , n42344 , n42345 , n42346 , n42347 , n42348 , n42349 , n42350 , n42351 , n42352 ,
     n42353 , n42354 , n42355 , n42356 , n42357 , n42358 , n42359 , n42360 , n42361 , n42362 ,
     n42363 , n42364 , n42365 , n42366 , n42367 , n42368 , n42369 , n42370 , n42371 , n42372 ,
     n42373 , n42374 , n42375 , n42376 , n42377 , n42378 , n42379 , n42380 , n42381 , n42382 ,
     n42383 , n42384 , n42385 , n42386 , n42387 , n42388 , n42389 , n42390 , n42391 , n42392 ,
     n42393 , n42394 , n42395 , n42396 , n42397 , n42398 , n42399 , n42400 , n42401 , n42402 ,
     n42403 , n42404 , n42405 , n42406 , n42407 , n42408 , n42409 , n42410 , n42411 , n42412 ,
     n42413 , n42414 , n42415 , n42416 , n42417 , n42418 , n42419 , n42420 , n42421 , n42422 ,
     n42423 , n42424 , n42425 , n42426 , n42427 , n42428 , n42429 , n42430 , n42431 , n42432 ,
     n42433 , n42434 , n42435 , n42436 , n42437 , n42438 , n42439 , n42440 , n42441 , n42442 ,
     n42443 , n42444 , n42445 , n42446 , n42447 , n42448 , n42449 , n42450 , n42451 , n42452 ,
     n42453 , n42454 , n42455 , n42456 , n42457 , n42458 , n42459 , n42460 , n42461 , n42462 ,
     n42463 , n42464 , n42465 , n42466 , n42467 , n42468 , n42469 , n42470 , n42471 , n42472 ,
     n42473 , n42474 , n42475 , n42476 , n42477 , n42478 , n42479 , n42480 , n42481 , n42482 ,
     n42483 , n42484 , n42485 , n42486 , n42487 , n42488 , n42489 , n42490 , n42491 , n42492 ,
     n42493 , n42494 , n42495 , n42496 , n42497 , n42498 , n42499 , n42500 , n42501 , n42502 ,
     n42503 , n42504 , n42505 , n42506 , n42507 , n42508 , n42509 , n42510 , n42511 , n42512 ,
     n42513 , n42514 , n42515 , n42516 , n42517 , n42518 , n42519 , n42520 , n42521 , n42522 ,
     n42523 , n42524 , n42525 , n42526 , n42527 , n42528 , n42529 , n42530 , n42531 , n42532 ,
     n42533 , n42534 , n42535 , n42536 , n42537 , n42538 , n42539 , n42540 , n42541 , n42542 ,
     n42543 , n42544 , n42545 , n42546 , n42547 , n42548 , n42549 , n42550 , n42551 , n42552 ,
     n42553 , n42554 , n42555 , n42556 , n42557 , n42558 , n42559 , n42560 , n42561 , n42562 ,
     n42563 , n42564 , n42565 , n42566 , n42567 , n42568 , n42569 , n42570 , n42571 , n42572 ,
     n42573 , n42574 , n42575 , n42576 , n42577 , n42578 , n42579 , n42580 , n42581 , n42582 ,
     n42583 , n42584 , n42585 , n42586 , n42587 , n42588 , n42589 , n42590 , n42591 , n42592 ,
     n42593 , n42594 , n42595 , n42596 , n42597 , n42598 , n42599 , n42600 , n42601 , n42602 ,
     n42603 , n42604 , n42605 , n42606 , n42607 , n42608 , n42609 , n42610 , n42611 , n42612 ,
     n42613 , n42614 , n42615 , n42616 , n42617 , n42618 , n42619 , n42620 , n42621 , n42622 ,
     n42623 , n42624 , n42625 , n42626 , n42627 , n42628 , n42629 , n42630 , n42631 , n42632 ,
     n42633 , n42634 , n42635 , n42636 , n42637 , n42638 , n42639 , n42640 , n42641 , n42642 ,
     n42643 , n42644 , n42645 , n42646 , n42647 , n42648 , n42649 , n42650 , n42651 , n42652 ,
     n42653 , n42654 , n42655 , n42656 , n42657 , n42658 , n42659 , n42660 , n42661 , n42662 ,
     n42663 , n42664 , n42665 , n42666 , n42667 , n42668 , n42669 , n42670 , n42671 , n42672 ,
     n42673 , n42674 , n42675 , n42676 , n42677 , n42678 , n42679 , n42680 , n42681 , n42682 ,
     n42683 , n42684 , n42685 , n42686 , n42687 , n42688 , n42689 , n42690 , n42691 , n42692 ,
     n42693 , n42694 , n42695 , n42696 , n42697 , n42698 , n42699 , n42700 , n42701 , n42702 ,
     n42703 , n42704 , n42705 , n42706 , n42707 , n42708 , n42709 , n42710 , n42711 , n42712 ,
     n42713 , n42714 , n42715 , n42716 , n42717 , n42718 , n42719 , n42720 , n42721 , n42722 ,
     n42723 , n42724 , n42725 , n42726 , n42727 , n42728 , n42729 , n42730 , n42731 , n42732 ,
     n42733 , n42734 , n42735 , n42736 , n42737 , n42738 , n42739 , n42740 , n42741 , n42742 ,
     n42743 , n42744 , n42745 , n42746 , n42747 , n42748 , n42749 , n42750 , n42751 , n42752 ,
     n42753 , n42754 , n42755 , n42756 , n42757 , n42758 , n42759 , n42760 , n42761 , n42762 ,
     n42763 , n42764 , n42765 , n42766 , n42767 , n42768 , n42769 , n42770 , n42771 , n42772 ,
     n42773 , n42774 , n42775 , n42776 , n42777 , n42778 , n42779 , n42780 , n42781 , n42782 ,
     n42783 , n42784 , n42785 , n42786 , n42787 , n42788 , n42789 , n42790 , n42791 , n42792 ,
     n42793 , n42794 , n42795 , n42796 , n42797 , n42798 , n42799 , n42800 , n42801 , n42802 ,
     n42803 , n42804 , n42805 , n42806 , n42807 , n42808 , n42809 , n42810 , n42811 , n42812 ,
     n42813 , n42814 , n42815 , n42816 , n42817 , n42818 , n42819 , n42820 , n42821 , n42822 ,
     n42823 , n42824 , n42825 , n42826 , n42827 , n42828 , n42829 , n42830 , n42831 , n42832 ,
     n42833 , n42834 , n42835 , n42836 , n42837 , n42838 , n42839 , n42840 , n42841 , n42842 ,
     n42843 , n42844 , n42845 , n42846 , n42847 , n42848 , n42849 , n42850 , n42851 , n42852 ,
     n42853 , n42854 , n42855 , n42856 , n42857 , n42858 , n42859 , n42860 , n42861 , n42862 ,
     n42863 , n42864 , n42865 , n42866 , n42867 , n42868 , n42869 , n42870 , n42871 , n42872 ,
     n42873 , n42874 , n42875 , n42876 , n42877 , n42878 , n42879 , n42880 , n42881 , n42882 ,
     n42883 , n42884 , n42885 , n42886 , n42887 , n42888 , n42889 , n42890 , n42891 , n42892 ,
     n42893 , n42894 , n42895 , n42896 , n42897 , n42898 , n42899 , n42900 , n42901 , n42902 ,
     n42903 , n42904 , n42905 , n42906 , n42907 , n42908 , n42909 , n42910 , n42911 , n42912 ,
     n42913 , n42914 , n42915 , n42916 , n42917 , n42918 , n42919 , n42920 , n42921 , n42922 ,
     n42923 , n42924 , n42925 , n42926 , n42927 , n42928 , n42929 , n42930 , n42931 , n42932 ,
     n42933 , n42934 , n42935 , n42936 , n42937 , n42938 , n42939 , n42940 , n42941 , n42942 ,
     n42943 , n42944 , n42945 , n42946 , n42947 , n42948 , n42949 , n42950 , n42951 , n42952 ,
     n42953 , n42954 , n42955 , n42956 , n42957 , n42958 , n42959 , n42960 , n42961 , n42962 ,
     n42963 , n42964 , n42965 , n42966 , n42967 , n42968 , n42969 , n42970 , n42971 , n42972 ,
     n42973 , n42974 , n42975 , n42976 , n42977 , n42978 , n42979 , n42980 , n42981 , n42982 ,
     n42983 , n42984 , n42985 , n42986 , n42987 , n42988 , n42989 , n42990 , n42991 , n42992 ,
     n42993 , n42994 , n42995 , n42996 , n42997 , n42998 , n42999 , n43000 , n43001 , n43002 ,
     n43003 , n43004 , n43005 , n43006 , n43007 , n43008 , n43009 , n43010 , n43011 , n43012 ,
     n43013 , n43014 , n43015 , n43016 , n43017 , n43018 , n43019 , n43020 , n43021 , n43022 ,
     n43023 , n43024 , n43025 , n43026 , n43027 , n43028 , n43029 , n43030 , n43031 , n43032 ,
     n43033 , n43034 , n43035 , n43036 , n43037 , n43038 , n43039 , n43040 , n43041 , n43042 ,
     n43043 , n43044 , n43045 , n43046 , n43047 , n43048 , n43049 , n43050 , n43051 , n43052 ,
     n43053 , n43054 , n43055 , n43056 , n43057 , n43058 , n43059 , n43060 , n43061 , n43062 ,
     n43063 , n43064 , n43065 , n43066 , n43067 , n43068 , n43069 , n43070 , n43071 , n43072 ,
     n43073 , n43074 , n43075 , n43076 , n43077 , n43078 , n43079 , n43080 , n43081 , n43082 ,
     n43083 , n43084 , n43085 , n43086 , n43087 , n43088 , n43089 , n43090 , n43091 , n43092 ,
     n43093 , n43094 , n43095 , n43096 , n43097 , n43098 , n43099 , n43100 , n43101 , n43102 ,
     n43103 , n43104 , n43105 , n43106 , n43107 , n43108 , n43109 , n43110 , n43111 , n43112 ,
     n43113 , n43114 , n43115 , n43116 , n43117 , n43118 , n43119 , n43120 , n43121 , n43122 ,
     n43123 , n43124 , n43125 , n43126 , n43127 , n43128 , n43129 , n43130 , n43131 , n43132 ,
     n43133 , n43134 , n43135 , n43136 , n43137 , n43138 , n43139 , n43140 , n43141 , n43142 ,
     n43143 , n43144 , n43145 , n43146 , n43147 , n43148 , n43149 , n43150 , n43151 , n43152 ,
     n43153 , n43154 , n43155 , n43156 , n43157 , n43158 , n43159 , n43160 , n43161 , n43162 ,
     n43163 , n43164 , n43165 , n43166 , n43167 , n43168 , n43169 , n43170 , n43171 , n43172 ,
     n43173 , n43174 , n43175 , n43176 , n43177 , n43178 , n43179 , n43180 , n43181 , n43182 ,
     n43183 , n43184 , n43185 , n43186 , n43187 , n43188 , n43189 , n43190 , n43191 , n43192 ,
     n43193 , n43194 , n43195 , n43196 , n43197 , n43198 , n43199 , n43200 , n43201 , n43202 ,
     n43203 , n43204 , n43205 , n43206 , n43207 , n43208 , n43209 , n43210 , n43211 , n43212 ,
     n43213 , n43214 , n43215 , n43216 , n43217 , n43218 , n43219 , n43220 , n43221 , n43222 ,
     n43223 , n43224 , n43225 , n43226 , n43227 , n43228 , n43229 , n43230 , n43231 , n43232 ,
     n43233 , n43234 , n43235 , n43236 , n43237 , n43238 , n43239 , n43240 , n43241 , n43242 ,
     n43243 , n43244 , n43245 , n43246 , n43247 , n43248 , n43249 , n43250 , n43251 , n43252 ,
     n43253 , n43254 , n43255 , n43256 , n43257 , n43258 , n43259 , n43260 , n43261 , n43262 ,
     n43263 , n43264 , n43265 , n43266 , n43267 , n43268 , n43269 , n43270 , n43271 , n43272 ,
     n43273 , n43274 , n43275 , n43276 , n43277 , n43278 , n43279 , n43280 , n43281 , n43282 ,
     n43283 , n43284 , n43285 , n43286 , n43287 , n43288 , n43289 , n43290 , n43291 , n43292 ,
     n43293 , n43294 , n43295 , n43296 , n43297 , n43298 , n43299 , n43300 , n43301 , n43302 ,
     n43303 , n43304 , n43305 , n43306 , n43307 , n43308 , n43309 , n43310 , n43311 , n43312 ,
     n43313 , n43314 , n43315 , n43316 , n43317 , n43318 , n43319 , n43320 , n43321 , n43322 ,
     n43323 , n43324 , n43325 , n43326 , n43327 , n43328 , n43329 , n43330 , n43331 , n43332 ,
     n43333 , n43334 , n43335 , n43336 , n43337 , n43338 , n43339 , n43340 , n43341 , n43342 ,
     n43343 , n43344 , n43345 , n43346 , n43347 , n43348 , n43349 , n43350 , n43351 , n43352 ,
     n43353 , n43354 , n43355 , n43356 , n43357 , n43358 , n43359 , n43360 , n43361 , n43362 ,
     n43363 , n43364 , n43365 , n43366 , n43367 , n43368 , n43369 , n43370 , n43371 , n43372 ,
     n43373 , n43374 , n43375 , n43376 , n43377 , n43378 , n43379 , n43380 , n43381 , n43382 ,
     n43383 , n43384 , n43385 , n43386 , n43387 , n43388 , n43389 , n43390 , n43391 , n43392 ,
     n43393 , n43394 , n43395 , n43396 , n43397 , n43398 , n43399 , n43400 , n43401 , n43402 ,
     n43403 , n43404 , n43405 , n43406 , n43407 , n43408 , n43409 , n43410 , n43411 , n43412 ,
     n43413 , n43414 , n43415 , n43416 , n43417 , n43418 , n43419 , n43420 , n43421 , n43422 ,
     n43423 , n43424 , n43425 , n43426 , n43427 , n43428 , n43429 , n43430 , n43431 , n43432 ,
     n43433 , n43434 , n43435 , n43436 , n43437 , n43438 , n43439 , n43440 , n43441 , n43442 ,
     n43443 , n43444 , n43445 , n43446 , n43447 , n43448 , n43449 , n43450 , n43451 , n43452 ,
     n43453 , n43454 , n43455 , n43456 , n43457 , n43458 , n43459 , n43460 , n43461 , n43462 ,
     n43463 , n43464 , n43465 , n43466 , n43467 , n43468 , n43469 , n43470 , n43471 , n43472 ,
     n43473 , n43474 , n43475 , n43476 , n43477 , n43478 , n43479 , n43480 , n43481 , n43482 ,
     n43483 , n43484 , n43485 , n43486 , n43487 , n43488 , n43489 , n43490 , n43491 , n43492 ,
     n43493 , n43494 , n43495 , n43496 , n43497 , n43498 , n43499 , n43500 , n43501 , n43502 ,
     n43503 , n43504 , n43505 , n43506 , n43507 , n43508 , n43509 , n43510 , n43511 , n43512 ,
     n43513 , n43514 , n43515 , n43516 , n43517 , n43518 , n43519 , n43520 , n43521 , n43522 ,
     n43523 , n43524 , n43525 , n43526 , n43527 , n43528 , n43529 , n43530 , n43531 , n43532 ,
     n43533 , n43534 , n43535 , n43536 , n43537 , n43538 , n43539 , n43540 , n43541 , n43542 ,
     n43543 , n43544 , n43545 , n43546 , n43547 , n43548 , n43549 , n43550 , n43551 , n43552 ,
     n43553 , n43554 , n43555 , n43556 , n43557 , n43558 , n43559 , n43560 , n43561 , n43562 ,
     n43563 , n43564 , n43565 , n43566 , n43567 , n43568 , n43569 , n43570 , n43571 , n43572 ,
     n43573 , n43574 , n43575 , n43576 , n43577 , n43578 , n43579 , n43580 , n43581 , n43582 ,
     n43583 , n43584 , n43585 , n43586 , n43587 , n43588 , n43589 , n43590 , n43591 , n43592 ,
     n43593 , n43594 , n43595 , n43596 , n43597 , n43598 , n43599 , n43600 , n43601 , n43602 ,
     n43603 , n43604 , n43605 , n43606 , n43607 , n43608 , n43609 , n43610 , n43611 , n43612 ,
     n43613 , n43614 , n43615 , n43616 , n43617 , n43618 , n43619 , n43620 , n43621 , n43622 ,
     n43623 , n43624 , n43625 , n43626 , n43627 , n43628 , n43629 , n43630 , n43631 , n43632 ,
     n43633 , n43634 , n43635 , n43636 , n43637 , n43638 , n43639 , n43640 , n43641 , n43642 ,
     n43643 , n43644 , n43645 , n43646 , n43647 , n43648 , n43649 , n43650 , n43651 , n43652 ,
     n43653 , n43654 , n43655 , n43656 , n43657 , n43658 , n43659 , n43660 , n43661 , n43662 ,
     n43663 , n43664 , n43665 , n43666 , n43667 , n43668 , n43669 , n43670 , n43671 , n43672 ,
     n43673 , n43674 , n43675 , n43676 , n43677 , n43678 , n43679 , n43680 , n43681 , n43682 ,
     n43683 , n43684 , n43685 , n43686 , n43687 , n43688 , n43689 , n43690 , n43691 , n43692 ,
     n43693 , n43694 , n43695 , n43696 , n43697 , n43698 , n43699 , n43700 , n43701 , n43702 ,
     n43703 , n43704 , n43705 , n43706 , n43707 , n43708 , n43709 , n43710 , n43711 , n43712 ,
     n43713 , n43714 , n43715 , n43716 , n43717 , n43718 , n43719 , n43720 , n43721 , n43722 ,
     n43723 , n43724 , n43725 , n43726 , n43727 , n43728 , n43729 , n43730 , n43731 , n43732 ,
     n43733 , n43734 , n43735 , n43736 , n43737 , n43738 , n43739 , n43740 , n43741 , n43742 ,
     n43743 , n43744 , n43745 , n43746 , n43747 , n43748 , n43749 , n43750 , n43751 , n43752 ,
     n43753 , n43754 , n43755 , n43756 , n43757 , n43758 , n43759 , n43760 , n43761 , n43762 ,
     n43763 , n43764 , n43765 , n43766 , n43767 , n43768 , n43769 , n43770 , n43771 , n43772 ,
     n43773 , n43774 , n43775 , n43776 , n43777 , n43778 , n43779 , n43780 , n43781 , n43782 ,
     n43783 , n43784 , n43785 , n43786 , n43787 , n43788 , n43789 , n43790 , n43791 , n43792 ,
     n43793 , n43794 , n43795 , n43796 , n43797 , n43798 , n43799 , n43800 , n43801 , n43802 ,
     n43803 , n43804 , n43805 , n43806 , n43807 , n43808 , n43809 , n43810 , n43811 , n43812 ,
     n43813 , n43814 , n43815 , n43816 , n43817 , n43818 , n43819 , n43820 , n43821 , n43822 ,
     n43823 , n43824 , n43825 , n43826 , n43827 , n43828 , n43829 , n43830 , n43831 , n43832 ,
     n43833 , n43834 , n43835 , n43836 , n43837 , n43838 , n43839 , n43840 , n43841 , n43842 ,
     n43843 , n43844 , n43845 , n43846 , n43847 , n43848 , n43849 , n43850 , n43851 , n43852 ,
     n43853 , n43854 , n43855 , n43856 , n43857 , n43858 , n43859 , n43860 , n43861 , n43862 ,
     n43863 , n43864 , n43865 , n43866 , n43867 , n43868 , n43869 , n43870 , n43871 , n43872 ,
     n43873 , n43874 , n43875 , n43876 , n43877 , n43878 , n43879 , n43880 , n43881 , n43882 ,
     n43883 , n43884 , n43885 , n43886 , n43887 , n43888 , n43889 , n43890 , n43891 , n43892 ,
     n43893 , n43894 , n43895 , n43896 , n43897 , n43898 , n43899 , n43900 , n43901 , n43902 ,
     n43903 , n43904 , n43905 , n43906 , n43907 , n43908 , n43909 , n43910 , n43911 , n43912 ,
     n43913 , n43914 , n43915 , n43916 , n43917 , n43918 , n43919 , n43920 , n43921 , n43922 ,
     n43923 , n43924 , n43925 , n43926 , n43927 , n43928 , n43929 , n43930 , n43931 , n43932 ,
     n43933 , n43934 , n43935 , n43936 , n43937 , n43938 , n43939 , n43940 , n43941 , n43942 ,
     n43943 , n43944 , n43945 , n43946 , n43947 , n43948 , n43949 , n43950 , n43951 , n43952 ,
     n43953 , n43954 , n43955 , n43956 , n43957 , n43958 , n43959 , n43960 , n43961 , n43962 ,
     n43963 , n43964 , n43965 , n43966 , n43967 , n43968 , n43969 , n43970 , n43971 , n43972 ,
     n43973 , n43974 , n43975 , n43976 , n43977 , n43978 , n43979 , n43980 , n43981 , n43982 ,
     n43983 , n43984 , n43985 , n43986 , n43987 , n43988 , n43989 , n43990 , n43991 , n43992 ,
     n43993 , n43994 , n43995 , n43996 , n43997 , n43998 , n43999 , n44000 , n44001 , n44002 ,
     n44003 , n44004 , n44005 , n44006 , n44007 , n44008 , n44009 , n44010 , n44011 , n44012 ,
     n44013 , n44014 , n44015 , n44016 , n44017 , n44018 , n44019 , n44020 , n44021 , n44022 ,
     n44023 , n44024 , n44025 , n44026 , n44027 , n44028 , n44029 , n44030 , n44031 , n44032 ,
     n44033 , n44034 , n44035 , n44036 , n44037 , n44038 , n44039 , n44040 , n44041 , n44042 ,
     n44043 , n44044 , n44045 , n44046 , n44047 , n44048 , n44049 , n44050 , n44051 , n44052 ,
     n44053 , n44054 , n44055 , n44056 , n44057 , n44058 , n44059 , n44060 , n44061 , n44062 ,
     n44063 , n44064 , n44065 , n44066 , n44067 , n44068 , n44069 , n44070 , n44071 , n44072 ,
     n44073 , n44074 , n44075 , n44076 , n44077 , n44078 , n44079 , n44080 , n44081 , n44082 ,
     n44083 , n44084 , n44085 , n44086 , n44087 , n44088 , n44089 , n44090 , n44091 , n44092 ,
     n44093 , n44094 , n44095 , n44096 , n44097 , n44098 , n44099 , n44100 , n44101 , n44102 ,
     n44103 , n44104 , n44105 , n44106 , n44107 , n44108 , n44109 , n44110 , n44111 , n44112 ,
     n44113 , n44114 , n44115 , n44116 , n44117 , n44118 , n44119 , n44120 , n44121 , n44122 ,
     n44123 , n44124 , n44125 , n44126 , n44127 , n44128 , n44129 , n44130 , n44131 , n44132 ,
     n44133 , n44134 , n44135 , n44136 , n44137 , n44138 , n44139 , n44140 , n44141 , n44142 ,
     n44143 , n44144 , n44145 , n44146 , n44147 , n44148 , n44149 , n44150 , n44151 , n44152 ,
     n44153 , n44154 , n44155 , n44156 , n44157 , n44158 , n44159 , n44160 , n44161 , n44162 ,
     n44163 , n44164 , n44165 , n44166 , n44167 , n44168 , n44169 , n44170 , n44171 , n44172 ,
     n44173 , n44174 , n44175 , n44176 , n44177 , n44178 , n44179 , n44180 , n44181 , n44182 ,
     n44183 , n44184 , n44185 , n44186 , n44187 , n44188 , n44189 , n44190 , n44191 , n44192 ,
     n44193 , n44194 , n44195 , n44196 , n44197 , n44198 , n44199 , n44200 , n44201 , n44202 ,
     n44203 , n44204 , n44205 , n44206 , n44207 , n44208 , n44209 , n44210 , n44211 , n44212 ,
     n44213 , n44214 , n44215 , n44216 , n44217 , n44218 , n44219 , n44220 , n44221 , n44222 ,
     n44223 , n44224 , n44225 , n44226 , n44227 , n44228 , n44229 , n44230 , n44231 , n44232 ,
     n44233 , n44234 , n44235 , n44236 , n44237 , n44238 , n44239 , n44240 , n44241 , n44242 ,
     n44243 , n44244 , n44245 , n44246 , n44247 , n44248 , n44249 , n44250 , n44251 , n44252 ,
     n44253 , n44254 , n44255 , n44256 , n44257 , n44258 , n44259 , n44260 , n44261 , n44262 ,
     n44263 , n44264 , n44265 , n44266 , n44267 , n44268 , n44269 , n44270 , n44271 , n44272 ,
     n44273 , n44274 , n44275 , n44276 , n44277 , n44278 , n44279 , n44280 , n44281 , n44282 ,
     n44283 , n44284 , n44285 , n44286 , n44287 , n44288 , n44289 , n44290 , n44291 , n44292 ,
     n44293 , n44294 , n44295 , n44296 , n44297 , n44298 , n44299 , n44300 , n44301 , n44302 ,
     n44303 , n44304 , n44305 , n44306 , n44307 , n44308 , n44309 , n44310 , n44311 , n44312 ,
     n44313 , n44314 , n44315 , n44316 , n44317 , n44318 , n44319 , n44320 , n44321 , n44322 ,
     n44323 , n44324 , n44325 , n44326 , n44327 , n44328 , n44329 , n44330 , n44331 , n44332 ,
     n44333 , n44334 , n44335 , n44336 , n44337 , n44338 , n44339 , n44340 , n44341 , n44342 ,
     n44343 , n44344 , n44345 , n44346 , n44347 , n44348 , n44349 , n44350 , n44351 , n44352 ,
     n44353 , n44354 , n44355 , n44356 , n44357 , n44358 , n44359 , n44360 , n44361 , n44362 ,
     n44363 , n44364 , n44365 , n44366 , n44367 , n44368 , n44369 , n44370 , n44371 , n44372 ,
     n44373 , n44374 , n44375 , n44376 , n44377 , n44378 , n44379 , n44380 , n44381 , n44382 ,
     n44383 , n44384 , n44385 , n44386 , n44387 , n44388 , n44389 , n44390 , n44391 , n44392 ,
     n44393 , n44394 , n44395 , n44396 , n44397 , n44398 , n44399 , n44400 , n44401 , n44402 ,
     n44403 , n44404 , n44405 , n44406 , n44407 , n44408 , n44409 , n44410 , n44411 , n44412 ,
     n44413 , n44414 , n44415 , n44416 , n44417 , n44418 , n44419 , n44420 , n44421 , n44422 ,
     n44423 , n44424 , n44425 , n44426 , n44427 , n44428 , n44429 , n44430 , n44431 , n44432 ,
     n44433 , n44434 , n44435 , n44436 , n44437 , n44438 , n44439 , n44440 , n44441 , n44442 ,
     n44443 , n44444 , n44445 , n44446 , n44447 , n44448 , n44449 , n44450 , n44451 , n44452 ,
     n44453 , n44454 , n44455 , n44456 , n44457 , n44458 , n44459 , n44460 , n44461 , n44462 ,
     n44463 , n44464 , n44465 , n44466 , n44467 , n44468 , n44469 , n44470 , n44471 , n44472 ,
     n44473 , n44474 , n44475 , n44476 , n44477 , n44478 , n44479 , n44480 , n44481 , n44482 ,
     n44483 , n44484 , n44485 , n44486 , n44487 , n44488 , n44489 , n44490 , n44491 , n44492 ,
     n44493 , n44494 , n44495 , n44496 , n44497 , n44498 , n44499 , n44500 , n44501 , n44502 ,
     n44503 , n44504 , n44505 , n44506 , n44507 , n44508 , n44509 , n44510 , n44511 , n44512 ,
     n44513 , n44514 , n44515 , n44516 , n44517 , n44518 , n44519 , n44520 , n44521 , n44522 ,
     n44523 , n44524 , n44525 , n44526 , n44527 , n44528 , n44529 , n44530 , n44531 , n44532 ,
     n44533 , n44534 , n44535 , n44536 , n44537 , n44538 , n44539 , n44540 , n44541 , n44542 ,
     n44543 , n44544 , n44545 , n44546 , n44547 , n44548 , n44549 , n44550 , n44551 , n44552 ,
     n44553 , n44554 , n44555 , n44556 , n44557 , n44558 , n44559 , n44560 , n44561 , n44562 ,
     n44563 , n44564 , n44565 , n44566 , n44567 , n44568 , n44569 , n44570 , n44571 , n44572 ,
     n44573 , n44574 , n44575 , n44576 , n44577 , n44578 , n44579 , n44580 , n44581 , n44582 ,
     n44583 , n44584 , n44585 , n44586 , n44587 , n44588 , n44589 , n44590 , n44591 , n44592 ,
     n44593 , n44594 , n44595 , n44596 , n44597 , n44598 , n44599 , n44600 , n44601 , n44602 ,
     n44603 , n44604 , n44605 , n44606 , n44607 , n44608 , n44609 , n44610 , n44611 , n44612 ,
     n44613 , n44614 , n44615 , n44616 , n44617 , n44618 , n44619 , n44620 , n44621 , n44622 ,
     n44623 , n44624 , n44625 , n44626 , n44627 , n44628 , n44629 , n44630 , n44631 , n44632 ,
     n44633 , n44634 , n44635 , n44636 , n44637 , n44638 , n44639 , n44640 , n44641 , n44642 ,
     n44643 , n44644 , n44645 , n44646 , n44647 , n44648 , n44649 , n44650 , n44651 , n44652 ,
     n44653 , n44654 , n44655 , n44656 , n44657 , n44658 , n44659 , n44660 , n44661 , n44662 ,
     n44663 , n44664 , n44665 , n44666 , n44667 , n44668 , n44669 , n44670 , n44671 , n44672 ,
     n44673 , n44674 , n44675 , n44676 , n44677 , n44678 , n44679 , n44680 , n44681 , n44682 ,
     n44683 , n44684 , n44685 , n44686 , n44687 , n44688 , n44689 , n44690 , n44691 , n44692 ,
     n44693 , n44694 , n44695 , n44696 , n44697 , n44698 , n44699 , n44700 , n44701 , n44702 ,
     n44703 , n44704 , n44705 , n44706 , n44707 , n44708 , n44709 , n44710 , n44711 , n44712 ,
     n44713 , n44714 , n44715 , n44716 , n44717 , n44718 , n44719 , n44720 , n44721 , n44722 ,
     n44723 , n44724 , n44725 , n44726 , n44727 , n44728 , n44729 , n44730 , n44731 , n44732 ,
     n44733 , n44734 , n44735 , n44736 , n44737 , n44738 , n44739 , n44740 , n44741 , n44742 ,
     n44743 , n44744 , n44745 , n44746 , n44747 , n44748 , n44749 , n44750 , n44751 , n44752 ,
     n44753 , n44754 , n44755 , n44756 , n44757 , n44758 , n44759 , n44760 , n44761 , n44762 ,
     n44763 , n44764 , n44765 , n44766 , n44767 , n44768 , n44769 , n44770 , n44771 , n44772 ,
     n44773 , n44774 , n44775 , n44776 , n44777 , n44778 , n44779 , n44780 , n44781 , n44782 ,
     n44783 , n44784 , n44785 , n44786 , n44787 , n44788 , n44789 , n44790 , n44791 , n44792 ,
     n44793 , n44794 , n44795 , n44796 , n44797 , n44798 , n44799 , n44800 , n44801 , n44802 ,
     n44803 , n44804 , n44805 , n44806 , n44807 , n44808 , n44809 , n44810 , n44811 , n44812 ,
     n44813 , n44814 , n44815 , n44816 , n44817 , n44818 , n44819 , n44820 , n44821 , n44822 ,
     n44823 , n44824 , n44825 , n44826 , n44827 , n44828 , n44829 , n44830 , n44831 , n44832 ,
     n44833 , n44834 , n44835 , n44836 , n44837 , n44838 , n44839 , n44840 , n44841 , n44842 ,
     n44843 , n44844 , n44845 , n44846 , n44847 , n44848 , n44849 , n44850 , n44851 , n44852 ,
     n44853 , n44854 , n44855 , n44856 , n44857 , n44858 , n44859 , n44860 , n44861 , n44862 ,
     n44863 , n44864 , n44865 , n44866 , n44867 , n44868 , n44869 , n44870 , n44871 , n44872 ,
     n44873 , n44874 , n44875 , n44876 , n44877 , n44878 , n44879 , n44880 , n44881 , n44882 ,
     n44883 , n44884 , n44885 , n44886 , n44887 , n44888 , n44889 , n44890 , n44891 , n44892 ,
     n44893 , n44894 , n44895 , n44896 , n44897 , n44898 , n44899 , n44900 , n44901 , n44902 ,
     n44903 , n44904 , n44905 , n44906 , n44907 , n44908 , n44909 , n44910 , n44911 , n44912 ,
     n44913 , n44914 , n44915 , n44916 , n44917 , n44918 , n44919 , n44920 , n44921 , n44922 ,
     n44923 , n44924 , n44925 , n44926 , n44927 , n44928 , n44929 , n44930 , n44931 , n44932 ,
     n44933 , n44934 , n44935 , n44936 , n44937 , n44938 , n44939 , n44940 , n44941 , n44942 ,
     n44943 , n44944 , n44945 , n44946 , n44947 , n44948 , n44949 , n44950 , n44951 , n44952 ,
     n44953 , n44954 , n44955 , n44956 , n44957 , n44958 , n44959 , n44960 , n44961 , n44962 ,
     n44963 , n44964 , n44965 , n44966 , n44967 , n44968 , n44969 , n44970 , n44971 , n44972 ,
     n44973 , n44974 , n44975 , n44976 , n44977 , n44978 , n44979 , n44980 , n44981 , n44982 ,
     n44983 , n44984 , n44985 , n44986 , n44987 , n44988 , n44989 , n44990 , n44991 , n44992 ,
     n44993 , n44994 , n44995 , n44996 , n44997 , n44998 , n44999 , n45000 , n45001 , n45002 ,
     n45003 , n45004 , n45005 , n45006 , n45007 , n45008 , n45009 , n45010 , n45011 , n45012 ,
     n45013 , n45014 , n45015 , n45016 , n45017 , n45018 , n45019 , n45020 , n45021 , n45022 ,
     n45023 , n45024 , n45025 , n45026 , n45027 , n45028 , n45029 , n45030 , n45031 , n45032 ,
     n45033 , n45034 , n45035 , n45036 , n45037 , n45038 , n45039 , n45040 , n45041 , n45042 ,
     n45043 , n45044 , n45045 , n45046 , n45047 , n45048 , n45049 , n45050 , n45051 , n45052 ,
     n45053 , n45054 , n45055 , n45056 , n45057 , n45058 , n45059 , n45060 , n45061 , n45062 ,
     n45063 , n45064 , n45065 , n45066 , n45067 , n45068 , n45069 , n45070 , n45071 , n45072 ,
     n45073 , n45074 , n45075 , n45076 , n45077 , n45078 , n45079 , n45080 , n45081 , n45082 ,
     n45083 , n45084 , n45085 , n45086 , n45087 , n45088 , n45089 , n45090 , n45091 , n45092 ,
     n45093 , n45094 , n45095 , n45096 , n45097 , n45098 , n45099 , n45100 , n45101 , n45102 ,
     n45103 , n45104 , n45105 , n45106 , n45107 , n45108 , n45109 , n45110 , n45111 , n45112 ,
     n45113 , n45114 , n45115 , n45116 , n45117 , n45118 , n45119 , n45120 , n45121 , n45122 ,
     n45123 , n45124 , n45125 , n45126 , n45127 , n45128 , n45129 , n45130 , n45131 , n45132 ,
     n45133 , n45134 , n45135 , n45136 , n45137 , n45138 , n45139 , n45140 , n45141 , n45142 ,
     n45143 , n45144 , n45145 , n45146 , n45147 , n45148 , n45149 , n45150 , n45151 , n45152 ,
     n45153 , n45154 , n45155 , n45156 , n45157 , n45158 , n45159 , n45160 , n45161 , n45162 ,
     n45163 , n45164 , n45165 , n45166 , n45167 , n45168 , n45169 , n45170 , n45171 , n45172 ,
     n45173 , n45174 , n45175 , n45176 , n45177 , n45178 , n45179 , n45180 , n45181 , n45182 ,
     n45183 , n45184 , n45185 , n45186 , n45187 , n45188 , n45189 , n45190 , n45191 , n45192 ,
     n45193 , n45194 , n45195 , n45196 , n45197 , n45198 , n45199 , n45200 , n45201 , n45202 ,
     n45203 , n45204 , n45205 , n45206 , n45207 , n45208 , n45209 , n45210 , n45211 , n45212 ,
     n45213 , n45214 , n45215 , n45216 , n45217 , n45218 , n45219 , n45220 , n45221 , n45222 ,
     n45223 , n45224 , n45225 , n45226 , n45227 , n45228 , n45229 , n45230 , n45231 , n45232 ,
     n45233 , n45234 , n45235 , n45236 , n45237 , n45238 , n45239 , n45240 , n45241 , n45242 ,
     n45243 , n45244 , n45245 , n45246 , n45247 , n45248 , n45249 , n45250 , n45251 , n45252 ,
     n45253 , n45254 , n45255 , n45256 , n45257 , n45258 , n45259 , n45260 , n45261 , n45262 ,
     n45263 , n45264 , n45265 , n45266 , n45267 , n45268 , n45269 , n45270 , n45271 , n45272 ,
     n45273 , n45274 , n45275 , n45276 , n45277 , n45278 , n45279 , n45280 , n45281 , n45282 ,
     n45283 , n45284 , n45285 , n45286 , n45287 , n45288 , n45289 , n45290 , n45291 , n45292 ,
     n45293 , n45294 , n45295 , n45296 , n45297 , n45298 , n45299 , n45300 , n45301 , n45302 ,
     n45303 , n45304 , n45305 , n45306 , n45307 , n45308 , n45309 , n45310 , n45311 , n45312 ,
     n45313 , n45314 , n45315 , n45316 , n45317 , n45318 , n45319 , n45320 , n45321 , n45322 ,
     n45323 , n45324 , n45325 , n45326 , n45327 , n45328 , n45329 , n45330 , n45331 , n45332 ,
     n45333 , n45334 , n45335 , n45336 , n45337 , n45338 , n45339 , n45340 , n45341 , n45342 ,
     n45343 , n45344 , n45345 , n45346 , n45347 , n45348 , n45349 , n45350 , n45351 , n45352 ,
     n45353 , n45354 , n45355 , n45356 , n45357 , n45358 , n45359 , n45360 , n45361 , n45362 ,
     n45363 , n45364 , n45365 , n45366 , n45367 , n45368 , n45369 , n45370 , n45371 , n45372 ,
     n45373 , n45374 , n45375 , n45376 , n45377 , n45378 , n45379 , n45380 , n45381 , n45382 ,
     n45383 , n45384 , n45385 , n45386 , n45387 , n45388 , n45389 , n45390 , n45391 , n45392 ,
     n45393 , n45394 , n45395 , n45396 , n45397 , n45398 , n45399 , n45400 , n45401 , n45402 ,
     n45403 , n45404 , n45405 , n45406 , n45407 , n45408 , n45409 , n45410 , n45411 , n45412 ,
     n45413 , n45414 , n45415 , n45416 , n45417 , n45418 , n45419 , n45420 , n45421 , n45422 ,
     n45423 , n45424 , n45425 , n45426 , n45427 , n45428 , n45429 , n45430 , n45431 , n45432 ,
     n45433 , n45434 , n45435 , n45436 , n45437 , n45438 , n45439 , n45440 , n45441 , n45442 ,
     n45443 , n45444 , n45445 , n45446 , n45447 , n45448 , n45449 , n45450 , n45451 , n45452 ,
     n45453 , n45454 , n45455 , n45456 , n45457 , n45458 , n45459 , n45460 , n45461 , n45462 ,
     n45463 , n45464 , n45465 , n45466 , n45467 , n45468 , n45469 , n45470 , n45471 , n45472 ,
     n45473 , n45474 , n45475 , n45476 , n45477 , n45478 , n45479 , n45480 , n45481 , n45482 ,
     n45483 , n45484 , n45485 , n45486 , n45487 , n45488 , n45489 , n45490 , n45491 , n45492 ,
     n45493 , n45494 , n45495 , n45496 , n45497 , n45498 , n45499 , n45500 , n45501 , n45502 ,
     n45503 , n45504 , n45505 , n45506 , n45507 , n45508 , n45509 , n45510 , n45511 , n45512 ,
     n45513 , n45514 , n45515 , n45516 , n45517 , n45518 , n45519 , n45520 , n45521 , n45522 ,
     n45523 , n45524 , n45525 , n45526 , n45527 , n45528 , n45529 , n45530 , n45531 , n45532 ,
     n45533 , n45534 , n45535 , n45536 , n45537 , n45538 , n45539 , n45540 , n45541 , n45542 ,
     n45543 , n45544 , n45545 , n45546 , n45547 , n45548 , n45549 , n45550 , n45551 , n45552 ,
     n45553 , n45554 , n45555 , n45556 , n45557 , n45558 , n45559 , n45560 , n45561 , n45562 ,
     n45563 , n45564 , n45565 , n45566 , n45567 , n45568 , n45569 , n45570 , n45571 , n45572 ,
     n45573 , n45574 , n45575 , n45576 , n45577 , n45578 , n45579 , n45580 , n45581 , n45582 ,
     n45583 , n45584 , n45585 , n45586 , n45587 , n45588 , n45589 , n45590 , n45591 , n45592 ,
     n45593 , n45594 , n45595 , n45596 , n45597 , n45598 , n45599 , n45600 , n45601 , n45602 ,
     n45603 , n45604 , n45605 , n45606 , n45607 , n45608 , n45609 , n45610 , n45611 , n45612 ,
     n45613 , n45614 , n45615 , n45616 , n45617 , n45618 , n45619 , n45620 , n45621 , n45622 ,
     n45623 , n45624 , n45625 , n45626 , n45627 , n45628 , n45629 , n45630 , n45631 , n45632 ,
     n45633 , n45634 , n45635 , n45636 , n45637 , n45638 , n45639 , n45640 , n45641 , n45642 ,
     n45643 , n45644 , n45645 , n45646 , n45647 , n45648 , n45649 , n45650 , n45651 , n45652 ,
     n45653 , n45654 , n45655 , n45656 , n45657 , n45658 , n45659 , n45660 , n45661 , n45662 ,
     n45663 , n45664 , n45665 , n45666 , n45667 , n45668 , n45669 , n45670 , n45671 , n45672 ,
     n45673 , n45674 , n45675 , n45676 , n45677 , n45678 , n45679 , n45680 , n45681 , n45682 ,
     n45683 , n45684 , n45685 , n45686 , n45687 , n45688 , n45689 , n45690 , n45691 , n45692 ,
     n45693 , n45694 , n45695 , n45696 , n45697 , n45698 , n45699 , n45700 , n45701 , n45702 ,
     n45703 , n45704 , n45705 , n45706 , n45707 , n45708 , n45709 , n45710 , n45711 , n45712 ,
     n45713 , n45714 , n45715 , n45716 , n45717 , n45718 , n45719 , n45720 , n45721 , n45722 ,
     n45723 , n45724 , n45725 , n45726 , n45727 , n45728 , n45729 , n45730 , n45731 , n45732 ,
     n45733 , n45734 , n45735 , n45736 , n45737 , n45738 , n45739 , n45740 , n45741 , n45742 ,
     n45743 , n45744 , n45745 , n45746 , n45747 , n45748 , n45749 , n45750 , n45751 , n45752 ,
     n45753 , n45754 , n45755 , n45756 , n45757 , n45758 , n45759 , n45760 , n45761 , n45762 ,
     n45763 , n45764 , n45765 , n45766 , n45767 , n45768 , n45769 , n45770 , n45771 , n45772 ,
     n45773 , n45774 , n45775 , n45776 , n45777 , n45778 , n45779 , n45780 , n45781 , n45782 ,
     n45783 , n45784 , n45785 , n45786 , n45787 , n45788 , n45789 , n45790 , n45791 , n45792 ,
     n45793 , n45794 , n45795 , n45796 , n45797 , n45798 , n45799 , n45800 , n45801 , n45802 ,
     n45803 , n45804 , n45805 , n45806 , n45807 , n45808 , n45809 , n45810 , n45811 , n45812 ,
     n45813 , n45814 , n45815 , n45816 , n45817 , n45818 , n45819 , n45820 , n45821 , n45822 ,
     n45823 , n45824 , n45825 , n45826 , n45827 , n45828 , n45829 , n45830 , n45831 , n45832 ,
     n45833 , n45834 , n45835 , n45836 , n45837 , n45838 , n45839 , n45840 , n45841 , n45842 ,
     n45843 , n45844 , n45845 , n45846 , n45847 , n45848 , n45849 , n45850 , n45851 , n45852 ,
     n45853 , n45854 , n45855 , n45856 , n45857 , n45858 , n45859 , n45860 , n45861 , n45862 ,
     n45863 , n45864 , n45865 , n45866 , n45867 , n45868 , n45869 , n45870 , n45871 , n45872 ,
     n45873 , n45874 , n45875 , n45876 , n45877 , n45878 , n45879 , n45880 , n45881 , n45882 ,
     n45883 , n45884 , n45885 , n45886 , n45887 , n45888 , n45889 , n45890 , n45891 , n45892 ,
     n45893 , n45894 , n45895 , n45896 , n45897 , n45898 , n45899 , n45900 , n45901 , n45902 ,
     n45903 , n45904 , n45905 , n45906 , n45907 , n45908 , n45909 , n45910 , n45911 , n45912 ,
     n45913 , n45914 , n45915 , n45916 , n45917 , n45918 , n45919 , n45920 , n45921 , n45922 ,
     n45923 , n45924 , n45925 , n45926 , n45927 , n45928 , n45929 , n45930 , n45931 , n45932 ,
     n45933 , n45934 , n45935 , n45936 , n45937 , n45938 , n45939 , n45940 , n45941 , n45942 ,
     n45943 , n45944 , n45945 , n45946 , n45947 , n45948 , n45949 , n45950 , n45951 , n45952 ,
     n45953 , n45954 , n45955 , n45956 , n45957 , n45958 , n45959 , n45960 , n45961 , n45962 ,
     n45963 , n45964 , n45965 , n45966 , n45967 , n45968 , n45969 , n45970 , n45971 , n45972 ,
     n45973 , n45974 , n45975 , n45976 , n45977 , n45978 , n45979 , n45980 , n45981 , n45982 ,
     n45983 , n45984 , n45985 , n45986 , n45987 , n45988 , n45989 , n45990 , n45991 , n45992 ,
     n45993 , n45994 , n45995 , n45996 , n45997 , n45998 , n45999 , n46000 , n46001 , n46002 ,
     n46003 , n46004 , n46005 , n46006 , n46007 , n46008 , n46009 , n46010 , n46011 , n46012 ,
     n46013 , n46014 , n46015 , n46016 , n46017 , n46018 , n46019 , n46020 , n46021 , n46022 ,
     n46023 , n46024 , n46025 , n46026 , n46027 , n46028 , n46029 , n46030 , n46031 , n46032 ,
     n46033 , n46034 , n46035 , n46036 , n46037 , n46038 , n46039 , n46040 , n46041 , n46042 ,
     n46043 , n46044 , n46045 , n46046 , n46047 , n46048 , n46049 , n46050 , n46051 , n46052 ,
     n46053 , n46054 , n46055 , n46056 , n46057 , n46058 , n46059 , n46060 , n46061 , n46062 ,
     n46063 , n46064 , n46065 , n46066 , n46067 , n46068 , n46069 , n46070 , n46071 , n46072 ,
     n46073 , n46074 , n46075 , n46076 , n46077 , n46078 , n46079 , n46080 , n46081 , n46082 ,
     n46083 , n46084 , n46085 , n46086 , n46087 , n46088 , n46089 , n46090 , n46091 , n46092 ,
     n46093 , n46094 , n46095 , n46096 , n46097 , n46098 , n46099 , n46100 , n46101 , n46102 ,
     n46103 , n46104 , n46105 , n46106 , n46107 , n46108 , n46109 , n46110 , n46111 , n46112 ,
     n46113 , n46114 , n46115 , n46116 , n46117 , n46118 , n46119 , n46120 , n46121 , n46122 ,
     n46123 , n46124 , n46125 , n46126 , n46127 , n46128 , n46129 , n46130 , n46131 , n46132 ,
     n46133 , n46134 , n46135 , n46136 , n46137 , n46138 , n46139 , n46140 , n46141 , n46142 ,
     n46143 , n46144 , n46145 , n46146 , n46147 , n46148 , n46149 , n46150 , n46151 , n46152 ,
     n46153 , n46154 , n46155 , n46156 , n46157 , n46158 , n46159 , n46160 , n46161 , n46162 ,
     n46163 , n46164 , n46165 , n46166 , n46167 , n46168 , n46169 , n46170 , n46171 , n46172 ,
     n46173 , n46174 , n46175 , n46176 , n46177 , n46178 , n46179 , n46180 , n46181 , n46182 ,
     n46183 , n46184 , n46185 , n46186 , n46187 , n46188 , n46189 , n46190 , n46191 , n46192 ,
     n46193 , n46194 , n46195 , n46196 , n46197 , n46198 , n46199 , n46200 , n46201 , n46202 ,
     n46203 , n46204 , n46205 , n46206 , n46207 , n46208 , n46209 , n46210 , n46211 , n46212 ,
     n46213 , n46214 , n46215 , n46216 , n46217 , n46218 , n46219 , n46220 , n46221 , n46222 ,
     n46223 , n46224 , n46225 , n46226 , n46227 , n46228 , n46229 , n46230 , n46231 , n46232 ,
     n46233 , n46234 , n46235 , n46236 , n46237 , n46238 , n46239 , n46240 , n46241 , n46242 ,
     n46243 , n46244 , n46245 , n46246 , n46247 , n46248 , n46249 , n46250 , n46251 , n46252 ,
     n46253 , n46254 , n46255 , n46256 , n46257 , n46258 , n46259 , n46260 , n46261 , n46262 ,
     n46263 , n46264 , n46265 , n46266 , n46267 , n46268 , n46269 , n46270 , n46271 , n46272 ,
     n46273 , n46274 , n46275 , n46276 , n46277 , n46278 , n46279 , n46280 , n46281 , n46282 ,
     n46283 , n46284 , n46285 , n46286 , n46287 , n46288 , n46289 , n46290 , n46291 , n46292 ,
     n46293 , n46294 , n46295 , n46296 , n46297 , n46298 , n46299 , n46300 , n46301 , n46302 ,
     n46303 , n46304 , n46305 , n46306 , n46307 , n46308 , n46309 , n46310 , n46311 , n46312 ,
     n46313 , n46314 , n46315 , n46316 , n46317 , n46318 , n46319 , n46320 , n46321 , n46322 ,
     n46323 , n46324 , n46325 , n46326 , n46327 , n46328 , n46329 , n46330 , n46331 , n46332 ,
     n46333 , n46334 , n46335 , n46336 , n46337 , n46338 , n46339 , n46340 , n46341 , n46342 ,
     n46343 , n46344 , n46345 , n46346 , n46347 , n46348 , n46349 , n46350 , n46351 , n46352 ,
     n46353 , n46354 , n46355 , n46356 , n46357 , n46358 , n46359 , n46360 , n46361 , n46362 ,
     n46363 , n46364 , n46365 , n46366 , n46367 , n46368 , n46369 , n46370 , n46371 , n46372 ,
     n46373 , n46374 , n46375 , n46376 , n46377 , n46378 , n46379 , n46380 , n46381 , n46382 ,
     n46383 , n46384 , n46385 , n46386 , n46387 , n46388 , n46389 , n46390 , n46391 , n46392 ,
     n46393 , n46394 , n46395 , n46396 , n46397 , n46398 , n46399 , n46400 , n46401 , n46402 ,
     n46403 , n46404 , n46405 , n46406 , n46407 , n46408 , n46409 , n46410 , n46411 , n46412 ,
     n46413 , n46414 , n46415 , n46416 , n46417 , n46418 , n46419 , n46420 , n46421 , n46422 ,
     n46423 , n46424 , n46425 , n46426 , n46427 , n46428 , n46429 , n46430 , n46431 , n46432 ,
     n46433 , n46434 , n46435 , n46436 , n46437 , n46438 , n46439 , n46440 , n46441 , n46442 ,
     n46443 , n46444 , n46445 , n46446 , n46447 , n46448 , n46449 , n46450 , n46451 , n46452 ,
     n46453 , n46454 , n46455 , n46456 , n46457 , n46458 , n46459 , n46460 , n46461 , n46462 ,
     n46463 , n46464 , n46465 , n46466 , n46467 , n46468 , n46469 , n46470 , n46471 , n46472 ,
     n46473 , n46474 , n46475 , n46476 , n46477 , n46478 , n46479 , n46480 , n46481 , n46482 ,
     n46483 , n46484 , n46485 , n46486 , n46487 , n46488 , n46489 , n46490 , n46491 , n46492 ,
     n46493 , n46494 , n46495 , n46496 , n46497 , n46498 , n46499 , n46500 , n46501 , n46502 ,
     n46503 , n46504 , n46505 , n46506 , n46507 , n46508 , n46509 , n46510 , n46511 , n46512 ,
     n46513 , n46514 , n46515 , n46516 , n46517 , n46518 , n46519 , n46520 , n46521 , n46522 ,
     n46523 , n46524 , n46525 , n46526 , n46527 , n46528 , n46529 , n46530 , n46531 , n46532 ,
     n46533 , n46534 , n46535 , n46536 , n46537 , n46538 , n46539 , n46540 , n46541 , n46542 ,
     n46543 , n46544 , n46545 , n46546 , n46547 , n46548 , n46549 , n46550 , n46551 , n46552 ,
     n46553 , n46554 , n46555 , n46556 , n46557 , n46558 , n46559 , n46560 , n46561 , n46562 ,
     n46563 , n46564 , n46565 , n46566 , n46567 , n46568 , n46569 , n46570 , n46571 , n46572 ,
     n46573 , n46574 , n46575 , n46576 , n46577 , n46578 , n46579 , n46580 , n46581 , n46582 ,
     n46583 , n46584 , n46585 , n46586 , n46587 , n46588 , n46589 , n46590 , n46591 , n46592 ,
     n46593 , n46594 , n46595 , n46596 , n46597 , n46598 , n46599 , n46600 , n46601 , n46602 ,
     n46603 , n46604 , n46605 , n46606 , n46607 , n46608 , n46609 , n46610 , n46611 , n46612 ,
     n46613 , n46614 , n46615 , n46616 , n46617 , n46618 , n46619 , n46620 , n46621 , n46622 ,
     n46623 , n46624 , n46625 , n46626 , n46627 , n46628 , n46629 , n46630 , n46631 , n46632 ,
     n46633 , n46634 , n46635 , n46636 , n46637 , n46638 , n46639 , n46640 , n46641 , n46642 ,
     n46643 , n46644 , n46645 , n46646 , n46647 , n46648 , n46649 , n46650 , n46651 , n46652 ,
     n46653 , n46654 , n46655 , n46656 , n46657 , n46658 , n46659 , n46660 , n46661 , n46662 ,
     n46663 , n46664 , n46665 , n46666 , n46667 , n46668 , n46669 , n46670 , n46671 , n46672 ,
     n46673 , n46674 , n46675 , n46676 , n46677 , n46678 , n46679 , n46680 , n46681 , n46682 ,
     n46683 , n46684 , n46685 , n46686 , n46687 , n46688 , n46689 , n46690 , n46691 , n46692 ,
     n46693 , n46694 , n46695 , n46696 , n46697 , n46698 , n46699 , n46700 , n46701 , n46702 ,
     n46703 , n46704 , n46705 , n46706 , n46707 , n46708 , n46709 , n46710 , n46711 , n46712 ,
     n46713 , n46714 , n46715 , n46716 , n46717 , n46718 , n46719 , n46720 , n46721 , n46722 ,
     n46723 , n46724 , n46725 , n46726 , n46727 , n46728 , n46729 , n46730 , n46731 , n46732 ,
     n46733 , n46734 , n46735 , n46736 , n46737 , n46738 , n46739 , n46740 , n46741 , n46742 ,
     n46743 , n46744 , n46745 , n46746 , n46747 , n46748 , n46749 , n46750 , n46751 , n46752 ,
     n46753 , n46754 , n46755 , n46756 , n46757 , n46758 , n46759 , n46760 , n46761 , n46762 ,
     n46763 , n46764 , n46765 , n46766 , n46767 , n46768 , n46769 , n46770 , n46771 , n46772 ,
     n46773 , n46774 , n46775 , n46776 , n46777 , n46778 , n46779 , n46780 , n46781 , n46782 ,
     n46783 , n46784 , n46785 , n46786 , n46787 , n46788 , n46789 , n46790 , n46791 , n46792 ,
     n46793 , n46794 , n46795 , n46796 , n46797 , n46798 , n46799 , n46800 , n46801 , n46802 ,
     n46803 , n46804 , n46805 , n46806 , n46807 , n46808 , n46809 , n46810 , n46811 , n46812 ,
     n46813 , n46814 , n46815 , n46816 , n46817 , n46818 , n46819 , n46820 , n46821 , n46822 ,
     n46823 , n46824 , n46825 , n46826 , n46827 , n46828 , n46829 , n46830 , n46831 , n46832 ,
     n46833 , n46834 , n46835 , n46836 , n46837 , n46838 , n46839 , n46840 , n46841 , n46842 ,
     n46843 , n46844 , n46845 , n46846 , n46847 , n46848 , n46849 , n46850 , n46851 , n46852 ,
     n46853 , n46854 , n46855 , n46856 , n46857 , n46858 , n46859 , n46860 , n46861 , n46862 ,
     n46863 , n46864 , n46865 , n46866 , n46867 , n46868 , n46869 , n46870 , n46871 , n46872 ,
     n46873 , n46874 , n46875 , n46876 , n46877 , n46878 , n46879 , n46880 , n46881 , n46882 ,
     n46883 , n46884 , n46885 , n46886 , n46887 , n46888 , n46889 , n46890 , n46891 , n46892 ,
     n46893 , n46894 , n46895 , n46896 , n46897 , n46898 , n46899 , n46900 , n46901 , n46902 ,
     n46903 , n46904 , n46905 , n46906 , n46907 , n46908 , n46909 , n46910 , n46911 , n46912 ,
     n46913 , n46914 , n46915 , n46916 , n46917 , n46918 , n46919 , n46920 , n46921 , n46922 ,
     n46923 , n46924 , n46925 , n46926 , n46927 , n46928 , n46929 , n46930 , n46931 , n46932 ,
     n46933 , n46934 , n46935 , n46936 , n46937 , n46938 , n46939 , n46940 , n46941 , n46942 ,
     n46943 , n46944 , n46945 , n46946 , n46947 , n46948 , n46949 , n46950 , n46951 , n46952 ,
     n46953 , n46954 , n46955 , n46956 , n46957 , n46958 , n46959 , n46960 , n46961 , n46962 ,
     n46963 , n46964 , n46965 , n46966 , n46967 , n46968 , n46969 , n46970 , n46971 , n46972 ,
     n46973 , n46974 , n46975 , n46976 , n46977 , n46978 , n46979 , n46980 , n46981 , n46982 ,
     n46983 , n46984 , n46985 , n46986 , n46987 , n46988 , n46989 , n46990 , n46991 , n46992 ,
     n46993 , n46994 , n46995 , n46996 , n46997 , n46998 , n46999 , n47000 , n47001 , n47002 ,
     n47003 , n47004 , n47005 , n47006 , n47007 , n47008 , n47009 , n47010 , n47011 , n47012 ,
     n47013 , n47014 , n47015 , n47016 , n47017 , n47018 , n47019 , n47020 , n47021 , n47022 ,
     n47023 , n47024 , n47025 , n47026 , n47027 , n47028 , n47029 , n47030 , n47031 , n47032 ,
     n47033 , n47034 , n47035 , n47036 , n47037 , n47038 , n47039 , n47040 , n47041 , n47042 ,
     n47043 , n47044 , n47045 , n47046 , n47047 , n47048 , n47049 , n47050 , n47051 , n47052 ,
     n47053 , n47054 , n47055 , n47056 , n47057 , n47058 , n47059 , n47060 , n47061 , n47062 ,
     n47063 , n47064 , n47065 , n47066 , n47067 , n47068 , n47069 , n47070 , n47071 , n47072 ,
     n47073 , n47074 , n47075 , n47076 , n47077 , n47078 , n47079 , n47080 , n47081 , n47082 ,
     n47083 , n47084 , n47085 , n47086 , n47087 , n47088 , n47089 , n47090 , n47091 , n47092 ,
     n47093 , n47094 , n47095 , n47096 , n47097 , n47098 , n47099 , n47100 , n47101 , n47102 ,
     n47103 , n47104 , n47105 , n47106 , n47107 , n47108 , n47109 , n47110 , n47111 , n47112 ,
     n47113 , n47114 , n47115 , n47116 , n47117 , n47118 , n47119 , n47120 , n47121 , n47122 ,
     n47123 , n47124 , n47125 , n47126 , n47127 , n47128 , n47129 , n47130 , n47131 , n47132 ,
     n47133 , n47134 , n47135 , n47136 , n47137 , n47138 , n47139 , n47140 , n47141 , n47142 ,
     n47143 , n47144 , n47145 , n47146 , n47147 , n47148 , n47149 , n47150 , n47151 , n47152 ,
     n47153 , n47154 , n47155 , n47156 , n47157 , n47158 , n47159 , n47160 , n47161 , n47162 ,
     n47163 , n47164 , n47165 , n47166 , n47167 , n47168 , n47169 , n47170 , n47171 , n47172 ,
     n47173 , n47174 , n47175 , n47176 , n47177 , n47178 , n47179 , n47180 , n47181 , n47182 ,
     n47183 , n47184 , n47185 , n47186 , n47187 , n47188 , n47189 , n47190 , n47191 , n47192 ,
     n47193 , n47194 , n47195 , n47196 , n47197 , n47198 , n47199 , n47200 , n47201 , n47202 ,
     n47203 , n47204 , n47205 , n47206 , n47207 , n47208 , n47209 , n47210 , n47211 , n47212 ,
     n47213 , n47214 , n47215 , n47216 , n47217 , n47218 , n47219 , n47220 , n47221 , n47222 ,
     n47223 , n47224 , n47225 , n47226 , n47227 , n47228 , n47229 , n47230 , n47231 , n47232 ,
     n47233 , n47234 , n47235 , n47236 , n47237 , n47238 , n47239 , n47240 , n47241 , n47242 ,
     n47243 , n47244 , n47245 , n47246 , n47247 , n47248 , n47249 , n47250 , n47251 , n47252 ,
     n47253 , n47254 , n47255 , n47256 , n47257 , n47258 , n47259 , n47260 , n47261 , n47262 ,
     n47263 , n47264 , n47265 , n47266 , n47267 , n47268 , n47269 , n47270 , n47271 , n47272 ,
     n47273 , n47274 , n47275 , n47276 , n47277 , n47278 , n47279 , n47280 , n47281 , n47282 ,
     n47283 , n47284 , n47285 , n47286 , n47287 , n47288 , n47289 , n47290 , n47291 , n47292 ,
     n47293 , n47294 , n47295 , n47296 , n47297 , n47298 , n47299 , n47300 , n47301 , n47302 ,
     n47303 , n47304 , n47305 , n47306 , n47307 , n47308 , n47309 , n47310 , n47311 , n47312 ,
     n47313 , n47314 , n47315 , n47316 , n47317 , n47318 , n47319 , n47320 , n47321 , n47322 ,
     n47323 , n47324 , n47325 , n47326 , n47327 , n47328 , n47329 , n47330 , n47331 , n47332 ,
     n47333 , n47334 , n47335 , n47336 , n47337 , n47338 , n47339 , n47340 , n47341 , n47342 ,
     n47343 , n47344 , n47345 , n47346 , n47347 , n47348 , n47349 , n47350 , n47351 , n47352 ,
     n47353 , n47354 , n47355 , n47356 , n47357 , n47358 , n47359 , n47360 , n47361 , n47362 ,
     n47363 , n47364 , n47365 , n47366 , n47367 , n47368 , n47369 , n47370 , n47371 , n47372 ,
     n47373 , n47374 , n47375 , n47376 , n47377 , n47378 , n47379 , n47380 , n47381 , n47382 ,
     n47383 , n47384 , n47385 , n47386 , n47387 , n47388 , n47389 , n47390 , n47391 , n47392 ,
     n47393 , n47394 , n47395 , n47396 , n47397 , n47398 , n47399 , n47400 , n47401 , n47402 ,
     n47403 , n47404 , n47405 , n47406 , n47407 , n47408 , n47409 , n47410 , n47411 , n47412 ,
     n47413 , n47414 , n47415 , n47416 , n47417 , n47418 , n47419 , n47420 , n47421 , n47422 ,
     n47423 , n47424 , n47425 , n47426 , n47427 , n47428 , n47429 , n47430 , n47431 , n47432 ,
     n47433 , n47434 , n47435 , n47436 , n47437 , n47438 , n47439 , n47440 , n47441 , n47442 ,
     n47443 , n47444 , n47445 , n47446 , n47447 , n47448 , n47449 , n47450 , n47451 , n47452 ,
     n47453 , n47454 , n47455 , n47456 , n47457 , n47458 , n47459 , n47460 , n47461 , n47462 ,
     n47463 , n47464 , n47465 , n47466 , n47467 , n47468 , n47469 , n47470 , n47471 , n47472 ,
     n47473 , n47474 , n47475 , n47476 , n47477 , n47478 , n47479 , n47480 , n47481 , n47482 ,
     n47483 , n47484 , n47485 , n47486 , n47487 , n47488 , n47489 , n47490 , n47491 , n47492 ,
     n47493 , n47494 , n47495 , n47496 , n47497 , n47498 , n47499 , n47500 , n47501 , n47502 ,
     n47503 , n47504 , n47505 , n47506 , n47507 , n47508 , n47509 , n47510 , n47511 , n47512 ,
     n47513 , n47514 , n47515 , n47516 , n47517 , n47518 , n47519 , n47520 , n47521 , n47522 ,
     n47523 , n47524 , n47525 , n47526 , n47527 , n47528 , n47529 , n47530 , n47531 , n47532 ,
     n47533 , n47534 , n47535 , n47536 , n47537 , n47538 , n47539 , n47540 , n47541 , n47542 ,
     n47543 , n47544 , n47545 , n47546 , n47547 , n47548 , n47549 , n47550 , n47551 , n47552 ,
     n47553 , n47554 , n47555 , n47556 , n47557 , n47558 , n47559 , n47560 , n47561 , n47562 ,
     n47563 , n47564 , n47565 , n47566 , n47567 , n47568 , n47569 , n47570 , n47571 , n47572 ,
     n47573 , n47574 , n47575 , n47576 , n47577 , n47578 , n47579 , n47580 , n47581 , n47582 ,
     n47583 , n47584 , n47585 , n47586 , n47587 , n47588 , n47589 , n47590 , n47591 , n47592 ,
     n47593 , n47594 , n47595 , n47596 , n47597 , n47598 , n47599 , n47600 , n47601 , n47602 ,
     n47603 , n47604 , n47605 , n47606 , n47607 , n47608 , n47609 , n47610 , n47611 , n47612 ,
     n47613 , n47614 , n47615 , n47616 , n47617 , n47618 , n47619 , n47620 , n47621 , n47622 ,
     n47623 , n47624 , n47625 , n47626 , n47627 , n47628 , n47629 , n47630 , n47631 , n47632 ,
     n47633 , n47634 , n47635 , n47636 , n47637 , n47638 , n47639 , n47640 , n47641 , n47642 ,
     n47643 , n47644 , n47645 , n47646 , n47647 , n47648 , n47649 , n47650 , n47651 , n47652 ,
     n47653 , n47654 , n47655 , n47656 , n47657 , n47658 , n47659 , n47660 , n47661 , n47662 ,
     n47663 , n47664 , n47665 , n47666 , n47667 , n47668 , n47669 , n47670 , n47671 , n47672 ,
     n47673 , n47674 , n47675 , n47676 , n47677 , n47678 , n47679 , n47680 , n47681 , n47682 ,
     n47683 , n47684 , n47685 , n47686 , n47687 , n47688 , n47689 , n47690 , n47691 , n47692 ,
     n47693 , n47694 , n47695 , n47696 , n47697 , n47698 , n47699 , n47700 , n47701 , n47702 ,
     n47703 , n47704 , n47705 , n47706 , n47707 , n47708 , n47709 , n47710 , n47711 , n47712 ,
     n47713 , n47714 , n47715 , n47716 , n47717 , n47718 , n47719 , n47720 , n47721 , n47722 ,
     n47723 , n47724 , n47725 , n47726 , n47727 , n47728 , n47729 , n47730 , n47731 , n47732 ,
     n47733 , n47734 , n47735 , n47736 , n47737 , n47738 , n47739 , n47740 , n47741 , n47742 ,
     n47743 , n47744 , n47745 , n47746 , n47747 , n47748 , n47749 , n47750 , n47751 , n47752 ,
     n47753 , n47754 , n47755 , n47756 , n47757 , n47758 , n47759 , n47760 , n47761 , n47762 ,
     n47763 , n47764 , n47765 , n47766 , n47767 , n47768 , n47769 , n47770 , n47771 , n47772 ,
     n47773 , n47774 , n47775 , n47776 , n47777 , n47778 , n47779 , n47780 , n47781 , n47782 ,
     n47783 , n47784 , n47785 , n47786 , n47787 , n47788 , n47789 , n47790 , n47791 , n47792 ,
     n47793 , n47794 , n47795 , n47796 , n47797 , n47798 , n47799 , n47800 , n47801 , n47802 ,
     n47803 , n47804 , n47805 , n47806 , n47807 , n47808 , n47809 , n47810 , n47811 , n47812 ,
     n47813 , n47814 , n47815 , n47816 , n47817 , n47818 , n47819 , n47820 , n47821 , n47822 ,
     n47823 , n47824 , n47825 , n47826 , n47827 , n47828 , n47829 , n47830 , n47831 , n47832 ,
     n47833 , n47834 , n47835 , n47836 , n47837 , n47838 , n47839 , n47840 , n47841 , n47842 ,
     n47843 , n47844 , n47845 , n47846 , n47847 , n47848 , n47849 , n47850 , n47851 , n47852 ,
     n47853 , n47854 , n47855 , n47856 , n47857 , n47858 , n47859 , n47860 , n47861 , n47862 ,
     n47863 , n47864 , n47865 , n47866 , n47867 , n47868 , n47869 , n47870 , n47871 , n47872 ,
     n47873 , n47874 , n47875 , n47876 , n47877 , n47878 , n47879 , n47880 , n47881 , n47882 ,
     n47883 , n47884 , n47885 , n47886 , n47887 , n47888 , n47889 , n47890 , n47891 , n47892 ,
     n47893 , n47894 , n47895 , n47896 , n47897 , n47898 , n47899 , n47900 , n47901 , n47902 ,
     n47903 , n47904 , n47905 , n47906 , n47907 , n47908 , n47909 , n47910 , n47911 , n47912 ,
     n47913 , n47914 , n47915 , n47916 , n47917 , n47918 , n47919 , n47920 , n47921 , n47922 ,
     n47923 , n47924 , n47925 , n47926 , n47927 , n47928 , n47929 , n47930 , n47931 , n47932 ,
     n47933 , n47934 , n47935 , n47936 , n47937 , n47938 , n47939 , n47940 , n47941 , n47942 ,
     n47943 , n47944 , n47945 , n47946 , n47947 , n47948 , n47949 , n47950 , n47951 , n47952 ,
     n47953 , n47954 , n47955 , n47956 , n47957 , n47958 , n47959 , n47960 , n47961 , n47962 ,
     n47963 , n47964 , n47965 , n47966 , n47967 , n47968 , n47969 , n47970 , n47971 , n47972 ,
     n47973 , n47974 , n47975 , n47976 , n47977 , n47978 , n47979 , n47980 , n47981 , n47982 ,
     n47983 , n47984 , n47985 , n47986 , n47987 , n47988 , n47989 , n47990 , n47991 , n47992 ,
     n47993 , n47994 , n47995 , n47996 , n47997 , n47998 , n47999 , n48000 , n48001 , n48002 ,
     n48003 , n48004 , n48005 , n48006 , n48007 , n48008 , n48009 , n48010 , n48011 , n48012 ,
     n48013 , n48014 , n48015 , n48016 , n48017 , n48018 , n48019 , n48020 , n48021 , n48022 ,
     n48023 , n48024 , n48025 , n48026 , n48027 , n48028 , n48029 , n48030 , n48031 , n48032 ,
     n48033 , n48034 , n48035 , n48036 , n48037 , n48038 , n48039 , n48040 , n48041 , n48042 ,
     n48043 , n48044 , n48045 , n48046 , n48047 , n48048 , n48049 , n48050 , n48051 , n48052 ,
     n48053 , n48054 , n48055 , n48056 , n48057 , n48058 , n48059 , n48060 , n48061 , n48062 ,
     n48063 , n48064 , n48065 , n48066 , n48067 , n48068 , n48069 , n48070 , n48071 , n48072 ,
     n48073 , n48074 , n48075 , n48076 , n48077 , n48078 , n48079 , n48080 , n48081 , n48082 ,
     n48083 , n48084 , n48085 , n48086 , n48087 , n48088 , n48089 , n48090 , n48091 , n48092 ,
     n48093 , n48094 , n48095 , n48096 , n48097 , n48098 , n48099 , n48100 , n48101 , n48102 ,
     n48103 , n48104 , n48105 , n48106 , n48107 , n48108 , n48109 , n48110 , n48111 , n48112 ,
     n48113 , n48114 , n48115 , n48116 , n48117 , n48118 , n48119 , n48120 , n48121 , n48122 ,
     n48123 , n48124 , n48125 , n48126 , n48127 , n48128 , n48129 , n48130 , n48131 , n48132 ,
     n48133 , n48134 , n48135 , n48136 , n48137 , n48138 , n48139 , n48140 , n48141 , n48142 ,
     n48143 , n48144 , n48145 , n48146 , n48147 , n48148 , n48149 , n48150 , n48151 , n48152 ,
     n48153 , n48154 , n48155 , n48156 , n48157 , n48158 , n48159 , n48160 , n48161 , n48162 ,
     n48163 , n48164 , n48165 , n48166 , n48167 , n48168 , n48169 , n48170 , n48171 , n48172 ,
     n48173 , n48174 , n48175 , n48176 , n48177 , n48178 , n48179 , n48180 , n48181 , n48182 ,
     n48183 , n48184 , n48185 , n48186 , n48187 , n48188 , n48189 , n48190 , n48191 , n48192 ,
     n48193 , n48194 , n48195 , n48196 , n48197 , n48198 , n48199 , n48200 , n48201 , n48202 ,
     n48203 , n48204 , n48205 , n48206 , n48207 , n48208 , n48209 , n48210 , n48211 , n48212 ,
     n48213 , n48214 , n48215 , n48216 , n48217 , n48218 , n48219 , n48220 , n48221 , n48222 ,
     n48223 , n48224 , n48225 , n48226 , n48227 , n48228 , n48229 , n48230 , n48231 , n48232 ,
     n48233 , n48234 , n48235 , n48236 , n48237 , n48238 , n48239 , n48240 , n48241 , n48242 ,
     n48243 , n48244 , n48245 , n48246 , n48247 , n48248 , n48249 , n48250 , n48251 , n48252 ,
     n48253 , n48254 , n48255 , n48256 , n48257 , n48258 , n48259 , n48260 , n48261 , n48262 ,
     n48263 , n48264 , n48265 , n48266 , n48267 , n48268 , n48269 , n48270 , n48271 , n48272 ,
     n48273 , n48274 , n48275 , n48276 , n48277 , n48278 , n48279 , n48280 , n48281 , n48282 ,
     n48283 , n48284 , n48285 , n48286 , n48287 , n48288 , n48289 , n48290 , n48291 , n48292 ,
     n48293 , n48294 , n48295 , n48296 , n48297 , n48298 , n48299 , n48300 , n48301 , n48302 ,
     n48303 , n48304 , n48305 , n48306 , n48307 , n48308 , n48309 , n48310 , n48311 , n48312 ,
     n48313 , n48314 , n48315 , n48316 , n48317 , n48318 , n48319 , n48320 , n48321 , n48322 ,
     n48323 , n48324 , n48325 , n48326 , n48327 , n48328 , n48329 , n48330 , n48331 , n48332 ,
     n48333 , n48334 , n48335 , n48336 , n48337 , n48338 , n48339 , n48340 , n48341 , n48342 ,
     n48343 , n48344 , n48345 , n48346 , n48347 , n48348 , n48349 , n48350 , n48351 , n48352 ,
     n48353 , n48354 , n48355 , n48356 , n48357 , n48358 , n48359 , n48360 , n48361 , n48362 ,
     n48363 , n48364 , n48365 , n48366 , n48367 , n48368 , n48369 , n48370 , n48371 , n48372 ,
     n48373 , n48374 , n48375 , n48376 , n48377 , n48378 , n48379 , n48380 , n48381 , n48382 ,
     n48383 , n48384 , n48385 , n48386 , n48387 , n48388 , n48389 , n48390 , n48391 , n48392 ,
     n48393 , n48394 , n48395 , n48396 , n48397 , n48398 , n48399 , n48400 , n48401 , n48402 ,
     n48403 , n48404 , n48405 , n48406 , n48407 , n48408 , n48409 , n48410 , n48411 , n48412 ,
     n48413 , n48414 , n48415 , n48416 , n48417 , n48418 , n48419 , n48420 , n48421 , n48422 ,
     n48423 , n48424 , n48425 , n48426 , n48427 , n48428 , n48429 , n48430 , n48431 , n48432 ,
     n48433 , n48434 , n48435 , n48436 , n48437 , n48438 , n48439 , n48440 , n48441 , n48442 ,
     n48443 , n48444 , n48445 , n48446 , n48447 , n48448 , n48449 , n48450 , n48451 , n48452 ,
     n48453 , n48454 , n48455 , n48456 , n48457 , n48458 , n48459 , n48460 , n48461 , n48462 ,
     n48463 , n48464 , n48465 , n48466 , n48467 , n48468 , n48469 , n48470 , n48471 , n48472 ,
     n48473 , n48474 , n48475 , n48476 , n48477 , n48478 , n48479 , n48480 , n48481 , n48482 ,
     n48483 , n48484 , n48485 , n48486 , n48487 , n48488 , n48489 , n48490 , n48491 , n48492 ,
     n48493 , n48494 , n48495 , n48496 , n48497 , n48498 , n48499 , n48500 , n48501 , n48502 ,
     n48503 , n48504 , n48505 , n48506 , n48507 , n48508 , n48509 , n48510 , n48511 , n48512 ,
     n48513 , n48514 , n48515 , n48516 , n48517 , n48518 , n48519 , n48520 , n48521 , n48522 ,
     n48523 , n48524 , n48525 , n48526 , n48527 , n48528 , n48529 , n48530 , n48531 , n48532 ,
     n48533 , n48534 , n48535 , n48536 , n48537 , n48538 , n48539 , n48540 , n48541 , n48542 ,
     n48543 , n48544 , n48545 , n48546 , n48547 , n48548 , n48549 , n48550 , n48551 , n48552 ,
     n48553 , n48554 , n48555 , n48556 , n48557 , n48558 , n48559 , n48560 , n48561 , n48562 ,
     n48563 , n48564 , n48565 , n48566 , n48567 , n48568 , n48569 , n48570 , n48571 , n48572 ,
     n48573 , n48574 , n48575 , n48576 , n48577 , n48578 , n48579 , n48580 , n48581 , n48582 ,
     n48583 , n48584 , n48585 , n48586 , n48587 , n48588 , n48589 , n48590 , n48591 , n48592 ,
     n48593 , n48594 , n48595 , n48596 , n48597 , n48598 , n48599 , n48600 , n48601 , n48602 ,
     n48603 , n48604 , n48605 , n48606 , n48607 , n48608 , n48609 , n48610 , n48611 , n48612 ,
     n48613 , n48614 , n48615 , n48616 , n48617 , n48618 , n48619 , n48620 , n48621 , n48622 ,
     n48623 , n48624 , n48625 , n48626 , n48627 , n48628 , n48629 , n48630 , n48631 , n48632 ,
     n48633 , n48634 , n48635 , n48636 , n48637 , n48638 , n48639 , n48640 , n48641 , n48642 ,
     n48643 , n48644 , n48645 , n48646 , n48647 , n48648 , n48649 , n48650 , n48651 , n48652 ,
     n48653 , n48654 , n48655 , n48656 , n48657 , n48658 , n48659 , n48660 , n48661 , n48662 ,
     n48663 , n48664 , n48665 , n48666 , n48667 , n48668 , n48669 , n48670 , n48671 , n48672 ,
     n48673 , n48674 , n48675 , n48676 , n48677 , n48678 , n48679 , n48680 , n48681 , n48682 ,
     n48683 , n48684 , n48685 , n48686 , n48687 , n48688 , n48689 , n48690 , n48691 , n48692 ,
     n48693 , n48694 , n48695 , n48696 , n48697 , n48698 , n48699 , n48700 , n48701 , n48702 ,
     n48703 , n48704 , n48705 , n48706 , n48707 , n48708 , n48709 , n48710 , n48711 , n48712 ,
     n48713 , n48714 , n48715 , n48716 , n48717 , n48718 , n48719 , n48720 , n48721 , n48722 ,
     n48723 , n48724 , n48725 , n48726 , n48727 , n48728 , n48729 , n48730 , n48731 , n48732 ,
     n48733 , n48734 , n48735 , n48736 , n48737 , n48738 , n48739 , n48740 , n48741 , n48742 ,
     n48743 , n48744 , n48745 , n48746 , n48747 , n48748 , n48749 , n48750 , n48751 , n48752 ,
     n48753 , n48754 , n48755 , n48756 , n48757 , n48758 , n48759 , n48760 , n48761 , n48762 ,
     n48763 , n48764 , n48765 , n48766 , n48767 , n48768 , n48769 , n48770 , n48771 , n48772 ,
     n48773 , n48774 , n48775 , n48776 , n48777 , n48778 , n48779 , n48780 , n48781 , n48782 ,
     n48783 , n48784 , n48785 , n48786 , n48787 , n48788 , n48789 , n48790 , n48791 , n48792 ,
     n48793 , n48794 , n48795 , n48796 , n48797 , n48798 , n48799 , n48800 , n48801 , n48802 ,
     n48803 , n48804 , n48805 , n48806 , n48807 , n48808 , n48809 , n48810 , n48811 , n48812 ,
     n48813 , n48814 , n48815 , n48816 , n48817 , n48818 , n48819 , n48820 , n48821 , n48822 ,
     n48823 , n48824 , n48825 , n48826 , n48827 , n48828 , n48829 , n48830 , n48831 , n48832 ,
     n48833 , n48834 , n48835 , n48836 , n48837 , n48838 , n48839 , n48840 , n48841 , n48842 ,
     n48843 , n48844 , n48845 , n48846 , n48847 , n48848 , n48849 , n48850 , n48851 , n48852 ,
     n48853 , n48854 , n48855 , n48856 , n48857 , n48858 , n48859 , n48860 , n48861 , n48862 ,
     n48863 , n48864 , n48865 , n48866 , n48867 , n48868 , n48869 , n48870 , n48871 , n48872 ,
     n48873 , n48874 , n48875 , n48876 , n48877 , n48878 , n48879 , n48880 , n48881 , n48882 ,
     n48883 , n48884 , n48885 , n48886 , n48887 , n48888 , n48889 , n48890 , n48891 , n48892 ,
     n48893 , n48894 , n48895 , n48896 , n48897 , n48898 , n48899 , n48900 , n48901 , n48902 ,
     n48903 , n48904 , n48905 , n48906 , n48907 , n48908 , n48909 , n48910 , n48911 , n48912 ,
     n48913 , n48914 , n48915 , n48916 , n48917 , n48918 , n48919 , n48920 , n48921 , n48922 ,
     n48923 , n48924 , n48925 , n48926 , n48927 , n48928 , n48929 , n48930 , n48931 , n48932 ,
     n48933 , n48934 , n48935 , n48936 , n48937 , n48938 , n48939 , n48940 , n48941 , n48942 ,
     n48943 , n48944 , n48945 , n48946 , n48947 , n48948 , n48949 , n48950 , n48951 , n48952 ,
     n48953 , n48954 , n48955 , n48956 , n48957 , n48958 , n48959 , n48960 , n48961 , n48962 ,
     n48963 , n48964 , n48965 , n48966 , n48967 , n48968 , n48969 , n48970 , n48971 , n48972 ,
     n48973 , n48974 , n48975 , n48976 , n48977 , n48978 , n48979 , n48980 , n48981 , n48982 ,
     n48983 , n48984 , n48985 , n48986 , n48987 , n48988 , n48989 , n48990 , n48991 , n48992 ,
     n48993 , n48994 , n48995 , n48996 , n48997 , n48998 , n48999 , n49000 , n49001 , n49002 ,
     n49003 , n49004 , n49005 , n49006 , n49007 , n49008 , n49009 , n49010 , n49011 , n49012 ,
     n49013 , n49014 , n49015 , n49016 , n49017 , n49018 , n49019 , n49020 , n49021 , n49022 ,
     n49023 , n49024 , n49025 , n49026 , n49027 , n49028 , n49029 , n49030 , n49031 , n49032 ,
     n49033 , n49034 , n49035 , n49036 , n49037 , n49038 , n49039 , n49040 , n49041 , n49042 ,
     n49043 , n49044 , n49045 , n49046 , n49047 , n49048 , n49049 , n49050 , n49051 , n49052 ,
     n49053 , n49054 , n49055 , n49056 , n49057 , n49058 , n49059 , n49060 , n49061 , n49062 ,
     n49063 , n49064 , n49065 , n49066 , n49067 , n49068 , n49069 , n49070 , n49071 , n49072 ,
     n49073 , n49074 , n49075 , n49076 , n49077 , n49078 , n49079 , n49080 , n49081 , n49082 ,
     n49083 , n49084 , n49085 , n49086 , n49087 , n49088 , n49089 , n49090 , n49091 , n49092 ,
     n49093 , n49094 , n49095 , n49096 , n49097 , n49098 , n49099 , n49100 , n49101 , n49102 ,
     n49103 , n49104 , n49105 , n49106 , n49107 , n49108 , n49109 , n49110 , n49111 , n49112 ,
     n49113 , n49114 , n49115 , n49116 , n49117 , n49118 , n49119 , n49120 , n49121 , n49122 ,
     n49123 , n49124 , n49125 , n49126 , n49127 , n49128 , n49129 , n49130 , n49131 , n49132 ,
     n49133 , n49134 , n49135 , n49136 , n49137 , n49138 , n49139 , n49140 , n49141 , n49142 ,
     n49143 , n49144 , n49145 , n49146 , n49147 , n49148 , n49149 , n49150 , n49151 , n49152 ,
     n49153 , n49154 , n49155 , n49156 , n49157 , n49158 , n49159 , n49160 , n49161 , n49162 ,
     n49163 , n49164 , n49165 , n49166 , n49167 , n49168 , n49169 , n49170 , n49171 , n49172 ,
     n49173 , n49174 , n49175 , n49176 , n49177 , n49178 , n49179 , n49180 , n49181 , n49182 ,
     n49183 , n49184 , n49185 , n49186 , n49187 , n49188 , n49189 , n49190 , n49191 , n49192 ,
     n49193 , n49194 , n49195 , n49196 , n49197 , n49198 , n49199 , n49200 , n49201 , n49202 ,
     n49203 , n49204 , n49205 , n49206 , n49207 , n49208 , n49209 , n49210 , n49211 , n49212 ,
     n49213 , n49214 , n49215 , n49216 , n49217 , n49218 , n49219 , n49220 , n49221 , n49222 ,
     n49223 , n49224 , n49225 , n49226 , n49227 , n49228 , n49229 , n49230 , n49231 , n49232 ,
     n49233 , n49234 , n49235 , n49236 , n49237 , n49238 , n49239 , n49240 , n49241 , n49242 ,
     n49243 , n49244 , n49245 , n49246 , n49247 , n49248 , n49249 , n49250 , n49251 , n49252 ,
     n49253 , n49254 , n49255 , n49256 , n49257 , n49258 , n49259 , n49260 , n49261 , n49262 ,
     n49263 , n49264 , n49265 , n49266 , n49267 , n49268 , n49269 , n49270 , n49271 , n49272 ,
     n49273 , n49274 , n49275 , n49276 , n49277 , n49278 , n49279 , n49280 , n49281 , n49282 ,
     n49283 , n49284 , n49285 , n49286 , n49287 , n49288 , n49289 , n49290 , n49291 , n49292 ,
     n49293 , n49294 , n49295 , n49296 , n49297 , n49298 , n49299 , n49300 , n49301 , n49302 ,
     n49303 , n49304 , n49305 , n49306 , n49307 , n49308 , n49309 , n49310 , n49311 , n49312 ,
     n49313 , n49314 , n49315 , n49316 , n49317 , n49318 , n49319 , n49320 , n49321 , n49322 ,
     n49323 , n49324 , n49325 , n49326 , n49327 , n49328 , n49329 , n49330 , n49331 , n49332 ,
     n49333 , n49334 , n49335 , n49336 , n49337 , n49338 , n49339 , n49340 , n49341 , n49342 ,
     n49343 , n49344 , n49345 , n49346 , n49347 , n49348 , n49349 , n49350 , n49351 , n49352 ,
     n49353 , n49354 , n49355 , n49356 , n49357 , n49358 , n49359 , n49360 , n49361 , n49362 ,
     n49363 , n49364 , n49365 , n49366 , n49367 , n49368 , n49369 , n49370 , n49371 , n49372 ,
     n49373 , n49374 , n49375 , n49376 , n49377 , n49378 , n49379 , n49380 , n49381 , n49382 ,
     n49383 , n49384 , n49385 , n49386 , n49387 , n49388 , n49389 , n49390 , n49391 , n49392 ,
     n49393 , n49394 , n49395 , n49396 , n49397 , n49398 , n49399 , n49400 , n49401 , n49402 ,
     n49403 , n49404 , n49405 , n49406 , n49407 , n49408 , n49409 , n49410 , n49411 , n49412 ,
     n49413 , n49414 , n49415 , n49416 , n49417 , n49418 , n49419 , n49420 , n49421 , n49422 ,
     n49423 , n49424 , n49425 , n49426 , n49427 , n49428 , n49429 , n49430 , n49431 , n49432 ,
     n49433 , n49434 , n49435 , n49436 , n49437 , n49438 , n49439 , n49440 , n49441 , n49442 ,
     n49443 , n49444 , n49445 , n49446 , n49447 , n49448 , n49449 , n49450 , n49451 , n49452 ,
     n49453 , n49454 , n49455 , n49456 , n49457 , n49458 , n49459 , n49460 , n49461 , n49462 ,
     n49463 , n49464 , n49465 , n49466 , n49467 , n49468 , n49469 , n49470 , n49471 , n49472 ,
     n49473 , n49474 , n49475 , n49476 , n49477 , n49478 , n49479 , n49480 , n49481 , n49482 ,
     n49483 , n49484 , n49485 , n49486 , n49487 , n49488 , n49489 , n49490 , n49491 , n49492 ,
     n49493 , n49494 , n49495 , n49496 , n49497 , n49498 , n49499 , n49500 , n49501 , n49502 ,
     n49503 , n49504 , n49505 , n49506 , n49507 , n49508 , n49509 , n49510 , n49511 , n49512 ,
     n49513 , n49514 , n49515 , n49516 , n49517 , n49518 , n49519 , n49520 , n49521 , n49522 ,
     n49523 , n49524 , n49525 , n49526 , n49527 , n49528 , n49529 , n49530 , n49531 , n49532 ,
     n49533 , n49534 , n49535 , n49536 , n49537 , n49538 , n49539 , n49540 , n49541 , n49542 ,
     n49543 , n49544 , n49545 , n49546 , n49547 , n49548 , n49549 , n49550 , n49551 , n49552 ,
     n49553 , n49554 , n49555 , n49556 , n49557 , n49558 , n49559 , n49560 , n49561 , n49562 ,
     n49563 , n49564 , n49565 , n49566 , n49567 , n49568 , n49569 , n49570 , n49571 , n49572 ,
     n49573 , n49574 , n49575 , n49576 , n49577 , n49578 , n49579 , n49580 , n49581 , n49582 ,
     n49583 , n49584 , n49585 , n49586 , n49587 , n49588 , n49589 , n49590 , n49591 , n49592 ,
     n49593 , n49594 , n49595 , n49596 , n49597 , n49598 , n49599 , n49600 , n49601 , n49602 ,
     n49603 , n49604 , n49605 , n49606 , n49607 , n49608 , n49609 , n49610 , n49611 , n49612 ,
     n49613 , n49614 , n49615 , n49616 , n49617 , n49618 , n49619 , n49620 , n49621 , n49622 ,
     n49623 , n49624 , n49625 , n49626 , n49627 , n49628 , n49629 , n49630 , n49631 , n49632 ,
     n49633 , n49634 , n49635 , n49636 , n49637 , n49638 , n49639 , n49640 , n49641 , n49642 ,
     n49643 , n49644 , n49645 , n49646 , n49647 , n49648 , n49649 , n49650 , n49651 , n49652 ,
     n49653 , n49654 , n49655 , n49656 , n49657 , n49658 , n49659 , n49660 , n49661 , n49662 ,
     n49663 , n49664 , n49665 , n49666 , n49667 , n49668 , n49669 , n49670 , n49671 , n49672 ,
     n49673 , n49674 , n49675 , n49676 , n49677 , n49678 , n49679 , n49680 , n49681 , n49682 ,
     n49683 , n49684 , n49685 , n49686 , n49687 , n49688 , n49689 , n49690 , n49691 , n49692 ,
     n49693 , n49694 , n49695 , n49696 , n49697 , n49698 , n49699 , n49700 , n49701 , n49702 ,
     n49703 , n49704 , n49705 , n49706 , n49707 , n49708 , n49709 , n49710 , n49711 , n49712 ,
     n49713 , n49714 , n49715 , n49716 , n49717 , n49718 , n49719 , n49720 , n49721 , n49722 ,
     n49723 , n49724 , n49725 , n49726 , n49727 , n49728 , n49729 , n49730 , n49731 , n49732 ,
     n49733 , n49734 , n49735 , n49736 , n49737 , n49738 , n49739 , n49740 , n49741 , n49742 ,
     n49743 , n49744 , n49745 , n49746 , n49747 , n49748 , n49749 , n49750 , n49751 , n49752 ,
     n49753 , n49754 , n49755 , n49756 , n49757 , n49758 , n49759 , n49760 , n49761 , n49762 ,
     n49763 , n49764 , n49765 , n49766 , n49767 , n49768 , n49769 , n49770 , n49771 , n49772 ,
     n49773 , n49774 , n49775 , n49776 , n49777 , n49778 , n49779 , n49780 , n49781 , n49782 ,
     n49783 , n49784 , n49785 , n49786 , n49787 , n49788 , n49789 , n49790 , n49791 , n49792 ,
     n49793 , n49794 , n49795 , n49796 , n49797 , n49798 , n49799 , n49800 , n49801 , n49802 ,
     n49803 , n49804 , n49805 , n49806 , n49807 , n49808 , n49809 , n49810 , n49811 , n49812 ,
     n49813 , n49814 , n49815 , n49816 , n49817 , n49818 , n49819 , n49820 , n49821 , n49822 ,
     n49823 , n49824 , n49825 , n49826 , n49827 , n49828 , n49829 , n49830 , n49831 , n49832 ,
     n49833 , n49834 , n49835 , n49836 , n49837 , n49838 , n49839 , n49840 , n49841 , n49842 ,
     n49843 , n49844 , n49845 , n49846 , n49847 , n49848 , n49849 , n49850 , n49851 , n49852 ,
     n49853 , n49854 , n49855 , n49856 , n49857 , n49858 , n49859 , n49860 , n49861 , n49862 ,
     n49863 , n49864 , n49865 , n49866 , n49867 , n49868 , n49869 , n49870 , n49871 , n49872 ,
     n49873 , n49874 , n49875 , n49876 , n49877 , n49878 , n49879 , n49880 , n49881 , n49882 ,
     n49883 , n49884 , n49885 , n49886 , n49887 , n49888 , n49889 , n49890 , n49891 , n49892 ,
     n49893 , n49894 , n49895 , n49896 , n49897 , n49898 , n49899 , n49900 , n49901 , n49902 ,
     n49903 , n49904 , n49905 , n49906 , n49907 , n49908 , n49909 , n49910 , n49911 , n49912 ,
     n49913 , n49914 , n49915 , n49916 , n49917 , n49918 , n49919 , n49920 , n49921 , n49922 ,
     n49923 , n49924 , n49925 , n49926 , n49927 , n49928 , n49929 , n49930 , n49931 , n49932 ,
     n49933 , n49934 , n49935 , n49936 , n49937 , n49938 , n49939 , n49940 , n49941 , n49942 ,
     n49943 , n49944 , n49945 , n49946 , n49947 , n49948 , n49949 , n49950 , n49951 , n49952 ,
     n49953 , n49954 , n49955 , n49956 , n49957 , n49958 , n49959 , n49960 , n49961 , n49962 ,
     n49963 , n49964 , n49965 , n49966 , n49967 , n49968 , n49969 , n49970 , n49971 , n49972 ,
     n49973 , n49974 , n49975 , n49976 , n49977 , n49978 , n49979 , n49980 , n49981 , n49982 ,
     n49983 , n49984 , n49985 , n49986 , n49987 , n49988 , n49989 , n49990 , n49991 , n49992 ,
     n49993 , n49994 , n49995 , n49996 , n49997 , n49998 , n49999 , n50000 , n50001 , n50002 ,
     n50003 , n50004 , n50005 , n50006 , n50007 , n50008 , n50009 , n50010 , n50011 , n50012 ,
     n50013 , n50014 , n50015 , n50016 , n50017 , n50018 , n50019 , n50020 , n50021 , n50022 ,
     n50023 , n50024 , n50025 , n50026 , n50027 , n50028 , n50029 , n50030 , n50031 , n50032 ,
     n50033 , n50034 , n50035 , n50036 , n50037 , n50038 , n50039 , n50040 , n50041 , n50042 ,
     n50043 , n50044 , n50045 , n50046 , n50047 , n50048 , n50049 , n50050 , n50051 , n50052 ,
     n50053 , n50054 , n50055 , n50056 , n50057 , n50058 , n50059 , n50060 , n50061 , n50062 ,
     n50063 , n50064 , n50065 , n50066 , n50067 , n50068 , n50069 , n50070 , n50071 , n50072 ,
     n50073 , n50074 , n50075 , n50076 , n50077 , n50078 , n50079 , n50080 , n50081 , n50082 ,
     n50083 , n50084 , n50085 , n50086 , n50087 , n50088 , n50089 , n50090 , n50091 , n50092 ,
     n50093 , n50094 , n50095 , n50096 , n50097 , n50098 , n50099 , n50100 , n50101 , n50102 ,
     n50103 , n50104 , n50105 , n50106 , n50107 , n50108 , n50109 , n50110 , n50111 , n50112 ,
     n50113 , n50114 , n50115 , n50116 , n50117 , n50118 , n50119 , n50120 , n50121 , n50122 ,
     n50123 , n50124 , n50125 , n50126 , n50127 , n50128 , n50129 , n50130 , n50131 , n50132 ,
     n50133 , n50134 , n50135 , n50136 , n50137 , n50138 , n50139 , n50140 , n50141 , n50142 ,
     n50143 , n50144 , n50145 , n50146 , n50147 , n50148 , n50149 , n50150 , n50151 , n50152 ,
     n50153 , n50154 , n50155 , n50156 , n50157 , n50158 , n50159 , n50160 , n50161 , n50162 ,
     n50163 , n50164 , n50165 , n50166 , n50167 , n50168 , n50169 , n50170 , n50171 , n50172 ,
     n50173 , n50174 , n50175 , n50176 , n50177 , n50178 , n50179 , n50180 , n50181 , n50182 ,
     n50183 , n50184 , n50185 , n50186 , n50187 , n50188 , n50189 , n50190 , n50191 , n50192 ,
     n50193 , n50194 , n50195 , n50196 , n50197 , n50198 , n50199 , n50200 , n50201 , n50202 ,
     n50203 , n50204 , n50205 , n50206 , n50207 , n50208 , n50209 , n50210 , n50211 , n50212 ,
     n50213 , n50214 , n50215 , n50216 , n50217 , n50218 , n50219 , n50220 , n50221 , n50222 ,
     n50223 , n50224 , n50225 , n50226 , n50227 , n50228 , n50229 , n50230 , n50231 , n50232 ,
     n50233 , n50234 , n50235 , n50236 , n50237 , n50238 , n50239 , n50240 , n50241 , n50242 ,
     n50243 , n50244 , n50245 , n50246 , n50247 , n50248 , n50249 , n50250 , n50251 , n50252 ,
     n50253 , n50254 , n50255 , n50256 , n50257 , n50258 , n50259 , n50260 , n50261 , n50262 ,
     n50263 , n50264 , n50265 , n50266 , n50267 , n50268 , n50269 , n50270 , n50271 , n50272 ,
     n50273 , n50274 , n50275 , n50276 , n50277 , n50278 , n50279 , n50280 , n50281 , n50282 ,
     n50283 , n50284 , n50285 , n50286 , n50287 , n50288 , n50289 , n50290 , n50291 , n50292 ,
     n50293 , n50294 , n50295 , n50296 , n50297 , n50298 , n50299 , n50300 , n50301 , n50302 ,
     n50303 , n50304 , n50305 , n50306 , n50307 , n50308 , n50309 , n50310 , n50311 , n50312 ,
     n50313 , n50314 , n50315 , n50316 , n50317 , n50318 , n50319 , n50320 , n50321 , n50322 ,
     n50323 , n50324 , n50325 , n50326 , n50327 , n50328 , n50329 , n50330 , n50331 , n50332 ,
     n50333 , n50334 , n50335 , n50336 , n50337 , n50338 , n50339 , n50340 , n50341 , n50342 ,
     n50343 , n50344 , n50345 , n50346 , n50347 , n50348 , n50349 , n50350 , n50351 , n50352 ,
     n50353 , n50354 , n50355 , n50356 , n50357 , n50358 , n50359 , n50360 , n50361 , n50362 ,
     n50363 , n50364 , n50365 , n50366 , n50367 , n50368 , n50369 , n50370 , n50371 , n50372 ,
     n50373 , n50374 , n50375 , n50376 , n50377 , n50378 , n50379 , n50380 , n50381 , n50382 ,
     n50383 , n50384 , n50385 , n50386 , n50387 , n50388 , n50389 , n50390 , n50391 , n50392 ,
     n50393 , n50394 , n50395 , n50396 , n50397 , n50398 , n50399 , n50400 , n50401 , n50402 ,
     n50403 , n50404 , n50405 , n50406 , n50407 , n50408 , n50409 , n50410 , n50411 , n50412 ,
     n50413 , n50414 , n50415 , n50416 , n50417 , n50418 , n50419 , n50420 , n50421 , n50422 ,
     n50423 , n50424 , n50425 , n50426 , n50427 , n50428 , n50429 , n50430 , n50431 , n50432 ,
     n50433 , n50434 , n50435 , n50436 , n50437 , n50438 , n50439 , n50440 , n50441 , n50442 ,
     n50443 , n50444 , n50445 , n50446 , n50447 , n50448 , n50449 , n50450 , n50451 , n50452 ,
     n50453 , n50454 , n50455 , n50456 , n50457 , n50458 , n50459 , n50460 , n50461 , n50462 ,
     n50463 , n50464 , n50465 , n50466 , n50467 , n50468 , n50469 , n50470 , n50471 , n50472 ,
     n50473 , n50474 , n50475 , n50476 , n50477 , n50478 , n50479 , n50480 , n50481 , n50482 ,
     n50483 , n50484 , n50485 , n50486 , n50487 , n50488 , n50489 , n50490 , n50491 , n50492 ,
     n50493 , n50494 , n50495 , n50496 , n50497 , n50498 , n50499 , n50500 , n50501 , n50502 ,
     n50503 , n50504 , n50505 , n50506 , n50507 , n50508 , n50509 , n50510 , n50511 , n50512 ,
     n50513 , n50514 , n50515 , n50516 , n50517 , n50518 , n50519 , n50520 , n50521 , n50522 ,
     n50523 , n50524 , n50525 , n50526 , n50527 , n50528 , n50529 , n50530 , n50531 , n50532 ,
     n50533 , n50534 , n50535 , n50536 , n50537 , n50538 , n50539 , n50540 , n50541 , n50542 ,
     n50543 , n50544 , n50545 , n50546 , n50547 , n50548 , n50549 , n50550 , n50551 , n50552 ,
     n50553 , n50554 , n50555 , n50556 , n50557 , n50558 , n50559 , n50560 , n50561 , n50562 ,
     n50563 , n50564 , n50565 , n50566 , n50567 , n50568 , n50569 , n50570 , n50571 , n50572 ,
     n50573 , n50574 , n50575 , n50576 , n50577 , n50578 , n50579 , n50580 , n50581 , n50582 ,
     n50583 , n50584 , n50585 , n50586 , n50587 , n50588 , n50589 , n50590 , n50591 , n50592 ,
     n50593 , n50594 , n50595 , n50596 , n50597 , n50598 , n50599 , n50600 , n50601 , n50602 ,
     n50603 , n50604 , n50605 , n50606 , n50607 , n50608 , n50609 , n50610 , n50611 , n50612 ,
     n50613 , n50614 , n50615 , n50616 , n50617 , n50618 , n50619 , n50620 , n50621 , n50622 ,
     n50623 , n50624 , n50625 , n50626 , n50627 , n50628 , n50629 , n50630 , n50631 , n50632 ,
     n50633 , n50634 , n50635 , n50636 , n50637 , n50638 , n50639 , n50640 , n50641 , n50642 ,
     n50643 , n50644 , n50645 , n50646 , n50647 , n50648 , n50649 , n50650 , n50651 , n50652 ,
     n50653 , n50654 , n50655 , n50656 , n50657 , n50658 , n50659 , n50660 , n50661 , n50662 ,
     n50663 , n50664 , n50665 , n50666 , n50667 , n50668 , n50669 , n50670 , n50671 , n50672 ,
     n50673 , n50674 , n50675 , n50676 , n50677 , n50678 , n50679 , n50680 , n50681 , n50682 ,
     n50683 , n50684 , n50685 , n50686 , n50687 , n50688 , n50689 , n50690 , n50691 , n50692 ,
     n50693 , n50694 , n50695 , n50696 , n50697 , n50698 , n50699 , n50700 , n50701 , n50702 ,
     n50703 , n50704 , n50705 , n50706 , n50707 , n50708 , n50709 , n50710 , n50711 , n50712 ,
     n50713 , n50714 , n50715 , n50716 , n50717 , n50718 , n50719 , n50720 , n50721 , n50722 ,
     n50723 , n50724 , n50725 , n50726 , n50727 , n50728 , n50729 , n50730 , n50731 , n50732 ,
     n50733 , n50734 , n50735 , n50736 , n50737 , n50738 , n50739 , n50740 , n50741 , n50742 ,
     n50743 , n50744 , n50745 , n50746 , n50747 , n50748 , n50749 , n50750 , n50751 , n50752 ,
     n50753 , n50754 , n50755 , n50756 , n50757 , n50758 , n50759 , n50760 , n50761 , n50762 ,
     n50763 , n50764 , n50765 , n50766 , n50767 , n50768 , n50769 , n50770 , n50771 , n50772 ,
     n50773 , n50774 , n50775 , n50776 , n50777 , n50778 , n50779 , n50780 , n50781 , n50782 ,
     n50783 , n50784 , n50785 , n50786 , n50787 , n50788 , n50789 , n50790 , n50791 , n50792 ,
     n50793 , n50794 , n50795 , n50796 , n50797 , n50798 , n50799 , n50800 , n50801 , n50802 ,
     n50803 , n50804 , n50805 , n50806 , n50807 , n50808 , n50809 , n50810 , n50811 , n50812 ,
     n50813 , n50814 , n50815 , n50816 , n50817 , n50818 , n50819 , n50820 , n50821 , n50822 ,
     n50823 , n50824 , n50825 , n50826 , n50827 , n50828 , n50829 , n50830 , n50831 , n50832 ,
     n50833 , n50834 , n50835 , n50836 , n50837 , n50838 , n50839 , n50840 , n50841 , n50842 ,
     n50843 , n50844 , n50845 , n50846 , n50847 , n50848 , n50849 , n50850 , n50851 , n50852 ,
     n50853 , n50854 , n50855 , n50856 , n50857 , n50858 , n50859 , n50860 , n50861 , n50862 ,
     n50863 , n50864 , n50865 , n50866 , n50867 , n50868 , n50869 , n50870 , n50871 , n50872 ,
     n50873 , n50874 , n50875 , n50876 , n50877 , n50878 , n50879 , n50880 , n50881 , n50882 ,
     n50883 , n50884 , n50885 , n50886 , n50887 , n50888 , n50889 , n50890 , n50891 , n50892 ,
     n50893 , n50894 , n50895 , n50896 , n50897 , n50898 , n50899 , n50900 , n50901 , n50902 ,
     n50903 , n50904 , n50905 , n50906 , n50907 , n50908 , n50909 , n50910 , n50911 , n50912 ,
     n50913 , n50914 , n50915 , n50916 , n50917 , n50918 , n50919 , n50920 , n50921 , n50922 ,
     n50923 , n50924 , n50925 , n50926 , n50927 , n50928 , n50929 , n50930 , n50931 , n50932 ,
     n50933 , n50934 , n50935 , n50936 , n50937 , n50938 , n50939 , n50940 , n50941 , n50942 ,
     n50943 , n50944 , n50945 , n50946 , n50947 , n50948 , n50949 , n50950 , n50951 , n50952 ,
     n50953 , n50954 , n50955 , n50956 , n50957 , n50958 , n50959 , n50960 , n50961 , n50962 ,
     n50963 , n50964 , n50965 , n50966 , n50967 , n50968 , n50969 , n50970 , n50971 , n50972 ,
     n50973 , n50974 , n50975 , n50976 , n50977 , n50978 , n50979 , n50980 , n50981 , n50982 ,
     n50983 , n50984 , n50985 , n50986 , n50987 , n50988 , n50989 , n50990 , n50991 , n50992 ,
     n50993 , n50994 , n50995 , n50996 , n50997 , n50998 , n50999 , n51000 , n51001 , n51002 ,
     n51003 , n51004 , n51005 , n51006 , n51007 , n51008 , n51009 , n51010 , n51011 , n51012 ,
     n51013 , n51014 , n51015 , n51016 , n51017 , n51018 , n51019 , n51020 , n51021 , n51022 ,
     n51023 , n51024 , n51025 , n51026 , n51027 , n51028 , n51029 , n51030 , n51031 , n51032 ,
     n51033 , n51034 , n51035 , n51036 , n51037 , n51038 , n51039 , n51040 , n51041 , n51042 ,
     n51043 , n51044 , n51045 , n51046 , n51047 , n51048 , n51049 , n51050 , n51051 , n51052 ,
     n51053 , n51054 , n51055 , n51056 , n51057 , n51058 , n51059 , n51060 , n51061 , n51062 ,
     n51063 , n51064 , n51065 , n51066 , n51067 , n51068 , n51069 , n51070 , n51071 , n51072 ,
     n51073 , n51074 , n51075 , n51076 , n51077 , n51078 , n51079 , n51080 , n51081 , n51082 ,
     n51083 , n51084 , n51085 , n51086 , n51087 , n51088 , n51089 , n51090 , n51091 , n51092 ,
     n51093 , n51094 , n51095 , n51096 , n51097 , n51098 , n51099 , n51100 , n51101 , n51102 ,
     n51103 , n51104 , n51105 , n51106 , n51107 , n51108 , n51109 , n51110 , n51111 , n51112 ,
     n51113 , n51114 , n51115 , n51116 , n51117 , n51118 , n51119 , n51120 , n51121 , n51122 ,
     n51123 , n51124 , n51125 , n51126 , n51127 , n51128 , n51129 , n51130 , n51131 , n51132 ,
     n51133 , n51134 , n51135 , n51136 , n51137 , n51138 , n51139 , n51140 , n51141 , n51142 ,
     n51143 , n51144 , n51145 , n51146 , n51147 , n51148 , n51149 , n51150 , n51151 , n51152 ,
     n51153 , n51154 , n51155 , n51156 , n51157 , n51158 , n51159 , n51160 , n51161 , n51162 ,
     n51163 , n51164 , n51165 , n51166 , n51167 , n51168 , n51169 , n51170 , n51171 , n51172 ,
     n51173 , n51174 , n51175 , n51176 , n51177 , n51178 , n51179 , n51180 , n51181 , n51182 ,
     n51183 , n51184 , n51185 , n51186 , n51187 , n51188 , n51189 , n51190 , n51191 , n51192 ,
     n51193 , n51194 , n51195 , n51196 , n51197 , n51198 , n51199 , n51200 , n51201 , n51202 ,
     n51203 , n51204 , n51205 , n51206 , n51207 , n51208 , n51209 , n51210 , n51211 , n51212 ,
     n51213 , n51214 , n51215 , n51216 , n51217 , n51218 , n51219 , n51220 , n51221 , n51222 ,
     n51223 , n51224 , n51225 , n51226 , n51227 , n51228 , n51229 , n51230 , n51231 , n51232 ,
     n51233 , n51234 , n51235 , n51236 , n51237 , n51238 , n51239 , n51240 , n51241 , n51242 ,
     n51243 , n51244 , n51245 , n51246 , n51247 , n51248 , n51249 , n51250 , n51251 , n51252 ,
     n51253 , n51254 , n51255 , n51256 , n51257 , n51258 , n51259 , n51260 , n51261 , n51262 ,
     n51263 , n51264 , n51265 , n51266 , n51267 , n51268 , n51269 , n51270 , n51271 , n51272 ,
     n51273 , n51274 , n51275 , n51276 , n51277 , n51278 , n51279 , n51280 , n51281 , n51282 ,
     n51283 , n51284 , n51285 , n51286 , n51287 , n51288 , n51289 , n51290 , n51291 , n51292 ,
     n51293 , n51294 , n51295 , n51296 , n51297 , n51298 , n51299 , n51300 , n51301 , n51302 ,
     n51303 , n51304 , n51305 , n51306 , n51307 , n51308 , n51309 , n51310 , n51311 , n51312 ,
     n51313 , n51314 , n51315 , n51316 , n51317 , n51318 , n51319 , n51320 , n51321 , n51322 ,
     n51323 , n51324 , n51325 , n51326 , n51327 , n51328 , n51329 , n51330 , n51331 , n51332 ,
     n51333 , n51334 , n51335 , n51336 , n51337 , n51338 , n51339 , n51340 , n51341 , n51342 ,
     n51343 , n51344 , n51345 , n51346 , n51347 , n51348 , n51349 , n51350 , n51351 , n51352 ,
     n51353 , n51354 , n51355 , n51356 , n51357 , n51358 , n51359 , n51360 , n51361 , n51362 ,
     n51363 , n51364 , n51365 , n51366 , n51367 , n51368 , n51369 , n51370 , n51371 , n51372 ,
     n51373 , n51374 , n51375 , n51376 , n51377 , n51378 , n51379 , n51380 , n51381 , n51382 ,
     n51383 , n51384 , n51385 , n51386 , n51387 , n51388 , n51389 , n51390 , n51391 , n51392 ,
     n51393 , n51394 , n51395 , n51396 , n51397 , n51398 , n51399 , n51400 , n51401 , n51402 ,
     n51403 , n51404 , n51405 , n51406 , n51407 , n51408 , n51409 , n51410 , n51411 , n51412 ,
     n51413 , n51414 , n51415 , n51416 , n51417 , n51418 , n51419 , n51420 , n51421 , n51422 ,
     n51423 , n51424 , n51425 , n51426 , n51427 , n51428 , n51429 , n51430 , n51431 , n51432 ,
     n51433 , n51434 , n51435 , n51436 , n51437 , n51438 , n51439 , n51440 , n51441 , n51442 ,
     n51443 , n51444 , n51445 , n51446 , n51447 , n51448 , n51449 , n51450 , n51451 , n51452 ,
     n51453 , n51454 , n51455 , n51456 , n51457 , n51458 , n51459 , n51460 , n51461 , n51462 ,
     n51463 , n51464 , n51465 , n51466 , n51467 , n51468 , n51469 , n51470 , n51471 , n51472 ,
     n51473 , n51474 , n51475 , n51476 , n51477 , n51478 , n51479 , n51480 , n51481 , n51482 ,
     n51483 , n51484 , n51485 , n51486 , n51487 , n51488 , n51489 , n51490 , n51491 , n51492 ,
     n51493 , n51494 , n51495 , n51496 , n51497 , n51498 , n51499 , n51500 , n51501 , n51502 ,
     n51503 , n51504 , n51505 , n51506 , n51507 , n51508 , n51509 , n51510 , n51511 , n51512 ,
     n51513 , n51514 , n51515 , n51516 , n51517 , n51518 , n51519 , n51520 , n51521 , n51522 ,
     n51523 , n51524 , n51525 , n51526 , n51527 , n51528 , n51529 , n51530 , n51531 , n51532 ,
     n51533 , n51534 , n51535 , n51536 , n51537 , n51538 , n51539 , n51540 , n51541 , n51542 ,
     n51543 , n51544 , n51545 , n51546 , n51547 , n51548 , n51549 , n51550 , n51551 , n51552 ,
     n51553 , n51554 , n51555 , n51556 , n51557 , n51558 , n51559 , n51560 , n51561 , n51562 ,
     n51563 , n51564 , n51565 , n51566 , n51567 , n51568 , n51569 , n51570 , n51571 , n51572 ,
     n51573 , n51574 , n51575 , n51576 , n51577 , n51578 , n51579 , n51580 , n51581 , n51582 ,
     n51583 , n51584 , n51585 , n51586 , n51587 , n51588 , n51589 , n51590 , n51591 , n51592 ,
     n51593 , n51594 , n51595 , n51596 , n51597 , n51598 , n51599 , n51600 , n51601 , n51602 ,
     n51603 , n51604 , n51605 , n51606 , n51607 , n51608 , n51609 , n51610 , n51611 , n51612 ,
     n51613 , n51614 , n51615 , n51616 , n51617 , n51618 , n51619 , n51620 , n51621 , n51622 ,
     n51623 , n51624 , n51625 , n51626 , n51627 , n51628 , n51629 , n51630 , n51631 , n51632 ,
     n51633 , n51634 , n51635 , n51636 , n51637 , n51638 , n51639 , n51640 , n51641 , n51642 ,
     n51643 , n51644 , n51645 , n51646 , n51647 , n51648 , n51649 , n51650 , n51651 , n51652 ,
     n51653 , n51654 , n51655 , n51656 , n51657 , n51658 , n51659 , n51660 , n51661 , n51662 ,
     n51663 , n51664 , n51665 , n51666 , n51667 , n51668 , n51669 , n51670 , n51671 , n51672 ,
     n51673 , n51674 , n51675 , n51676 , n51677 , n51678 , n51679 , n51680 , n51681 , n51682 ,
     n51683 , n51684 , n51685 , n51686 , n51687 , n51688 , n51689 , n51690 , n51691 , n51692 ,
     n51693 , n51694 , n51695 , n51696 , n51697 , n51698 , n51699 , n51700 , n51701 , n51702 ,
     n51703 , n51704 , n51705 , n51706 , n51707 , n51708 , n51709 , n51710 , n51711 , n51712 ,
     n51713 , n51714 , n51715 , n51716 , n51717 , n51718 , n51719 , n51720 , n51721 , n51722 ,
     n51723 , n51724 , n51725 , n51726 , n51727 , n51728 , n51729 , n51730 , n51731 , n51732 ,
     n51733 , n51734 , n51735 , n51736 , n51737 , n51738 , n51739 , n51740 , n51741 , n51742 ,
     n51743 , n51744 , n51745 , n51746 , n51747 , n51748 , n51749 , n51750 , n51751 , n51752 ,
     n51753 , n51754 , n51755 , n51756 , n51757 , n51758 , n51759 , n51760 , n51761 , n51762 ,
     n51763 , n51764 , n51765 , n51766 , n51767 , n51768 , n51769 , n51770 , n51771 , n51772 ,
     n51773 , n51774 , n51775 , n51776 , n51777 , n51778 , n51779 , n51780 , n51781 , n51782 ,
     n51783 , n51784 , n51785 , n51786 , n51787 , n51788 , n51789 , n51790 , n51791 , n51792 ,
     n51793 , n51794 , n51795 , n51796 , n51797 , n51798 , n51799 , n51800 , n51801 , n51802 ,
     n51803 , n51804 , n51805 , n51806 , n51807 , n51808 , n51809 , n51810 , n51811 , n51812 ,
     n51813 , n51814 , n51815 , n51816 , n51817 , n51818 , n51819 , n51820 , n51821 , n51822 ,
     n51823 , n51824 , n51825 , n51826 , n51827 , n51828 , n51829 , n51830 , n51831 , n51832 ,
     n51833 , n51834 , n51835 , n51836 , n51837 , n51838 , n51839 , n51840 , n51841 , n51842 ,
     n51843 , n51844 , n51845 , n51846 , n51847 , n51848 , n51849 , n51850 , n51851 , n51852 ,
     n51853 , n51854 , n51855 , n51856 , n51857 , n51858 , n51859 , n51860 , n51861 , n51862 ,
     n51863 , n51864 , n51865 , n51866 , n51867 , n51868 , n51869 , n51870 , n51871 , n51872 ,
     n51873 , n51874 , n51875 , n51876 , n51877 , n51878 , n51879 , n51880 , n51881 , n51882 ,
     n51883 , n51884 , n51885 , n51886 , n51887 , n51888 , n51889 , n51890 , n51891 , n51892 ,
     n51893 , n51894 , n51895 , n51896 , n51897 , n51898 , n51899 , n51900 , n51901 , n51902 ,
     n51903 , n51904 , n51905 , n51906 , n51907 , n51908 , n51909 , n51910 , n51911 , n51912 ,
     n51913 , n51914 , n51915 , n51916 , n51917 , n51918 , n51919 , n51920 , n51921 , n51922 ,
     n51923 , n51924 , n51925 , n51926 , n51927 , n51928 , n51929 , n51930 , n51931 , n51932 ,
     n51933 , n51934 , n51935 , n51936 , n51937 , n51938 , n51939 , n51940 , n51941 , n51942 ,
     n51943 , n51944 , n51945 , n51946 , n51947 , n51948 , n51949 , n51950 , n51951 , n51952 ,
     n51953 , n51954 , n51955 , n51956 , n51957 , n51958 , n51959 , n51960 , n51961 , n51962 ,
     n51963 , n51964 , n51965 , n51966 , n51967 , n51968 , n51969 , n51970 , n51971 , n51972 ,
     n51973 , n51974 , n51975 , n51976 , n51977 , n51978 , n51979 , n51980 , n51981 , n51982 ,
     n51983 , n51984 , n51985 , n51986 , n51987 , n51988 , n51989 , n51990 , n51991 , n51992 ,
     n51993 , n51994 , n51995 , n51996 , n51997 , n51998 , n51999 , n52000 , n52001 , n52002 ,
     n52003 , n52004 , n52005 , n52006 , n52007 , n52008 , n52009 , n52010 , n52011 , n52012 ,
     n52013 , n52014 , n52015 , n52016 , n52017 , n52018 , n52019 , n52020 , n52021 , n52022 ,
     n52023 , n52024 , n52025 , n52026 , n52027 , n52028 , n52029 , n52030 , n52031 , n52032 ,
     n52033 , n52034 , n52035 , n52036 , n52037 , n52038 , n52039 , n52040 , n52041 , n52042 ,
     n52043 , n52044 , n52045 , n52046 , n52047 , n52048 , n52049 , n52050 , n52051 , n52052 ,
     n52053 , n52054 , n52055 , n52056 , n52057 , n52058 , n52059 , n52060 , n52061 , n52062 ,
     n52063 , n52064 , n52065 , n52066 , n52067 , n52068 , n52069 , n52070 , n52071 , n52072 ,
     n52073 , n52074 , n52075 , n52076 , n52077 , n52078 , n52079 , n52080 , n52081 , n52082 ,
     n52083 , n52084 , n52085 , n52086 , n52087 , n52088 , n52089 , n52090 , n52091 , n52092 ,
     n52093 , n52094 , n52095 , n52096 , n52097 , n52098 , n52099 , n52100 , n52101 , n52102 ,
     n52103 , n52104 , n52105 , n52106 , n52107 , n52108 , n52109 , n52110 , n52111 , n52112 ,
     n52113 , n52114 , n52115 , n52116 , n52117 , n52118 , n52119 , n52120 , n52121 , n52122 ,
     n52123 , n52124 , n52125 , n52126 , n52127 , n52128 , n52129 , n52130 , n52131 , n52132 ,
     n52133 , n52134 , n52135 , n52136 , n52137 , n52138 , n52139 , n52140 , n52141 , n52142 ,
     n52143 , n52144 , n52145 , n52146 , n52147 , n52148 , n52149 , n52150 , n52151 , n52152 ,
     n52153 , n52154 , n52155 , n52156 , n52157 , n52158 , n52159 , n52160 , n52161 , n52162 ,
     n52163 , n52164 , n52165 , n52166 , n52167 , n52168 , n52169 , n52170 , n52171 , n52172 ,
     n52173 , n52174 , n52175 , n52176 , n52177 , n52178 , n52179 , n52180 , n52181 , n52182 ,
     n52183 , n52184 , n52185 , n52186 , n52187 , n52188 , n52189 , n52190 , n52191 , n52192 ,
     n52193 , n52194 , n52195 , n52196 , n52197 , n52198 , n52199 , n52200 , n52201 , n52202 ,
     n52203 , n52204 , n52205 , n52206 , n52207 , n52208 , n52209 , n52210 , n52211 , n52212 ,
     n52213 , n52214 , n52215 , n52216 , n52217 , n52218 , n52219 , n52220 , n52221 , n52222 ,
     n52223 , n52224 , n52225 , n52226 , n52227 , n52228 , n52229 , n52230 , n52231 , n52232 ,
     n52233 , n52234 , n52235 , n52236 , n52237 , n52238 , n52239 , n52240 , n52241 , n52242 ,
     n52243 , n52244 , n52245 , n52246 , n52247 , n52248 , n52249 , n52250 , n52251 , n52252 ,
     n52253 , n52254 , n52255 , n52256 , n52257 , n52258 , n52259 , n52260 , n52261 , n52262 ,
     n52263 , n52264 , n52265 , n52266 , n52267 , n52268 , n52269 , n52270 , n52271 , n52272 ,
     n52273 , n52274 , n52275 , n52276 , n52277 , n52278 , n52279 , n52280 , n52281 , n52282 ,
     n52283 , n52284 , n52285 , n52286 , n52287 , n52288 , n52289 , n52290 , n52291 , n52292 ,
     n52293 , n52294 , n52295 , n52296 , n52297 , n52298 , n52299 , n52300 , n52301 , n52302 ,
     n52303 , n52304 , n52305 , n52306 , n52307 , n52308 , n52309 , n52310 , n52311 , n52312 ,
     n52313 , n52314 , n52315 , n52316 , n52317 , n52318 , n52319 , n52320 , n52321 , n52322 ,
     n52323 , n52324 , n52325 , n52326 , n52327 , n52328 , n52329 , n52330 , n52331 , n52332 ,
     n52333 , n52334 , n52335 , n52336 , n52337 , n52338 , n52339 , n52340 , n52341 , n52342 ,
     n52343 , n52344 , n52345 , n52346 , n52347 , n52348 , n52349 , n52350 , n52351 , n52352 ,
     n52353 , n52354 , n52355 , n52356 , n52357 , n52358 , n52359 , n52360 , n52361 , n52362 ,
     n52363 , n52364 , n52365 , n52366 , n52367 , n52368 , n52369 , n52370 , n52371 , n52372 ,
     n52373 , n52374 , n52375 , n52376 , n52377 , n52378 , n52379 , n52380 , n52381 , n52382 ,
     n52383 , n52384 , n52385 , n52386 , n52387 , n52388 , n52389 , n52390 , n52391 , n52392 ,
     n52393 , n52394 , n52395 , n52396 , n52397 , n52398 , n52399 , n52400 , n52401 , n52402 ,
     n52403 , n52404 , n52405 , n52406 , n52407 , n52408 , n52409 , n52410 , n52411 , n52412 ,
     n52413 , n52414 , n52415 , n52416 , n52417 , n52418 , n52419 , n52420 , n52421 , n52422 ,
     n52423 , n52424 , n52425 , n52426 , n52427 , n52428 , n52429 , n52430 , n52431 , n52432 ,
     n52433 , n52434 , n52435 , n52436 , n52437 , n52438 , n52439 , n52440 , n52441 , n52442 ,
     n52443 , n52444 , n52445 , n52446 , n52447 , n52448 , n52449 , n52450 , n52451 , n52452 ,
     n52453 , n52454 , n52455 , n52456 , n52457 , n52458 , n52459 , n52460 , n52461 , n52462 ,
     n52463 , n52464 , n52465 , n52466 , n52467 , n52468 , n52469 , n52470 , n52471 , n52472 ,
     n52473 , n52474 , n52475 , n52476 , n52477 , n52478 , n52479 , n52480 , n52481 , n52482 ,
     n52483 , n52484 , n52485 , n52486 , n52487 , n52488 , n52489 , n52490 , n52491 , n52492 ,
     n52493 , n52494 , n52495 , n52496 , n52497 , n52498 , n52499 , n52500 , n52501 , n52502 ,
     n52503 , n52504 , n52505 , n52506 , n52507 , n52508 , n52509 , n52510 , n52511 , n52512 ,
     n52513 , n52514 , n52515 , n52516 , n52517 , n52518 , n52519 , n52520 , n52521 , n52522 ,
     n52523 , n52524 , n52525 , n52526 , n52527 , n52528 , n52529 , n52530 , n52531 , n52532 ,
     n52533 , n52534 , n52535 , n52536 , n52537 , n52538 , n52539 , n52540 , n52541 , n52542 ,
     n52543 , n52544 , n52545 , n52546 , n52547 , n52548 , n52549 , n52550 , n52551 , n52552 ,
     n52553 , n52554 , n52555 , n52556 , n52557 , n52558 , n52559 , n52560 , n52561 , n52562 ,
     n52563 , n52564 , n52565 , n52566 , n52567 , n52568 , n52569 , n52570 , n52571 , n52572 ,
     n52573 , n52574 , n52575 , n52576 , n52577 , n52578 , n52579 , n52580 , n52581 , n52582 ,
     n52583 , n52584 , n52585 , n52586 , n52587 , n52588 , n52589 , n52590 , n52591 , n52592 ,
     n52593 , n52594 , n52595 , n52596 , n52597 , n52598 , n52599 , n52600 , n52601 , n52602 ,
     n52603 , n52604 , n52605 , n52606 , n52607 , n52608 , n52609 , n52610 , n52611 , n52612 ,
     n52613 , n52614 , n52615 , n52616 , n52617 , n52618 , n52619 , n52620 , n52621 , n52622 ,
     n52623 , n52624 , n52625 , n52626 , n52627 , n52628 , n52629 , n52630 , n52631 , n52632 ,
     n52633 , n52634 , n52635 , n52636 , n52637 , n52638 , n52639 , n52640 , n52641 , n52642 ,
     n52643 , n52644 , n52645 , n52646 , n52647 , n52648 , n52649 , n52650 , n52651 , n52652 ,
     n52653 , n52654 , n52655 , n52656 , n52657 , n52658 , n52659 , n52660 , n52661 , n52662 ,
     n52663 , n52664 , n52665 , n52666 , n52667 , n52668 , n52669 , n52670 , n52671 , n52672 ,
     n52673 , n52674 , n52675 , n52676 , n52677 , n52678 , n52679 , n52680 , n52681 , n52682 ,
     n52683 , n52684 , n52685 , n52686 , n52687 , n52688 , n52689 , n52690 , n52691 , n52692 ,
     n52693 , n52694 , n52695 , n52696 , n52697 , n52698 , n52699 , n52700 , n52701 , n52702 ,
     n52703 , n52704 , n52705 , n52706 , n52707 , n52708 , n52709 , n52710 , n52711 , n52712 ,
     n52713 , n52714 , n52715 , n52716 , n52717 , n52718 , n52719 , n52720 , n52721 , n52722 ,
     n52723 , n52724 , n52725 , n52726 , n52727 , n52728 , n52729 , n52730 , n52731 , n52732 ,
     n52733 , n52734 , n52735 , n52736 , n52737 , n52738 , n52739 , n52740 , n52741 , n52742 ,
     n52743 , n52744 , n52745 , n52746 , n52747 , n52748 , n52749 , n52750 , n52751 , n52752 ,
     n52753 , n52754 , n52755 , n52756 , n52757 , n52758 , n52759 , n52760 , n52761 , n52762 ,
     n52763 , n52764 , n52765 , n52766 , n52767 , n52768 , n52769 , n52770 , n52771 , n52772 ,
     n52773 , n52774 , n52775 , n52776 , n52777 , n52778 , n52779 , n52780 , n52781 , n52782 ,
     n52783 , n52784 , n52785 , n52786 , n52787 , n52788 , n52789 , n52790 , n52791 , n52792 ,
     n52793 , n52794 , n52795 , n52796 , n52797 , n52798 , n52799 , n52800 , n52801 , n52802 ,
     n52803 , n52804 , n52805 , n52806 , n52807 , n52808 , n52809 , n52810 , n52811 , n52812 ,
     n52813 , n52814 , n52815 , n52816 , n52817 , n52818 , n52819 , n52820 , n52821 , n52822 ,
     n52823 , n52824 , n52825 , n52826 , n52827 , n52828 , n52829 , n52830 , n52831 , n52832 ,
     n52833 , n52834 , n52835 , n52836 , n52837 , n52838 , n52839 , n52840 , n52841 , n52842 ,
     n52843 , n52844 , n52845 , n52846 , n52847 , n52848 , n52849 , n52850 , n52851 , n52852 ,
     n52853 , n52854 , n52855 , n52856 , n52857 , n52858 , n52859 , n52860 , n52861 , n52862 ,
     n52863 , n52864 , n52865 , n52866 , n52867 , n52868 , n52869 , n52870 , n52871 , n52872 ,
     n52873 , n52874 , n52875 , n52876 , n52877 , n52878 , n52879 , n52880 , n52881 , n52882 ,
     n52883 , n52884 , n52885 , n52886 , n52887 , n52888 , n52889 , n52890 , n52891 , n52892 ,
     n52893 , n52894 , n52895 , n52896 , n52897 , n52898 , n52899 , n52900 , n52901 , n52902 ,
     n52903 , n52904 , n52905 , n52906 , n52907 , n52908 , n52909 , n52910 , n52911 , n52912 ,
     n52913 , n52914 , n52915 , n52916 , n52917 , n52918 , n52919 , n52920 , n52921 , n52922 ,
     n52923 , n52924 , n52925 , n52926 , n52927 , n52928 , n52929 , n52930 , n52931 , n52932 ,
     n52933 , n52934 , n52935 , n52936 , n52937 , n52938 , n52939 , n52940 , n52941 , n52942 ,
     n52943 , n52944 , n52945 , n52946 , n52947 , n52948 , n52949 , n52950 , n52951 , n52952 ,
     n52953 , n52954 , n52955 , n52956 , n52957 , n52958 , n52959 , n52960 , n52961 , n52962 ,
     n52963 , n52964 , n52965 , n52966 , n52967 , n52968 , n52969 , n52970 , n52971 , n52972 ,
     n52973 , n52974 , n52975 , n52976 , n52977 , n52978 , n52979 , n52980 , n52981 , n52982 ,
     n52983 , n52984 , n52985 , n52986 , n52987 , n52988 , n52989 , n52990 , n52991 , n52992 ,
     n52993 , n52994 , n52995 , n52996 , n52997 , n52998 , n52999 , n53000 , n53001 , n53002 ,
     n53003 , n53004 , n53005 , n53006 , n53007 , n53008 , n53009 , n53010 , n53011 , n53012 ,
     n53013 , n53014 , n53015 , n53016 , n53017 , n53018 , n53019 , n53020 , n53021 , n53022 ,
     n53023 , n53024 , n53025 , n53026 , n53027 , n53028 , n53029 , n53030 , n53031 , n53032 ,
     n53033 , n53034 , n53035 , n53036 , n53037 , n53038 , n53039 , n53040 , n53041 , n53042 ,
     n53043 , n53044 , n53045 , n53046 , n53047 , n53048 , n53049 , n53050 , n53051 , n53052 ,
     n53053 , n53054 , n53055 , n53056 , n53057 , n53058 , n53059 , n53060 , n53061 , n53062 ,
     n53063 , n53064 , n53065 , n53066 , n53067 , n53068 , n53069 , n53070 , n53071 , n53072 ,
     n53073 , n53074 , n53075 , n53076 , n53077 , n53078 , n53079 , n53080 , n53081 , n53082 ,
     n53083 , n53084 , n53085 , n53086 , n53087 , n53088 , n53089 , n53090 , n53091 , n53092 ,
     n53093 , n53094 , n53095 , n53096 , n53097 , n53098 , n53099 , n53100 , n53101 , n53102 ,
     n53103 , n53104 , n53105 , n53106 , n53107 , n53108 , n53109 , n53110 , n53111 , n53112 ,
     n53113 , n53114 , n53115 , n53116 , n53117 , n53118 , n53119 , n53120 , n53121 , n53122 ,
     n53123 , n53124 , n53125 , n53126 , n53127 , n53128 , n53129 , n53130 , n53131 , n53132 ,
     n53133 , n53134 , n53135 , n53136 , n53137 , n53138 , n53139 , n53140 , n53141 , n53142 ,
     n53143 , n53144 , n53145 , n53146 , n53147 , n53148 , n53149 , n53150 , n53151 , n53152 ,
     n53153 , n53154 , n53155 , n53156 , n53157 , n53158 , n53159 , n53160 , n53161 , n53162 ,
     n53163 , n53164 , n53165 , n53166 , n53167 , n53168 , n53169 , n53170 , n53171 , n53172 ,
     n53173 , n53174 , n53175 , n53176 , n53177 , n53178 , n53179 , n53180 , n53181 , n53182 ,
     n53183 , n53184 , n53185 , n53186 , n53187 , n53188 , n53189 , n53190 , n53191 , n53192 ,
     n53193 , n53194 , n53195 , n53196 , n53197 , n53198 , n53199 , n53200 , n53201 , n53202 ,
     n53203 , n53204 , n53205 , n53206 , n53207 , n53208 , n53209 , n53210 , n53211 , n53212 ,
     n53213 , n53214 , n53215 , n53216 , n53217 , n53218 , n53219 , n53220 , n53221 , n53222 ,
     n53223 , n53224 , n53225 , n53226 , n53227 , n53228 , n53229 , n53230 , n53231 , n53232 ,
     n53233 , n53234 , n53235 , n53236 , n53237 , n53238 , n53239 , n53240 , n53241 , n53242 ,
     n53243 , n53244 , n53245 , n53246 , n53247 , n53248 , n53249 , n53250 , n53251 , n53252 ,
     n53253 , n53254 , n53255 , n53256 , n53257 , n53258 , n53259 , n53260 , n53261 , n53262 ,
     n53263 , n53264 , n53265 , n53266 , n53267 , n53268 , n53269 , n53270 , n53271 , n53272 ,
     n53273 , n53274 , n53275 , n53276 , n53277 , n53278 , n53279 , n53280 , n53281 , n53282 ,
     n53283 , n53284 , n53285 , n53286 , n53287 , n53288 , n53289 , n53290 , n53291 , n53292 ,
     n53293 , n53294 , n53295 , n53296 , n53297 , n53298 , n53299 , n53300 , n53301 , n53302 ,
     n53303 , n53304 , n53305 , n53306 , n53307 , n53308 , n53309 , n53310 , n53311 , n53312 ,
     n53313 , n53314 , n53315 , n53316 , n53317 , n53318 , n53319 , n53320 , n53321 , n53322 ,
     n53323 , n53324 , n53325 , n53326 , n53327 , n53328 , n53329 , n53330 , n53331 , n53332 ,
     n53333 , n53334 , n53335 , n53336 , n53337 , n53338 , n53339 , n53340 , n53341 , n53342 ,
     n53343 , n53344 , n53345 , n53346 , n53347 , n53348 , n53349 , n53350 , n53351 , n53352 ,
     n53353 , n53354 , n53355 , n53356 , n53357 , n53358 , n53359 , n53360 , n53361 , n53362 ,
     n53363 , n53364 , n53365 , n53366 , n53367 , n53368 , n53369 , n53370 , n53371 , n53372 ,
     n53373 , n53374 , n53375 , n53376 , n53377 , n53378 , n53379 , n53380 , n53381 , n53382 ,
     n53383 , n53384 , n53385 , n53386 , n53387 , n53388 , n53389 , n53390 , n53391 , n53392 ,
     n53393 , n53394 , n53395 , n53396 , n53397 , n53398 , n53399 , n53400 , n53401 , n53402 ,
     n53403 , n53404 , n53405 , n53406 , n53407 , n53408 , n53409 , n53410 , n53411 , n53412 ,
     n53413 , n53414 , n53415 , n53416 , n53417 , n53418 , n53419 , n53420 , n53421 , n53422 ,
     n53423 , n53424 , n53425 , n53426 , n53427 , n53428 , n53429 , n53430 , n53431 , n53432 ,
     n53433 , n53434 , n53435 , n53436 , n53437 , n53438 , n53439 , n53440 , n53441 , n53442 ,
     n53443 , n53444 , n53445 , n53446 , n53447 , n53448 , n53449 , n53450 , n53451 , n53452 ,
     n53453 , n53454 , n53455 , n53456 , n53457 , n53458 , n53459 , n53460 , n53461 , n53462 ,
     n53463 , n53464 , n53465 , n53466 , n53467 , n53468 , n53469 , n53470 , n53471 , n53472 ,
     n53473 , n53474 , n53475 , n53476 , n53477 , n53478 , n53479 , n53480 , n53481 , n53482 ,
     n53483 , n53484 , n53485 , n53486 , n53487 , n53488 , n53489 , n53490 , n53491 , n53492 ,
     n53493 , n53494 , n53495 , n53496 , n53497 , n53498 , n53499 , n53500 , n53501 , n53502 ,
     n53503 , n53504 , n53505 , n53506 , n53507 , n53508 , n53509 , n53510 , n53511 , n53512 ,
     n53513 , n53514 , n53515 , n53516 , n53517 , n53518 , n53519 , n53520 , n53521 , n53522 ,
     n53523 , n53524 , n53525 , n53526 , n53527 , n53528 , n53529 , n53530 , n53531 , n53532 ,
     n53533 , n53534 , n53535 , n53536 , n53537 , n53538 , n53539 , n53540 , n53541 , n53542 ,
     n53543 , n53544 , n53545 , n53546 , n53547 , n53548 , n53549 , n53550 , n53551 , n53552 ,
     n53553 , n53554 , n53555 , n53556 , n53557 , n53558 , n53559 , n53560 , n53561 , n53562 ,
     n53563 , n53564 , n53565 , n53566 , n53567 , n53568 , n53569 , n53570 , n53571 , n53572 ,
     n53573 , n53574 , n53575 , n53576 , n53577 , n53578 , n53579 , n53580 , n53581 , n53582 ,
     n53583 , n53584 , n53585 , n53586 , n53587 , n53588 , n53589 , n53590 , n53591 , n53592 ,
     n53593 , n53594 , n53595 , n53596 , n53597 , n53598 , n53599 , n53600 , n53601 , n53602 ,
     n53603 , n53604 , n53605 , n53606 , n53607 , n53608 , n53609 , n53610 , n53611 , n53612 ,
     n53613 , n53614 , n53615 , n53616 , n53617 , n53618 , n53619 , n53620 , n53621 , n53622 ,
     n53623 , n53624 , n53625 , n53626 , n53627 , n53628 , n53629 , n53630 , n53631 , n53632 ,
     n53633 , n53634 , n53635 , n53636 , n53637 , n53638 , n53639 , n53640 , n53641 , n53642 ,
     n53643 , n53644 , n53645 , n53646 , n53647 , n53648 , n53649 , n53650 , n53651 , n53652 ,
     n53653 , n53654 , n53655 , n53656 , n53657 , n53658 , n53659 , n53660 , n53661 , n53662 ,
     n53663 , n53664 , n53665 , n53666 , n53667 , n53668 , n53669 , n53670 , n53671 , n53672 ,
     n53673 , n53674 , n53675 , n53676 , n53677 , n53678 , n53679 , n53680 , n53681 , n53682 ,
     n53683 , n53684 , n53685 , n53686 , n53687 , n53688 , n53689 , n53690 , n53691 , n53692 ,
     n53693 , n53694 , n53695 , n53696 , n53697 , n53698 , n53699 , n53700 , n53701 , n53702 ,
     n53703 , n53704 , n53705 , n53706 , n53707 , n53708 , n53709 , n53710 , n53711 , n53712 ,
     n53713 , n53714 , n53715 , n53716 , n53717 , n53718 , n53719 , n53720 , n53721 , n53722 ,
     n53723 , n53724 , n53725 , n53726 , n53727 , n53728 , n53729 , n53730 , n53731 , n53732 ,
     n53733 , n53734 , n53735 , n53736 , n53737 , n53738 , n53739 , n53740 , n53741 , n53742 ,
     n53743 , n53744 , n53745 , n53746 , n53747 , n53748 , n53749 , n53750 , n53751 , n53752 ,
     n53753 , n53754 , n53755 , n53756 , n53757 , n53758 , n53759 , n53760 , n53761 , n53762 ,
     n53763 , n53764 , n53765 , n53766 , n53767 , n53768 , n53769 , n53770 , n53771 , n53772 ,
     n53773 , n53774 , n53775 , n53776 , n53777 , n53778 , n53779 , n53780 , n53781 , n53782 ,
     n53783 , n53784 , n53785 , n53786 , n53787 , n53788 , n53789 , n53790 , n53791 , n53792 ,
     n53793 , n53794 , n53795 , n53796 , n53797 , n53798 , n53799 , n53800 , n53801 , n53802 ,
     n53803 , n53804 , n53805 , n53806 , n53807 , n53808 , n53809 , n53810 , n53811 , n53812 ,
     n53813 , n53814 , n53815 , n53816 , n53817 , n53818 , n53819 , n53820 , n53821 , n53822 ,
     n53823 , n53824 , n53825 , n53826 , n53827 , n53828 , n53829 , n53830 , n53831 , n53832 ,
     n53833 , n53834 , n53835 , n53836 , n53837 , n53838 , n53839 , n53840 , n53841 , n53842 ,
     n53843 , n53844 , n53845 , n53846 , n53847 , n53848 , n53849 , n53850 , n53851 , n53852 ,
     n53853 , n53854 , n53855 , n53856 , n53857 , n53858 , n53859 , n53860 , n53861 , n53862 ,
     n53863 , n53864 , n53865 , n53866 , n53867 , n53868 , n53869 , n53870 , n53871 , n53872 ,
     n53873 , n53874 , n53875 , n53876 , n53877 , n53878 , n53879 , n53880 , n53881 , n53882 ,
     n53883 , n53884 , n53885 , n53886 , n53887 , n53888 , n53889 , n53890 , n53891 , n53892 ,
     n53893 , n53894 , n53895 , n53896 , n53897 , n53898 , n53899 , n53900 , n53901 , n53902 ,
     n53903 , n53904 , n53905 , n53906 , n53907 , n53908 , n53909 , n53910 , n53911 , n53912 ,
     n53913 , n53914 , n53915 , n53916 , n53917 , n53918 , n53919 , n53920 , n53921 , n53922 ,
     n53923 , n53924 , n53925 , n53926 , n53927 , n53928 , n53929 , n53930 , n53931 , n53932 ,
     n53933 , n53934 , n53935 , n53936 , n53937 , n53938 , n53939 , n53940 , n53941 , n53942 ,
     n53943 , n53944 , n53945 , n53946 , n53947 , n53948 , n53949 , n53950 , n53951 , n53952 ,
     n53953 , n53954 , n53955 , n53956 , n53957 , n53958 , n53959 , n53960 , n53961 , n53962 ,
     n53963 , n53964 , n53965 , n53966 , n53967 , n53968 , n53969 , n53970 , n53971 , n53972 ,
     n53973 , n53974 , n53975 , n53976 , n53977 , n53978 , n53979 , n53980 , n53981 , n53982 ,
     n53983 , n53984 , n53985 , n53986 , n53987 , n53988 , n53989 , n53990 , n53991 , n53992 ,
     n53993 , n53994 , n53995 , n53996 , n53997 , n53998 , n53999 , n54000 , n54001 , n54002 ,
     n54003 , n54004 , n54005 , n54006 , n54007 , n54008 , n54009 , n54010 , n54011 , n54012 ,
     n54013 , n54014 , n54015 , n54016 , n54017 , n54018 , n54019 , n54020 , n54021 , n54022 ,
     n54023 , n54024 , n54025 , n54026 , n54027 , n54028 , n54029 , n54030 , n54031 , n54032 ,
     n54033 , n54034 , n54035 , n54036 , n54037 , n54038 , n54039 , n54040 , n54041 , n54042 ,
     n54043 , n54044 , n54045 , n54046 , n54047 , n54048 , n54049 , n54050 , n54051 , n54052 ,
     n54053 , n54054 , n54055 , n54056 , n54057 , n54058 , n54059 , n54060 , n54061 , n54062 ,
     n54063 , n54064 , n54065 , n54066 , n54067 , n54068 , n54069 , n54070 , n54071 , n54072 ,
     n54073 , n54074 , n54075 , n54076 , n54077 , n54078 , n54079 , n54080 , n54081 , n54082 ,
     n54083 , n54084 , n54085 , n54086 , n54087 , n54088 , n54089 , n54090 , n54091 , n54092 ,
     n54093 , n54094 , n54095 , n54096 , n54097 , n54098 , n54099 , n54100 , n54101 , n54102 ,
     n54103 , n54104 , n54105 , n54106 , n54107 , n54108 , n54109 , n54110 , n54111 , n54112 ,
     n54113 , n54114 , n54115 , n54116 , n54117 , n54118 , n54119 , n54120 , n54121 , n54122 ,
     n54123 , n54124 , n54125 , n54126 , n54127 , n54128 , n54129 , n54130 , n54131 , n54132 ,
     n54133 , n54134 , n54135 , n54136 , n54137 , n54138 , n54139 , n54140 , n54141 , n54142 ,
     n54143 , n54144 , n54145 , n54146 , n54147 , n54148 , n54149 , n54150 , n54151 , n54152 ,
     n54153 , n54154 , n54155 , n54156 , n54157 , n54158 , n54159 , n54160 , n54161 , n54162 ,
     n54163 , n54164 , n54165 , n54166 , n54167 , n54168 , n54169 , n54170 , n54171 , n54172 ,
     n54173 , n54174 , n54175 , n54176 , n54177 , n54178 , n54179 , n54180 , n54181 , n54182 ,
     n54183 , n54184 , n54185 , n54186 , n54187 , n54188 , n54189 , n54190 , n54191 , n54192 ,
     n54193 , n54194 , n54195 , n54196 , n54197 , n54198 , n54199 , n54200 , n54201 , n54202 ,
     n54203 , n54204 , n54205 , n54206 , n54207 , n54208 , n54209 , n54210 , n54211 , n54212 ,
     n54213 , n54214 , n54215 , n54216 , n54217 , n54218 , n54219 , n54220 , n54221 , n54222 ,
     n54223 , n54224 , n54225 , n54226 , n54227 , n54228 , n54229 , n54230 , n54231 , n54232 ,
     n54233 , n54234 , n54235 , n54236 , n54237 , n54238 , n54239 , n54240 , n54241 , n54242 ,
     n54243 , n54244 , n54245 , n54246 , n54247 , n54248 , n54249 , n54250 , n54251 , n54252 ,
     n54253 , n54254 , n54255 , n54256 , n54257 , n54258 , n54259 , n54260 , n54261 , n54262 ,
     n54263 , n54264 , n54265 , n54266 , n54267 , n54268 , n54269 , n54270 , n54271 , n54272 ,
     n54273 , n54274 , n54275 , n54276 , n54277 , n54278 , n54279 , n54280 , n54281 , n54282 ,
     n54283 , n54284 , n54285 , n54286 , n54287 , n54288 , n54289 , n54290 , n54291 , n54292 ,
     n54293 , n54294 , n54295 , n54296 , n54297 , n54298 , n54299 , n54300 , n54301 , n54302 ,
     n54303 , n54304 , n54305 , n54306 , n54307 , n54308 , n54309 , n54310 , n54311 , n54312 ,
     n54313 , n54314 , n54315 , n54316 , n54317 , n54318 , n54319 , n54320 , n54321 , n54322 ,
     n54323 , n54324 , n54325 , n54326 , n54327 , n54328 , n54329 , n54330 , n54331 , n54332 ,
     n54333 , n54334 , n54335 , n54336 , n54337 , n54338 , n54339 , n54340 , n54341 , n54342 ,
     n54343 , n54344 , n54345 , n54346 , n54347 , n54348 , n54349 , n54350 , n54351 , n54352 ,
     n54353 , n54354 , n54355 , n54356 , n54357 , n54358 , n54359 , n54360 , n54361 , n54362 ,
     n54363 , n54364 , n54365 , n54366 , n54367 , n54368 , n54369 , n54370 , n54371 , n54372 ,
     n54373 , n54374 , n54375 , n54376 , n54377 , n54378 , n54379 , n54380 , n54381 , n54382 ,
     n54383 , n54384 , n54385 , n54386 , n54387 , n54388 , n54389 , n54390 , n54391 , n54392 ,
     n54393 , n54394 , n54395 , n54396 , n54397 , n54398 , n54399 , n54400 , n54401 , n54402 ,
     n54403 , n54404 , n54405 , n54406 , n54407 , n54408 , n54409 , n54410 , n54411 , n54412 ,
     n54413 , n54414 , n54415 , n54416 , n54417 , n54418 , n54419 , n54420 , n54421 , n54422 ,
     n54423 , n54424 , n54425 , n54426 , n54427 , n54428 , n54429 , n54430 , n54431 , n54432 ,
     n54433 , n54434 , n54435 , n54436 , n54437 , n54438 , n54439 , n54440 , n54441 , n54442 ,
     n54443 , n54444 , n54445 , n54446 , n54447 , n54448 , n54449 , n54450 , n54451 , n54452 ,
     n54453 , n54454 , n54455 , n54456 , n54457 , n54458 , n54459 , n54460 , n54461 , n54462 ,
     n54463 , n54464 , n54465 , n54466 , n54467 , n54468 , n54469 , n54470 , n54471 , n54472 ,
     n54473 , n54474 , n54475 , n54476 , n54477 , n54478 , n54479 , n54480 , n54481 , n54482 ,
     n54483 , n54484 , n54485 , n54486 , n54487 , n54488 , n54489 , n54490 , n54491 , n54492 ,
     n54493 , n54494 , n54495 , n54496 , n54497 , n54498 , n54499 , n54500 , n54501 , n54502 ,
     n54503 , n54504 , n54505 , n54506 , n54507 , n54508 , n54509 , n54510 , n54511 , n54512 ,
     n54513 , n54514 , n54515 , n54516 , n54517 , n54518 , n54519 , n54520 , n54521 , n54522 ,
     n54523 , n54524 , n54525 , n54526 , n54527 , n54528 , n54529 , n54530 , n54531 , n54532 ,
     n54533 , n54534 , n54535 , n54536 , n54537 , n54538 , n54539 , n54540 , n54541 , n54542 ,
     n54543 , n54544 , n54545 , n54546 , n54547 , n54548 , n54549 , n54550 , n54551 , n54552 ,
     n54553 , n54554 , n54555 , n54556 , n54557 , n54558 , n54559 , n54560 , n54561 , n54562 ,
     n54563 , n54564 , n54565 , n54566 , n54567 , n54568 , n54569 , n54570 , n54571 , n54572 ,
     n54573 , n54574 , n54575 , n54576 , n54577 , n54578 , n54579 , n54580 , n54581 , n54582 ,
     n54583 , n54584 , n54585 , n54586 , n54587 , n54588 , n54589 , n54590 , n54591 , n54592 ,
     n54593 , n54594 , n54595 , n54596 , n54597 , n54598 , n54599 , n54600 , n54601 , n54602 ,
     n54603 , n54604 , n54605 , n54606 , n54607 , n54608 , n54609 , n54610 , n54611 , n54612 ,
     n54613 , n54614 , n54615 , n54616 , n54617 , n54618 , n54619 , n54620 , n54621 , n54622 ,
     n54623 , n54624 , n54625 , n54626 , n54627 , n54628 , n54629 , n54630 , n54631 , n54632 ,
     n54633 , n54634 , n54635 , n54636 , n54637 , n54638 , n54639 , n54640 , n54641 , n54642 ,
     n54643 , n54644 , n54645 , n54646 , n54647 , n54648 , n54649 , n54650 , n54651 , n54652 ,
     n54653 , n54654 , n54655 , n54656 , n54657 , n54658 , n54659 , n54660 , n54661 , n54662 ,
     n54663 , n54664 , n54665 , n54666 , n54667 , n54668 , n54669 , n54670 , n54671 , n54672 ,
     n54673 , n54674 , n54675 , n54676 , n54677 , n54678 , n54679 , n54680 , n54681 , n54682 ,
     n54683 , n54684 , n54685 , n54686 , n54687 , n54688 , n54689 , n54690 , n54691 , n54692 ,
     n54693 , n54694 , n54695 , n54696 , n54697 , n54698 , n54699 , n54700 , n54701 , n54702 ,
     n54703 , n54704 , n54705 , n54706 , n54707 , n54708 , n54709 , n54710 , n54711 , n54712 ,
     n54713 , n54714 , n54715 , n54716 , n54717 , n54718 , n54719 , n54720 , n54721 , n54722 ,
     n54723 , n54724 , n54725 , n54726 , n54727 , n54728 , n54729 , n54730 , n54731 , n54732 ,
     n54733 , n54734 , n54735 , n54736 , n54737 , n54738 , n54739 , n54740 , n54741 , n54742 ,
     n54743 , n54744 , n54745 , n54746 , n54747 , n54748 , n54749 , n54750 , n54751 , n54752 ,
     n54753 , n54754 , n54755 , n54756 , n54757 , n54758 , n54759 , n54760 , n54761 , n54762 ,
     n54763 , n54764 , n54765 , n54766 , n54767 , n54768 , n54769 , n54770 , n54771 , n54772 ,
     n54773 , n54774 , n54775 , n54776 , n54777 , n54778 , n54779 , n54780 , n54781 , n54782 ,
     n54783 , n54784 , n54785 , n54786 , n54787 , n54788 , n54789 , n54790 , n54791 , n54792 ,
     n54793 , n54794 , n54795 , n54796 , n54797 , n54798 , n54799 , n54800 , n54801 , n54802 ,
     n54803 , n54804 , n54805 , n54806 , n54807 , n54808 , n54809 , n54810 , n54811 , n54812 ,
     n54813 , n54814 , n54815 , n54816 , n54817 , n54818 , n54819 , n54820 , n54821 , n54822 ,
     n54823 , n54824 , n54825 , n54826 , n54827 , n54828 , n54829 , n54830 , n54831 , n54832 ,
     n54833 , n54834 , n54835 , n54836 , n54837 , n54838 , n54839 , n54840 , n54841 , n54842 ,
     n54843 , n54844 , n54845 , n54846 , n54847 , n54848 , n54849 , n54850 , n54851 , n54852 ,
     n54853 , n54854 , n54855 , n54856 , n54857 , n54858 , n54859 , n54860 , n54861 , n54862 ,
     n54863 , n54864 , n54865 , n54866 , n54867 , n54868 , n54869 , n54870 , n54871 , n54872 ,
     n54873 , n54874 , n54875 , n54876 , n54877 , n54878 , n54879 , n54880 , n54881 , n54882 ,
     n54883 , n54884 , n54885 , n54886 , n54887 , n54888 , n54889 , n54890 , n54891 , n54892 ,
     n54893 , n54894 , n54895 , n54896 , n54897 , n54898 , n54899 , n54900 , n54901 , n54902 ,
     n54903 , n54904 , n54905 , n54906 , n54907 , n54908 , n54909 , n54910 , n54911 , n54912 ,
     n54913 , n54914 , n54915 , n54916 , n54917 , n54918 , n54919 , n54920 , n54921 , n54922 ,
     n54923 , n54924 , n54925 , n54926 , n54927 , n54928 , n54929 , n54930 , n54931 , n54932 ,
     n54933 , n54934 , n54935 , n54936 , n54937 , n54938 , n54939 , n54940 , n54941 , n54942 ,
     n54943 , n54944 , n54945 , n54946 , n54947 , n54948 , n54949 , n54950 , n54951 , n54952 ,
     n54953 , n54954 , n54955 , n54956 , n54957 , n54958 , n54959 , n54960 , n54961 , n54962 ,
     n54963 , n54964 , n54965 , n54966 , n54967 , n54968 , n54969 , n54970 , n54971 , n54972 ,
     n54973 , n54974 , n54975 , n54976 , n54977 , n54978 , n54979 , n54980 , n54981 , n54982 ,
     n54983 , n54984 , n54985 , n54986 , n54987 , n54988 , n54989 , n54990 , n54991 , n54992 ,
     n54993 , n54994 , n54995 , n54996 , n54997 , n54998 , n54999 , n55000 , n55001 , n55002 ,
     n55003 , n55004 , n55005 , n55006 , n55007 , n55008 , n55009 , n55010 , n55011 , n55012 ,
     n55013 , n55014 , n55015 , n55016 , n55017 , n55018 , n55019 , n55020 , n55021 , n55022 ,
     n55023 , n55024 , n55025 , n55026 , n55027 , n55028 , n55029 , n55030 , n55031 , n55032 ,
     n55033 , n55034 , n55035 , n55036 , n55037 , n55038 , n55039 , n55040 , n55041 , n55042 ,
     n55043 , n55044 , n55045 , n55046 , n55047 , n55048 , n55049 , n55050 , n55051 , n55052 ,
     n55053 , n55054 , n55055 , n55056 , n55057 , n55058 , n55059 , n55060 , n55061 , n55062 ,
     n55063 , n55064 , n55065 , n55066 , n55067 , n55068 , n55069 , n55070 , n55071 , n55072 ,
     n55073 , n55074 , n55075 , n55076 , n55077 , n55078 , n55079 , n55080 , n55081 , n55082 ,
     n55083 , n55084 , n55085 , n55086 , n55087 , n55088 , n55089 , n55090 , n55091 , n55092 ,
     n55093 , n55094 , n55095 , n55096 , n55097 , n55098 , n55099 , n55100 , n55101 , n55102 ,
     n55103 , n55104 , n55105 , n55106 , n55107 , n55108 , n55109 , n55110 , n55111 , n55112 ,
     n55113 , n55114 , n55115 , n55116 , n55117 , n55118 , n55119 , n55120 , n55121 , n55122 ,
     n55123 , n55124 , n55125 , n55126 , n55127 , n55128 , n55129 , n55130 , n55131 , n55132 ,
     n55133 , n55134 , n55135 , n55136 , n55137 , n55138 , n55139 , n55140 , n55141 , n55142 ,
     n55143 , n55144 , n55145 , n55146 , n55147 , n55148 , n55149 , n55150 , n55151 , n55152 ,
     n55153 , n55154 , n55155 , n55156 , n55157 , n55158 , n55159 , n55160 , n55161 , n55162 ,
     n55163 , n55164 , n55165 , n55166 , n55167 , n55168 , n55169 , n55170 , n55171 , n55172 ,
     n55173 , n55174 , n55175 , n55176 , n55177 , n55178 , n55179 , n55180 , n55181 , n55182 ,
     n55183 , n55184 , n55185 , n55186 , n55187 , n55188 , n55189 , n55190 , n55191 , n55192 ,
     n55193 , n55194 , n55195 , n55196 , n55197 , n55198 , n55199 , n55200 , n55201 , n55202 ,
     n55203 , n55204 , n55205 , n55206 , n55207 , n55208 , n55209 , n55210 , n55211 , n55212 ,
     n55213 , n55214 , n55215 , n55216 , n55217 , n55218 , n55219 , n55220 , n55221 , n55222 ,
     n55223 , n55224 , n55225 , n55226 , n55227 , n55228 , n55229 , n55230 , n55231 , n55232 ,
     n55233 , n55234 , n55235 , n55236 , n55237 , n55238 , n55239 , n55240 , n55241 , n55242 ,
     n55243 , n55244 , n55245 , n55246 , n55247 , n55248 , n55249 , n55250 , n55251 , n55252 ,
     n55253 , n55254 , n55255 , n55256 , n55257 , n55258 , n55259 , n55260 , n55261 , n55262 ,
     n55263 , n55264 , n55265 , n55266 , n55267 , n55268 , n55269 , n55270 , n55271 , n55272 ,
     n55273 , n55274 , n55275 , n55276 , n55277 , n55278 , n55279 , n55280 , n55281 , n55282 ,
     n55283 , n55284 , n55285 , n55286 , n55287 , n55288 , n55289 , n55290 , n55291 , n55292 ,
     n55293 , n55294 , n55295 , n55296 , n55297 , n55298 , n55299 , n55300 , n55301 , n55302 ,
     n55303 , n55304 , n55305 , n55306 , n55307 , n55308 , n55309 , n55310 , n55311 , n55312 ,
     n55313 , n55314 , n55315 , n55316 , n55317 , n55318 , n55319 , n55320 , n55321 , n55322 ,
     n55323 , n55324 , n55325 , n55326 , n55327 , n55328 , n55329 , n55330 , n55331 , n55332 ,
     n55333 , n55334 , n55335 , n55336 , n55337 , n55338 , n55339 , n55340 , n55341 , n55342 ,
     n55343 , n55344 , n55345 , n55346 , n55347 , n55348 , n55349 , n55350 , n55351 , n55352 ,
     n55353 , n55354 , n55355 , n55356 , n55357 , n55358 , n55359 , n55360 , n55361 , n55362 ,
     n55363 , n55364 , n55365 , n55366 , n55367 , n55368 , n55369 , n55370 , n55371 , n55372 ,
     n55373 , n55374 , n55375 , n55376 , n55377 , n55378 , n55379 , n55380 , n55381 , n55382 ,
     n55383 , n55384 , n55385 , n55386 , n55387 , n55388 , n55389 , n55390 , n55391 , n55392 ,
     n55393 , n55394 , n55395 , n55396 , n55397 , n55398 , n55399 , n55400 , n55401 , n55402 ,
     n55403 , n55404 , n55405 , n55406 , n55407 , n55408 , n55409 , n55410 , n55411 , n55412 ,
     n55413 , n55414 , n55415 , n55416 , n55417 , n55418 , n55419 , n55420 , n55421 , n55422 ,
     n55423 , n55424 , n55425 , n55426 , n55427 , n55428 , n55429 , n55430 , n55431 , n55432 ,
     n55433 , n55434 , n55435 , n55436 , n55437 , n55438 , n55439 , n55440 , n55441 , n55442 ,
     n55443 , n55444 , n55445 , n55446 , n55447 , n55448 , n55449 , n55450 , n55451 , n55452 ,
     n55453 , n55454 , n55455 , n55456 , n55457 , n55458 , n55459 , n55460 , n55461 , n55462 ,
     n55463 , n55464 , n55465 , n55466 , n55467 , n55468 , n55469 , n55470 , n55471 , n55472 ,
     n55473 , n55474 , n55475 , n55476 , n55477 , n55478 , n55479 , n55480 , n55481 , n55482 ,
     n55483 , n55484 , n55485 , n55486 , n55487 , n55488 , n55489 , n55490 , n55491 , n55492 ,
     n55493 , n55494 , n55495 , n55496 , n55497 , n55498 , n55499 , n55500 , n55501 , n55502 ,
     n55503 , n55504 , n55505 , n55506 , n55507 , n55508 , n55509 , n55510 , n55511 , n55512 ,
     n55513 , n55514 , n55515 , n55516 , n55517 , n55518 , n55519 , n55520 , n55521 , n55522 ,
     n55523 , n55524 , n55525 , n55526 , n55527 , n55528 , n55529 , n55530 , n55531 , n55532 ,
     n55533 , n55534 , n55535 , n55536 , n55537 , n55538 , n55539 , n55540 , n55541 , n55542 ,
     n55543 , n55544 , n55545 , n55546 , n55547 , n55548 , n55549 , n55550 , n55551 , n55552 ,
     n55553 , n55554 , n55555 , n55556 , n55557 , n55558 , n55559 , n55560 , n55561 , n55562 ,
     n55563 , n55564 , n55565 , n55566 , n55567 , n55568 , n55569 , n55570 , n55571 , n55572 ,
     n55573 , n55574 , n55575 , n55576 , n55577 , n55578 , n55579 , n55580 , n55581 , n55582 ,
     n55583 , n55584 , n55585 , n55586 , n55587 , n55588 , n55589 , n55590 , n55591 , n55592 ,
     n55593 , n55594 , n55595 , n55596 , n55597 , n55598 , n55599 , n55600 , n55601 , n55602 ,
     n55603 , n55604 , n55605 , n55606 , n55607 , n55608 , n55609 , n55610 , n55611 , n55612 ,
     n55613 , n55614 , n55615 , n55616 , n55617 , n55618 , n55619 , n55620 , n55621 , n55622 ,
     n55623 , n55624 , n55625 , n55626 , n55627 , n55628 , n55629 , n55630 , n55631 , n55632 ,
     n55633 , n55634 , n55635 , n55636 , n55637 , n55638 , n55639 , n55640 , n55641 , n55642 ,
     n55643 , n55644 , n55645 , n55646 , n55647 , n55648 , n55649 , n55650 , n55651 , n55652 ,
     n55653 , n55654 , n55655 , n55656 , n55657 , n55658 , n55659 , n55660 , n55661 , n55662 ,
     n55663 , n55664 , n55665 , n55666 , n55667 , n55668 , n55669 , n55670 , n55671 , n55672 ,
     n55673 , n55674 , n55675 , n55676 , n55677 , n55678 , n55679 , n55680 , n55681 , n55682 ,
     n55683 , n55684 , n55685 , n55686 , n55687 , n55688 , n55689 , n55690 , n55691 , n55692 ,
     n55693 , n55694 , n55695 , n55696 , n55697 , n55698 , n55699 , n55700 , n55701 , n55702 ,
     n55703 , n55704 , n55705 , n55706 , n55707 , n55708 , n55709 , n55710 , n55711 , n55712 ,
     n55713 , n55714 , n55715 , n55716 , n55717 , n55718 , n55719 , n55720 , n55721 , n55722 ,
     n55723 , n55724 , n55725 , n55726 , n55727 , n55728 , n55729 , n55730 , n55731 , n55732 ,
     n55733 , n55734 , n55735 , n55736 , n55737 , n55738 , n55739 , n55740 , n55741 , n55742 ,
     n55743 , n55744 , n55745 , n55746 , n55747 , n55748 , n55749 , n55750 , n55751 , n55752 ,
     n55753 , n55754 , n55755 , n55756 , n55757 , n55758 , n55759 , n55760 , n55761 , n55762 ,
     n55763 , n55764 , n55765 , n55766 , n55767 , n55768 , n55769 , n55770 , n55771 , n55772 ,
     n55773 , n55774 , n55775 , n55776 , n55777 , n55778 , n55779 , n55780 , n55781 , n55782 ,
     n55783 , n55784 , n55785 , n55786 , n55787 , n55788 , n55789 , n55790 , n55791 , n55792 ,
     n55793 , n55794 , n55795 , n55796 , n55797 , n55798 , n55799 , n55800 , n55801 , n55802 ,
     n55803 , n55804 , n55805 , n55806 , n55807 , n55808 , n55809 , n55810 , n55811 , n55812 ,
     n55813 , n55814 , n55815 , n55816 , n55817 , n55818 , n55819 , n55820 , n55821 , n55822 ,
     n55823 , n55824 , n55825 , n55826 , n55827 , n55828 , n55829 , n55830 , n55831 , n55832 ,
     n55833 , n55834 , n55835 , n55836 , n55837 , n55838 , n55839 , n55840 , n55841 , n55842 ,
     n55843 , n55844 , n55845 , n55846 , n55847 , n55848 , n55849 , n55850 , n55851 , n55852 ,
     n55853 , n55854 , n55855 , n55856 , n55857 , n55858 , n55859 , n55860 , n55861 , n55862 ,
     n55863 , n55864 , n55865 , n55866 , n55867 , n55868 , n55869 , n55870 , n55871 , n55872 ,
     n55873 , n55874 , n55875 , n55876 , n55877 , n55878 , n55879 , n55880 , n55881 , n55882 ,
     n55883 , n55884 , n55885 , n55886 , n55887 , n55888 , n55889 , n55890 , n55891 , n55892 ,
     n55893 , n55894 , n55895 , n55896 , n55897 , n55898 , n55899 , n55900 , n55901 , n55902 ,
     n55903 , n55904 , n55905 , n55906 , n55907 , n55908 , n55909 , n55910 , n55911 , n55912 ,
     n55913 , n55914 , n55915 , n55916 , n55917 , n55918 , n55919 , n55920 , n55921 , n55922 ,
     n55923 , n55924 , n55925 , n55926 , n55927 , n55928 , n55929 , n55930 , n55931 , n55932 ,
     n55933 , n55934 , n55935 , n55936 , n55937 , n55938 , n55939 , n55940 , n55941 , n55942 ,
     n55943 , n55944 , n55945 , n55946 , n55947 , n55948 , n55949 , n55950 , n55951 , n55952 ,
     n55953 , n55954 , n55955 , n55956 , n55957 , n55958 , n55959 , n55960 , n55961 , n55962 ,
     n55963 , n55964 , n55965 , n55966 , n55967 , n55968 , n55969 , n55970 , n55971 , n55972 ,
     n55973 , n55974 , n55975 , n55976 , n55977 , n55978 , n55979 , n55980 , n55981 , n55982 ,
     n55983 , n55984 , n55985 , n55986 , n55987 , n55988 , n55989 , n55990 , n55991 , n55992 ,
     n55993 , n55994 , n55995 , n55996 , n55997 , n55998 , n55999 , n56000 , n56001 , n56002 ,
     n56003 , n56004 , n56005 , n56006 , n56007 , n56008 , n56009 , n56010 , n56011 , n56012 ,
     n56013 , n56014 , n56015 , n56016 , n56017 , n56018 , n56019 , n56020 , n56021 , n56022 ,
     n56023 , n56024 , n56025 , n56026 , n56027 , n56028 , n56029 , n56030 , n56031 , n56032 ,
     n56033 , n56034 , n56035 , n56036 , n56037 , n56038 , n56039 , n56040 , n56041 , n56042 ,
     n56043 , n56044 , n56045 , n56046 , n56047 , n56048 , n56049 , n56050 , n56051 , n56052 ,
     n56053 , n56054 , n56055 , n56056 , n56057 , n56058 , n56059 , n56060 , n56061 , n56062 ,
     n56063 , n56064 , n56065 , n56066 , n56067 , n56068 , n56069 , n56070 , n56071 , n56072 ,
     n56073 , n56074 , n56075 , n56076 , n56077 , n56078 , n56079 , n56080 , n56081 , n56082 ,
     n56083 , n56084 , n56085 , n56086 , n56087 , n56088 , n56089 , n56090 , n56091 , n56092 ,
     n56093 , n56094 , n56095 , n56096 , n56097 , n56098 , n56099 , n56100 , n56101 , n56102 ,
     n56103 , n56104 , n56105 , n56106 , n56107 , n56108 , n56109 , n56110 , n56111 , n56112 ,
     n56113 , n56114 , n56115 , n56116 , n56117 , n56118 , n56119 , n56120 , n56121 , n56122 ,
     n56123 , n56124 , n56125 , n56126 , n56127 , n56128 , n56129 , n56130 , n56131 , n56132 ,
     n56133 , n56134 , n56135 , n56136 , n56137 , n56138 , n56139 , n56140 , n56141 , n56142 ,
     n56143 , n56144 , n56145 , n56146 , n56147 , n56148 , n56149 , n56150 , n56151 , n56152 ,
     n56153 , n56154 , n56155 , n56156 , n56157 , n56158 , n56159 , n56160 , n56161 , n56162 ,
     n56163 , n56164 , n56165 , n56166 , n56167 , n56168 , n56169 , n56170 , n56171 , n56172 ,
     n56173 , n56174 , n56175 , n56176 , n56177 , n56178 , n56179 , n56180 , n56181 , n56182 ,
     n56183 , n56184 , n56185 , n56186 , n56187 , n56188 , n56189 , n56190 , n56191 , n56192 ,
     n56193 , n56194 , n56195 , n56196 , n56197 , n56198 , n56199 , n56200 , n56201 , n56202 ,
     n56203 , n56204 , n56205 , n56206 , n56207 , n56208 , n56209 , n56210 , n56211 , n56212 ,
     n56213 , n56214 , n56215 , n56216 , n56217 , n56218 , n56219 , n56220 , n56221 , n56222 ,
     n56223 , n56224 , n56225 , n56226 , n56227 , n56228 , n56229 , n56230 , n56231 , n56232 ,
     n56233 , n56234 , n56235 , n56236 , n56237 , n56238 , n56239 , n56240 , n56241 , n56242 ,
     n56243 , n56244 , n56245 , n56246 , n56247 , n56248 , n56249 , n56250 , n56251 , n56252 ,
     n56253 , n56254 , n56255 , n56256 , n56257 , n56258 , n56259 , n56260 , n56261 , n56262 ,
     n56263 , n56264 , n56265 , n56266 , n56267 , n56268 , n56269 , n56270 , n56271 , n56272 ,
     n56273 , n56274 , n56275 , n56276 , n56277 , n56278 , n56279 , n56280 , n56281 , n56282 ,
     n56283 , n56284 , n56285 , n56286 , n56287 , n56288 , n56289 , n56290 , n56291 , n56292 ,
     n56293 , n56294 , n56295 , n56296 , n56297 , n56298 , n56299 , n56300 , n56301 , n56302 ,
     n56303 , n56304 , n56305 , n56306 , n56307 , n56308 , n56309 , n56310 , n56311 , n56312 ,
     n56313 , n56314 , n56315 , n56316 , n56317 , n56318 , n56319 , n56320 , n56321 , n56322 ,
     n56323 , n56324 , n56325 , n56326 , n56327 , n56328 , n56329 , n56330 , n56331 , n56332 ,
     n56333 , n56334 , n56335 , n56336 , n56337 , n56338 , n56339 , n56340 , n56341 , n56342 ,
     n56343 , n56344 , n56345 , n56346 , n56347 , n56348 , n56349 , n56350 , n56351 , n56352 ,
     n56353 , n56354 , n56355 , n56356 , n56357 , n56358 , n56359 , n56360 , n56361 , n56362 ,
     n56363 , n56364 , n56365 , n56366 , n56367 , n56368 , n56369 , n56370 , n56371 , n56372 ,
     n56373 , n56374 , n56375 , n56376 , n56377 , n56378 , n56379 , n56380 , n56381 , n56382 ,
     n56383 , n56384 , n56385 , n56386 , n56387 , n56388 , n56389 , n56390 , n56391 , n56392 ,
     n56393 , n56394 , n56395 , n56396 , n56397 , n56398 , n56399 , n56400 , n56401 , n56402 ,
     n56403 , n56404 , n56405 , n56406 , n56407 , n56408 , n56409 , n56410 , n56411 , n56412 ,
     n56413 , n56414 , n56415 , n56416 , n56417 , n56418 , n56419 , n56420 , n56421 , n56422 ,
     n56423 , n56424 , n56425 , n56426 , n56427 , n56428 , n56429 , n56430 , n56431 , n56432 ,
     n56433 , n56434 , n56435 , n56436 , n56437 , n56438 , n56439 , n56440 , n56441 , n56442 ,
     n56443 , n56444 , n56445 , n56446 , n56447 , n56448 , n56449 , n56450 , n56451 , n56452 ,
     n56453 , n56454 , n56455 , n56456 , n56457 , n56458 , n56459 , n56460 , n56461 , n56462 ,
     n56463 , n56464 , n56465 , n56466 , n56467 , n56468 , n56469 , n56470 , n56471 , n56472 ,
     n56473 , n56474 , n56475 , n56476 , n56477 , n56478 , n56479 , n56480 , n56481 , n56482 ,
     n56483 , n56484 , n56485 , n56486 , n56487 , n56488 , n56489 , n56490 , n56491 , n56492 ,
     n56493 , n56494 , n56495 , n56496 , n56497 , n56498 , n56499 , n56500 , n56501 , n56502 ,
     n56503 , n56504 , n56505 , n56506 , n56507 , n56508 , n56509 , n56510 , n56511 , n56512 ,
     n56513 , n56514 , n56515 , n56516 , n56517 , n56518 , n56519 , n56520 , n56521 , n56522 ,
     n56523 , n56524 , n56525 , n56526 , n56527 , n56528 , n56529 , n56530 , n56531 , n56532 ,
     n56533 , n56534 , n56535 , n56536 , n56537 , n56538 , n56539 , n56540 , n56541 , n56542 ,
     n56543 , n56544 , n56545 , n56546 , n56547 , n56548 , n56549 , n56550 , n56551 , n56552 ,
     n56553 , n56554 , n56555 , n56556 , n56557 , n56558 , n56559 , n56560 , n56561 , n56562 ,
     n56563 , n56564 , n56565 , n56566 , n56567 , n56568 , n56569 , n56570 , n56571 , n56572 ,
     n56573 , n56574 , n56575 , n56576 , n56577 , n56578 , n56579 , n56580 , n56581 , n56582 ,
     n56583 , n56584 , n56585 , n56586 , n56587 , n56588 , n56589 , n56590 , n56591 , n56592 ,
     n56593 , n56594 , n56595 , n56596 , n56597 , n56598 , n56599 , n56600 , n56601 , n56602 ,
     n56603 , n56604 , n56605 , n56606 , n56607 , n56608 , n56609 , n56610 , n56611 , n56612 ,
     n56613 , n56614 , n56615 , n56616 , n56617 , n56618 , n56619 , n56620 , n56621 , n56622 ,
     n56623 , n56624 , n56625 , n56626 , n56627 , n56628 , n56629 , n56630 , n56631 , n56632 ,
     n56633 , n56634 , n56635 , n56636 , n56637 , n56638 , n56639 , n56640 , n56641 , n56642 ,
     n56643 , n56644 , n56645 , n56646 , n56647 , n56648 , n56649 , n56650 , n56651 , n56652 ,
     n56653 , n56654 , n56655 , n56656 , n56657 , n56658 , n56659 , n56660 , n56661 , n56662 ,
     n56663 , n56664 , n56665 , n56666 , n56667 , n56668 , n56669 , n56670 , n56671 , n56672 ,
     n56673 , n56674 , n56675 , n56676 , n56677 , n56678 , n56679 , n56680 , n56681 , n56682 ,
     n56683 , n56684 , n56685 , n56686 , n56687 , n56688 , n56689 , n56690 , n56691 , n56692 ,
     n56693 , n56694 , n56695 , n56696 , n56697 , n56698 , n56699 , n56700 , n56701 , n56702 ,
     n56703 , n56704 , n56705 , n56706 , n56707 , n56708 , n56709 , n56710 , n56711 , n56712 ,
     n56713 , n56714 , n56715 , n56716 , n56717 , n56718 , n56719 , n56720 , n56721 , n56722 ,
     n56723 , n56724 , n56725 , n56726 , n56727 , n56728 , n56729 , n56730 , n56731 , n56732 ,
     n56733 , n56734 , n56735 , n56736 , n56737 , n56738 , n56739 , n56740 , n56741 , n56742 ,
     n56743 , n56744 , n56745 , n56746 , n56747 , n56748 , n56749 , n56750 , n56751 , n56752 ,
     n56753 , n56754 , n56755 , n56756 , n56757 , n56758 , n56759 , n56760 , n56761 , n56762 ,
     n56763 , n56764 , n56765 , n56766 , n56767 , n56768 , n56769 , n56770 , n56771 , n56772 ,
     n56773 , n56774 , n56775 , n56776 , n56777 , n56778 , n56779 , n56780 , n56781 , n56782 ,
     n56783 , n56784 , n56785 , n56786 , n56787 , n56788 , n56789 , n56790 , n56791 , n56792 ,
     n56793 , n56794 , n56795 , n56796 , n56797 , n56798 , n56799 , n56800 , n56801 , n56802 ,
     n56803 , n56804 , n56805 , n56806 , n56807 , n56808 , n56809 , n56810 , n56811 , n56812 ,
     n56813 , n56814 , n56815 , n56816 , n56817 , n56818 , n56819 , n56820 , n56821 , n56822 ,
     n56823 , n56824 , n56825 , n56826 , n56827 , n56828 , n56829 , n56830 , n56831 , n56832 ,
     n56833 , n56834 , n56835 , n56836 , n56837 , n56838 , n56839 , n56840 , n56841 , n56842 ,
     n56843 , n56844 , n56845 , n56846 , n56847 , n56848 , n56849 , n56850 , n56851 , n56852 ,
     n56853 , n56854 , n56855 , n56856 , n56857 , n56858 , n56859 , n56860 , n56861 , n56862 ,
     n56863 , n56864 , n56865 , n56866 , n56867 , n56868 , n56869 , n56870 , n56871 , n56872 ,
     n56873 , n56874 , n56875 , n56876 , n56877 , n56878 , n56879 , n56880 , n56881 , n56882 ,
     n56883 , n56884 , n56885 , n56886 , n56887 , n56888 , n56889 , n56890 , n56891 , n56892 ,
     n56893 , n56894 , n56895 , n56896 , n56897 , n56898 , n56899 , n56900 , n56901 , n56902 ,
     n56903 , n56904 , n56905 , n56906 , n56907 , n56908 , n56909 , n56910 , n56911 , n56912 ,
     n56913 , n56914 , n56915 , n56916 , n56917 , n56918 , n56919 , n56920 , n56921 , n56922 ,
     n56923 , n56924 , n56925 , n56926 , n56927 , n56928 , n56929 , n56930 , n56931 , n56932 ,
     n56933 , n56934 , n56935 , n56936 , n56937 , n56938 , n56939 , n56940 , n56941 , n56942 ,
     n56943 , n56944 , n56945 , n56946 , n56947 , n56948 , n56949 , n56950 , n56951 , n56952 ,
     n56953 , n56954 , n56955 , n56956 , n56957 , n56958 , n56959 , n56960 , n56961 , n56962 ,
     n56963 , n56964 , n56965 , n56966 , n56967 , n56968 , n56969 , n56970 , n56971 , n56972 ,
     n56973 , n56974 , n56975 , n56976 , n56977 , n56978 , n56979 , n56980 , n56981 , n56982 ,
     n56983 , n56984 , n56985 , n56986 , n56987 , n56988 , n56989 , n56990 , n56991 , n56992 ,
     n56993 , n56994 , n56995 , n56996 , n56997 , n56998 , n56999 , n57000 , n57001 , n57002 ,
     n57003 , n57004 , n57005 , n57006 , n57007 , n57008 , n57009 , n57010 , n57011 , n57012 ,
     n57013 , n57014 , n57015 , n57016 , n57017 , n57018 , n57019 , n57020 , n57021 , n57022 ,
     n57023 , n57024 , n57025 , n57026 , n57027 , n57028 , n57029 , n57030 , n57031 , n57032 ,
     n57033 , n57034 , n57035 , n57036 , n57037 , n57038 , n57039 , n57040 , n57041 , n57042 ,
     n57043 , n57044 , n57045 , n57046 , n57047 , n57048 , n57049 , n57050 , n57051 , n57052 ,
     n57053 , n57054 , n57055 , n57056 , n57057 , n57058 , n57059 , n57060 , n57061 , n57062 ,
     n57063 , n57064 , n57065 , n57066 , n57067 , n57068 , n57069 , n57070 , n57071 , n57072 ,
     n57073 , n57074 , n57075 , n57076 , n57077 , n57078 , n57079 , n57080 , n57081 , n57082 ,
     n57083 , n57084 , n57085 , n57086 , n57087 , n57088 , n57089 , n57090 , n57091 , n57092 ,
     n57093 , n57094 , n57095 , n57096 , n57097 , n57098 , n57099 , n57100 , n57101 , n57102 ,
     n57103 , n57104 , n57105 , n57106 , n57107 , n57108 , n57109 , n57110 , n57111 , n57112 ,
     n57113 , n57114 , n57115 , n57116 , n57117 , n57118 , n57119 , n57120 , n57121 , n57122 ,
     n57123 , n57124 , n57125 , n57126 , n57127 , n57128 , n57129 , n57130 , n57131 , n57132 ,
     n57133 , n57134 , n57135 , n57136 , n57137 , n57138 , n57139 , n57140 , n57141 , n57142 ,
     n57143 , n57144 , n57145 , n57146 , n57147 , n57148 , n57149 , n57150 , n57151 , n57152 ,
     n57153 , n57154 , n57155 , n57156 , n57157 , n57158 , n57159 , n57160 , n57161 , n57162 ,
     n57163 , n57164 , n57165 , n57166 , n57167 , n57168 , n57169 , n57170 , n57171 , n57172 ,
     n57173 , n57174 , n57175 , n57176 , n57177 , n57178 , n57179 , n57180 , n57181 , n57182 ,
     n57183 , n57184 , n57185 , n57186 , n57187 , n57188 , n57189 , n57190 , n57191 , n57192 ,
     n57193 , n57194 , n57195 , n57196 , n57197 , n57198 , n57199 , n57200 , n57201 , n57202 ,
     n57203 , n57204 , n57205 , n57206 , n57207 , n57208 , n57209 , n57210 , n57211 , n57212 ,
     n57213 , n57214 , n57215 , n57216 , n57217 , n57218 , n57219 , n57220 , n57221 , n57222 ,
     n57223 , n57224 , n57225 , n57226 , n57227 , n57228 , n57229 , n57230 , n57231 , n57232 ,
     n57233 , n57234 , n57235 , n57236 , n57237 , n57238 , n57239 , n57240 , n57241 , n57242 ,
     n57243 , n57244 , n57245 , n57246 , n57247 , n57248 , n57249 , n57250 , n57251 , n57252 ,
     n57253 , n57254 , n57255 , n57256 , n57257 , n57258 , n57259 , n57260 , n57261 , n57262 ,
     n57263 , n57264 , n57265 , n57266 , n57267 , n57268 , n57269 , n57270 , n57271 , n57272 ,
     n57273 , n57274 , n57275 , n57276 , n57277 , n57278 , n57279 , n57280 , n57281 , n57282 ,
     n57283 , n57284 , n57285 , n57286 , n57287 , n57288 , n57289 , n57290 , n57291 , n57292 ,
     n57293 , n57294 , n57295 , n57296 , n57297 , n57298 , n57299 , n57300 , n57301 , n57302 ,
     n57303 , n57304 , n57305 , n57306 , n57307 , n57308 , n57309 , n57310 , n57311 , n57312 ,
     n57313 , n57314 , n57315 , n57316 , n57317 , n57318 , n57319 , n57320 , n57321 , n57322 ,
     n57323 , n57324 , n57325 , n57326 , n57327 , n57328 , n57329 , n57330 , n57331 , n57332 ,
     n57333 , n57334 , n57335 , n57336 , n57337 , n57338 , n57339 , n57340 , n57341 , n57342 ,
     n57343 , n57344 , n57345 , n57346 , n57347 , n57348 , n57349 , n57350 , n57351 , n57352 ,
     n57353 , n57354 , n57355 , n57356 , n57357 , n57358 , n57359 , n57360 , n57361 , n57362 ,
     n57363 , n57364 , n57365 , n57366 , n57367 , n57368 , n57369 , n57370 , n57371 , n57372 ,
     n57373 , n57374 , n57375 , n57376 , n57377 , n57378 , n57379 , n57380 , n57381 , n57382 ,
     n57383 , n57384 , n57385 , n57386 , n57387 , n57388 , n57389 , n57390 , n57391 , n57392 ,
     n57393 , n57394 , n57395 , n57396 , n57397 , n57398 , n57399 , n57400 , n57401 , n57402 ,
     n57403 , n57404 , n57405 , n57406 , n57407 , n57408 , n57409 , n57410 , n57411 , n57412 ,
     n57413 , n57414 , n57415 , n57416 , n57417 , n57418 , n57419 , n57420 , n57421 , n57422 ,
     n57423 , n57424 , n57425 , n57426 , n57427 , n57428 , n57429 , n57430 , n57431 , n57432 ,
     n57433 , n57434 , n57435 , n57436 , n57437 , n57438 , n57439 , n57440 , n57441 , n57442 ,
     n57443 , n57444 , n57445 , n57446 , n57447 , n57448 , n57449 , n57450 , n57451 , n57452 ,
     n57453 , n57454 , n57455 , n57456 , n57457 , n57458 , n57459 , n57460 , n57461 , n57462 ,
     n57463 , n57464 , n57465 , n57466 , n57467 , n57468 , n57469 , n57470 , n57471 , n57472 ,
     n57473 , n57474 , n57475 , n57476 , n57477 , n57478 , n57479 , n57480 , n57481 , n57482 ,
     n57483 , n57484 , n57485 , n57486 , n57487 , n57488 , n57489 , n57490 , n57491 , n57492 ,
     n57493 , n57494 , n57495 , n57496 , n57497 , n57498 , n57499 , n57500 , n57501 , n57502 ,
     n57503 , n57504 , n57505 , n57506 , n57507 , n57508 , n57509 , n57510 , n57511 , n57512 ,
     n57513 , n57514 , n57515 , n57516 , n57517 , n57518 , n57519 , n57520 , n57521 , n57522 ,
     n57523 , n57524 , n57525 , n57526 , n57527 , n57528 , n57529 , n57530 , n57531 , n57532 ,
     n57533 , n57534 , n57535 , n57536 , n57537 , n57538 , n57539 , n57540 , n57541 , n57542 ,
     n57543 , n57544 , n57545 , n57546 , n57547 , n57548 , n57549 , n57550 , n57551 , n57552 ,
     n57553 , n57554 , n57555 , n57556 , n57557 , n57558 , n57559 , n57560 , n57561 , n57562 ,
     n57563 , n57564 , n57565 , n57566 , n57567 , n57568 , n57569 , n57570 , n57571 , n57572 ,
     n57573 , n57574 , n57575 , n57576 , n57577 , n57578 , n57579 , n57580 , n57581 , n57582 ,
     n57583 , n57584 , n57585 , n57586 , n57587 , n57588 , n57589 , n57590 , n57591 , n57592 ,
     n57593 , n57594 , n57595 , n57596 , n57597 , n57598 , n57599 , n57600 , n57601 , n57602 ,
     n57603 , n57604 , n57605 , n57606 , n57607 , n57608 , n57609 , n57610 , n57611 , n57612 ,
     n57613 , n57614 , n57615 , n57616 , n57617 , n57618 , n57619 , n57620 , n57621 , n57622 ,
     n57623 , n57624 , n57625 , n57626 , n57627 , n57628 , n57629 , n57630 , n57631 , n57632 ,
     n57633 , n57634 , n57635 , n57636 , n57637 , n57638 , n57639 , n57640 , n57641 , n57642 ,
     n57643 , n57644 , n57645 , n57646 , n57647 , n57648 , n57649 , n57650 , n57651 , n57652 ,
     n57653 , n57654 , n57655 , n57656 , n57657 , n57658 , n57659 , n57660 , n57661 , n57662 ,
     n57663 , n57664 , n57665 , n57666 , n57667 , n57668 , n57669 , n57670 , n57671 , n57672 ,
     n57673 , n57674 , n57675 , n57676 , n57677 , n57678 , n57679 , n57680 , n57681 , n57682 ,
     n57683 , n57684 , n57685 , n57686 , n57687 , n57688 , n57689 , n57690 , n57691 , n57692 ,
     n57693 , n57694 , n57695 , n57696 , n57697 , n57698 , n57699 , n57700 , n57701 , n57702 ,
     n57703 , n57704 , n57705 , n57706 , n57707 , n57708 , n57709 , n57710 , n57711 , n57712 ,
     n57713 , n57714 , n57715 , n57716 , n57717 , n57718 , n57719 , n57720 , n57721 , n57722 ,
     n57723 , n57724 , n57725 , n57726 , n57727 , n57728 , n57729 , n57730 , n57731 , n57732 ,
     n57733 , n57734 , n57735 , n57736 , n57737 , n57738 , n57739 , n57740 , n57741 , n57742 ,
     n57743 , n57744 , n57745 , n57746 , n57747 , n57748 , n57749 , n57750 , n57751 , n57752 ,
     n57753 , n57754 , n57755 , n57756 , n57757 , n57758 , n57759 , n57760 , n57761 , n57762 ,
     n57763 , n57764 , n57765 , n57766 , n57767 , n57768 , n57769 , n57770 , n57771 , n57772 ,
     n57773 , n57774 , n57775 , n57776 , n57777 , n57778 , n57779 , n57780 , n57781 , n57782 ,
     n57783 , n57784 , n57785 , n57786 , n57787 , n57788 , n57789 , n57790 , n57791 , n57792 ,
     n57793 , n57794 , n57795 , n57796 , n57797 , n57798 , n57799 , n57800 , n57801 , n57802 ,
     n57803 , n57804 , n57805 , n57806 , n57807 , n57808 , n57809 , n57810 , n57811 , n57812 ,
     n57813 , n57814 , n57815 , n57816 , n57817 , n57818 , n57819 , n57820 , n57821 , n57822 ,
     n57823 , n57824 , n57825 , n57826 , n57827 , n57828 , n57829 , n57830 , n57831 , n57832 ,
     n57833 , n57834 , n57835 , n57836 , n57837 , n57838 , n57839 , n57840 , n57841 , n57842 ,
     n57843 , n57844 , n57845 , n57846 , n57847 , n57848 , n57849 , n57850 , n57851 , n57852 ,
     n57853 , n57854 , n57855 , n57856 , n57857 , n57858 , n57859 , n57860 , n57861 , n57862 ,
     n57863 , n57864 , n57865 , n57866 , n57867 , n57868 , n57869 , n57870 , n57871 , n57872 ,
     n57873 , n57874 , n57875 , n57876 , n57877 , n57878 , n57879 , n57880 , n57881 , n57882 ,
     n57883 , n57884 , n57885 , n57886 , n57887 , n57888 , n57889 , n57890 , n57891 , n57892 ,
     n57893 , n57894 , n57895 , n57896 , n57897 , n57898 , n57899 , n57900 , n57901 , n57902 ,
     n57903 , n57904 , n57905 , n57906 , n57907 , n57908 , n57909 , n57910 , n57911 , n57912 ,
     n57913 , n57914 , n57915 , n57916 , n57917 , n57918 , n57919 , n57920 , n57921 , n57922 ,
     n57923 , n57924 , n57925 , n57926 , n57927 , n57928 , n57929 , n57930 , n57931 , n57932 ,
     n57933 , n57934 , n57935 , n57936 , n57937 , n57938 , n57939 , n57940 , n57941 , n57942 ,
     n57943 , n57944 , n57945 , n57946 , n57947 , n57948 , n57949 , n57950 , n57951 , n57952 ,
     n57953 , n57954 , n57955 , n57956 , n57957 , n57958 , n57959 , n57960 , n57961 , n57962 ,
     n57963 , n57964 , n57965 , n57966 , n57967 , n57968 , n57969 , n57970 , n57971 , n57972 ,
     n57973 , n57974 , n57975 , n57976 , n57977 , n57978 , n57979 , n57980 , n57981 , n57982 ,
     n57983 , n57984 , n57985 , n57986 , n57987 , n57988 , n57989 , n57990 , n57991 , n57992 ,
     n57993 , n57994 , n57995 , n57996 , n57997 , n57998 , n57999 , n58000 , n58001 , n58002 ,
     n58003 , n58004 , n58005 , n58006 , n58007 , n58008 , n58009 , n58010 , n58011 , n58012 ,
     n58013 , n58014 , n58015 , n58016 , n58017 , n58018 , n58019 , n58020 , n58021 , n58022 ,
     n58023 , n58024 , n58025 , n58026 , n58027 , n58028 , n58029 , n58030 , n58031 , n58032 ,
     n58033 , n58034 , n58035 , n58036 , n58037 , n58038 , n58039 , n58040 , n58041 , n58042 ,
     n58043 , n58044 , n58045 , n58046 , n58047 , n58048 , n58049 , n58050 , n58051 , n58052 ,
     n58053 , n58054 , n58055 , n58056 , n58057 , n58058 , n58059 , n58060 , n58061 , n58062 ,
     n58063 , n58064 , n58065 , n58066 , n58067 , n58068 , n58069 , n58070 , n58071 , n58072 ,
     n58073 , n58074 , n58075 , n58076 , n58077 , n58078 , n58079 , n58080 , n58081 , n58082 ,
     n58083 , n58084 , n58085 , n58086 , n58087 , n58088 , n58089 , n58090 , n58091 , n58092 ,
     n58093 , n58094 , n58095 , n58096 , n58097 , n58098 , n58099 , n58100 , n58101 , n58102 ,
     n58103 , n58104 , n58105 , n58106 , n58107 , n58108 , n58109 , n58110 , n58111 , n58112 ,
     n58113 , n58114 , n58115 , n58116 , n58117 , n58118 , n58119 , n58120 , n58121 , n58122 ,
     n58123 , n58124 , n58125 , n58126 , n58127 , n58128 , n58129 , n58130 , n58131 , n58132 ,
     n58133 , n58134 , n58135 , n58136 , n58137 , n58138 , n58139 , n58140 , n58141 , n58142 ,
     n58143 , n58144 , n58145 , n58146 , n58147 , n58148 , n58149 , n58150 , n58151 , n58152 ,
     n58153 , n58154 , n58155 , n58156 , n58157 , n58158 , n58159 , n58160 , n58161 , n58162 ,
     n58163 , n58164 , n58165 , n58166 , n58167 , n58168 , n58169 , n58170 , n58171 , n58172 ,
     n58173 , n58174 , n58175 , n58176 , n58177 , n58178 , n58179 , n58180 , n58181 , n58182 ,
     n58183 , n58184 , n58185 , n58186 , n58187 , n58188 , n58189 , n58190 , n58191 , n58192 ,
     n58193 , n58194 , n58195 , n58196 , n58197 , n58198 , n58199 , n58200 , n58201 , n58202 ,
     n58203 , n58204 , n58205 , n58206 , n58207 , n58208 , n58209 , n58210 , n58211 , n58212 ,
     n58213 , n58214 , n58215 , n58216 , n58217 , n58218 , n58219 , n58220 , n58221 , n58222 ,
     n58223 , n58224 , n58225 , n58226 , n58227 , n58228 , n58229 , n58230 , n58231 , n58232 ,
     n58233 , n58234 , n58235 , n58236 , n58237 , n58238 , n58239 , n58240 , n58241 , n58242 ,
     n58243 , n58244 , n58245 , n58246 , n58247 , n58248 , n58249 , n58250 , n58251 , n58252 ,
     n58253 , n58254 , n58255 , n58256 , n58257 , n58258 , n58259 , n58260 , n58261 , n58262 ,
     n58263 , n58264 , n58265 , n58266 , n58267 , n58268 , n58269 , n58270 , n58271 , n58272 ,
     n58273 , n58274 , n58275 , n58276 , n58277 , n58278 , n58279 , n58280 , n58281 , n58282 ,
     n58283 , n58284 , n58285 , n58286 , n58287 , n58288 , n58289 , n58290 , n58291 , n58292 ,
     n58293 , n58294 , n58295 , n58296 , n58297 , n58298 , n58299 , n58300 , n58301 , n58302 ,
     n58303 , n58304 , n58305 , n58306 , n58307 , n58308 , n58309 , n58310 , n58311 , n58312 ,
     n58313 , n58314 , n58315 , n58316 , n58317 , n58318 , n58319 , n58320 , n58321 , n58322 ,
     n58323 , n58324 , n58325 , n58326 , n58327 , n58328 , n58329 , n58330 , n58331 , n58332 ,
     n58333 , n58334 , n58335 , n58336 , n58337 , n58338 , n58339 , n58340 , n58341 , n58342 ,
     n58343 , n58344 , n58345 , n58346 , n58347 , n58348 , n58349 , n58350 , n58351 , n58352 ,
     n58353 , n58354 , n58355 , n58356 , n58357 , n58358 , n58359 , n58360 , n58361 , n58362 ,
     n58363 , n58364 , n58365 , n58366 , n58367 , n58368 , n58369 , n58370 , n58371 , n58372 ,
     n58373 , n58374 , n58375 , n58376 , n58377 , n58378 , n58379 , n58380 , n58381 , n58382 ,
     n58383 , n58384 , n58385 , n58386 , n58387 , n58388 , n58389 , n58390 , n58391 , n58392 ,
     n58393 , n58394 , n58395 , n58396 , n58397 , n58398 , n58399 , n58400 , n58401 , n58402 ,
     n58403 , n58404 , n58405 , n58406 , n58407 , n58408 , n58409 , n58410 , n58411 , n58412 ,
     n58413 , n58414 , n58415 , n58416 , n58417 , n58418 , n58419 , n58420 , n58421 , n58422 ,
     n58423 , n58424 , n58425 , n58426 , n58427 , n58428 , n58429 , n58430 , n58431 , n58432 ,
     n58433 , n58434 , n58435 , n58436 , n58437 , n58438 , n58439 , n58440 , n58441 , n58442 ,
     n58443 , n58444 , n58445 , n58446 , n58447 , n58448 , n58449 , n58450 , n58451 , n58452 ,
     n58453 , n58454 , n58455 , n58456 , n58457 , n58458 , n58459 , n58460 , n58461 , n58462 ,
     n58463 , n58464 , n58465 , n58466 , n58467 , n58468 , n58469 , n58470 , n58471 , n58472 ,
     n58473 , n58474 , n58475 , n58476 , n58477 , n58478 , n58479 , n58480 , n58481 , n58482 ,
     n58483 , n58484 , n58485 , n58486 , n58487 , n58488 , n58489 , n58490 , n58491 , n58492 ,
     n58493 , n58494 , n58495 , n58496 , n58497 , n58498 , n58499 , n58500 , n58501 , n58502 ,
     n58503 , n58504 , n58505 , n58506 , n58507 , n58508 , n58509 , n58510 , n58511 , n58512 ,
     n58513 , n58514 , n58515 , n58516 , n58517 , n58518 , n58519 , n58520 , n58521 , n58522 ,
     n58523 , n58524 , n58525 , n58526 , n58527 , n58528 , n58529 , n58530 , n58531 , n58532 ,
     n58533 , n58534 , n58535 , n58536 , n58537 , n58538 , n58539 , n58540 , n58541 , n58542 ,
     n58543 , n58544 , n58545 , n58546 , n58547 , n58548 , n58549 , n58550 , n58551 , n58552 ,
     n58553 , n58554 , n58555 , n58556 , n58557 , n58558 , n58559 , n58560 , n58561 , n58562 ,
     n58563 , n58564 , n58565 , n58566 , n58567 , n58568 , n58569 , n58570 , n58571 , n58572 ,
     n58573 , n58574 , n58575 , n58576 , n58577 , n58578 , n58579 , n58580 , n58581 , n58582 ,
     n58583 , n58584 , n58585 , n58586 , n58587 , n58588 , n58589 , n58590 , n58591 , n58592 ,
     n58593 , n58594 , n58595 , n58596 , n58597 , n58598 , n58599 , n58600 , n58601 , n58602 ,
     n58603 , n58604 , n58605 , n58606 , n58607 , n58608 , n58609 , n58610 , n58611 , n58612 ,
     n58613 , n58614 , n58615 , n58616 , n58617 , n58618 , n58619 , n58620 , n58621 , n58622 ,
     n58623 , n58624 , n58625 , n58626 , n58627 , n58628 , n58629 , n58630 , n58631 , n58632 ,
     n58633 , n58634 , n58635 , n58636 , n58637 , n58638 , n58639 , n58640 , n58641 , n58642 ,
     n58643 , n58644 , n58645 , n58646 , n58647 , n58648 , n58649 , n58650 , n58651 , n58652 ,
     n58653 , n58654 , n58655 , n58656 , n58657 , n58658 , n58659 , n58660 , n58661 , n58662 ,
     n58663 , n58664 , n58665 , n58666 , n58667 , n58668 , n58669 , n58670 , n58671 , n58672 ,
     n58673 , n58674 , n58675 , n58676 , n58677 , n58678 , n58679 , n58680 , n58681 , n58682 ,
     n58683 , n58684 , n58685 , n58686 , n58687 , n58688 , n58689 , n58690 , n58691 , n58692 ,
     n58693 , n58694 , n58695 , n58696 , n58697 , n58698 , n58699 , n58700 , n58701 , n58702 ,
     n58703 , n58704 , n58705 , n58706 , n58707 , n58708 , n58709 , n58710 , n58711 , n58712 ,
     n58713 , n58714 , n58715 , n58716 , n58717 , n58718 , n58719 , n58720 , n58721 , n58722 ,
     n58723 , n58724 , n58725 , n58726 , n58727 , n58728 , n58729 , n58730 , n58731 , n58732 ,
     n58733 , n58734 , n58735 , n58736 , n58737 , n58738 , n58739 , n58740 , n58741 , n58742 ,
     n58743 , n58744 , n58745 , n58746 , n58747 , n58748 , n58749 , n58750 , n58751 , n58752 ,
     n58753 , n58754 , n58755 , n58756 , n58757 , n58758 , n58759 , n58760 , n58761 , n58762 ,
     n58763 , n58764 , n58765 , n58766 , n58767 , n58768 , n58769 , n58770 , n58771 , n58772 ,
     n58773 , n58774 , n58775 , n58776 , n58777 , n58778 , n58779 , n58780 , n58781 , n58782 ,
     n58783 , n58784 , n58785 , n58786 , n58787 , n58788 , n58789 , n58790 , n58791 , n58792 ,
     n58793 , n58794 , n58795 , n58796 , n58797 , n58798 , n58799 , n58800 , n58801 , n58802 ,
     n58803 , n58804 , n58805 , n58806 , n58807 , n58808 , n58809 , n58810 , n58811 , n58812 ,
     n58813 , n58814 , n58815 , n58816 , n58817 , n58818 , n58819 , n58820 , n58821 , n58822 ,
     n58823 , n58824 , n58825 , n58826 , n58827 , n58828 , n58829 , n58830 , n58831 , n58832 ,
     n58833 , n58834 , n58835 , n58836 , n58837 , n58838 , n58839 , n58840 , n58841 , n58842 ,
     n58843 , n58844 , n58845 , n58846 , n58847 , n58848 , n58849 , n58850 , n58851 , n58852 ,
     n58853 , n58854 , n58855 , n58856 , n58857 , n58858 , n58859 , n58860 , n58861 , n58862 ,
     n58863 , n58864 , n58865 , n58866 , n58867 , n58868 , n58869 , n58870 , n58871 , n58872 ,
     n58873 , n58874 , n58875 , n58876 , n58877 , n58878 , n58879 , n58880 , n58881 , n58882 ,
     n58883 , n58884 , n58885 , n58886 , n58887 , n58888 , n58889 , n58890 , n58891 , n58892 ,
     n58893 , n58894 , n58895 , n58896 , n58897 , n58898 , n58899 , n58900 , n58901 , n58902 ,
     n58903 , n58904 , n58905 , n58906 , n58907 , n58908 , n58909 , n58910 , n58911 , n58912 ,
     n58913 , n58914 , n58915 , n58916 , n58917 , n58918 , n58919 , n58920 , n58921 , n58922 ,
     n58923 , n58924 , n58925 , n58926 , n58927 , n58928 , n58929 , n58930 , n58931 , n58932 ,
     n58933 , n58934 , n58935 , n58936 , n58937 , n58938 , n58939 , n58940 , n58941 , n58942 ,
     n58943 , n58944 , n58945 , n58946 , n58947 , n58948 , n58949 , n58950 , n58951 , n58952 ,
     n58953 , n58954 , n58955 , n58956 , n58957 , n58958 , n58959 , n58960 , n58961 , n58962 ,
     n58963 , n58964 , n58965 , n58966 , n58967 , n58968 , n58969 , n58970 , n58971 , n58972 ,
     n58973 , n58974 , n58975 , n58976 , n58977 , n58978 , n58979 , n58980 , n58981 , n58982 ,
     n58983 , n58984 , n58985 , n58986 , n58987 , n58988 , n58989 , n58990 , n58991 , n58992 ,
     n58993 , n58994 , n58995 , n58996 , n58997 , n58998 , n58999 , n59000 , n59001 , n59002 ,
     n59003 , n59004 , n59005 , n59006 , n59007 , n59008 , n59009 , n59010 , n59011 , n59012 ,
     n59013 , n59014 , n59015 , n59016 , n59017 , n59018 , n59019 , n59020 , n59021 , n59022 ,
     n59023 , n59024 , n59025 , n59026 , n59027 , n59028 , n59029 , n59030 , n59031 , n59032 ,
     n59033 , n59034 , n59035 , n59036 , n59037 , n59038 , n59039 , n59040 , n59041 , n59042 ,
     n59043 , n59044 , n59045 , n59046 , n59047 , n59048 , n59049 , n59050 , n59051 , n59052 ,
     n59053 , n59054 , n59055 , n59056 , n59057 , n59058 , n59059 , n59060 , n59061 , n59062 ,
     n59063 , n59064 , n59065 , n59066 , n59067 , n59068 , n59069 , n59070 , n59071 , n59072 ,
     n59073 , n59074 , n59075 , n59076 , n59077 , n59078 , n59079 , n59080 , n59081 , n59082 ,
     n59083 , n59084 , n59085 , n59086 , n59087 , n59088 , n59089 , n59090 , n59091 , n59092 ,
     n59093 , n59094 , n59095 , n59096 , n59097 , n59098 , n59099 , n59100 , n59101 , n59102 ,
     n59103 , n59104 , n59105 , n59106 , n59107 , n59108 , n59109 , n59110 , n59111 , n59112 ,
     n59113 , n59114 , n59115 , n59116 , n59117 , n59118 , n59119 , n59120 , n59121 , n59122 ,
     n59123 , n59124 , n59125 , n59126 , n59127 , n59128 , n59129 , n59130 , n59131 , n59132 ,
     n59133 , n59134 , n59135 , n59136 , n59137 , n59138 , n59139 , n59140 , n59141 , n59142 ,
     n59143 , n59144 , n59145 , n59146 , n59147 , n59148 , n59149 , n59150 , n59151 , n59152 ,
     n59153 , n59154 , n59155 , n59156 , n59157 , n59158 , n59159 , n59160 , n59161 , n59162 ,
     n59163 , n59164 , n59165 , n59166 , n59167 , n59168 , n59169 , n59170 , n59171 , n59172 ,
     n59173 , n59174 , n59175 , n59176 , n59177 , n59178 , n59179 , n59180 , n59181 , n59182 ,
     n59183 , n59184 , n59185 , n59186 , n59187 , n59188 , n59189 , n59190 , n59191 , n59192 ,
     n59193 , n59194 , n59195 , n59196 , n59197 , n59198 , n59199 , n59200 , n59201 , n59202 ,
     n59203 , n59204 , n59205 , n59206 , n59207 , n59208 , n59209 , n59210 , n59211 , n59212 ,
     n59213 , n59214 , n59215 , n59216 , n59217 , n59218 , n59219 , n59220 , n59221 , n59222 ,
     n59223 , n59224 , n59225 , n59226 , n59227 , n59228 , n59229 , n59230 , n59231 , n59232 ,
     n59233 , n59234 , n59235 , n59236 , n59237 , n59238 , n59239 , n59240 , n59241 , n59242 ,
     n59243 , n59244 , n59245 , n59246 , n59247 , n59248 , n59249 , n59250 , n59251 , n59252 ,
     n59253 , n59254 , n59255 , n59256 , n59257 , n59258 , n59259 , n59260 , n59261 , n59262 ,
     n59263 , n59264 , n59265 , n59266 , n59267 , n59268 , n59269 , n59270 , n59271 , n59272 ,
     n59273 , n59274 , n59275 , n59276 , n59277 , n59278 , n59279 , n59280 , n59281 , n59282 ,
     n59283 , n59284 , n59285 , n59286 , n59287 , n59288 , n59289 , n59290 , n59291 , n59292 ,
     n59293 , n59294 , n59295 , n59296 , n59297 , n59298 , n59299 , n59300 , n59301 , n59302 ,
     n59303 , n59304 , n59305 , n59306 , n59307 , n59308 , n59309 , n59310 , n59311 , n59312 ,
     n59313 , n59314 , n59315 , n59316 , n59317 , n59318 , n59319 , n59320 , n59321 , n59322 ,
     n59323 , n59324 , n59325 , n59326 , n59327 , n59328 , n59329 , n59330 , n59331 , n59332 ,
     n59333 , n59334 , n59335 , n59336 , n59337 , n59338 , n59339 , n59340 , n59341 , n59342 ,
     n59343 , n59344 , n59345 , n59346 , n59347 , n59348 , n59349 , n59350 , n59351 , n59352 ,
     n59353 , n59354 , n59355 , n59356 , n59357 , n59358 , n59359 , n59360 , n59361 , n59362 ,
     n59363 , n59364 , n59365 , n59366 , n59367 , n59368 , n59369 , n59370 , n59371 , n59372 ,
     n59373 , n59374 , n59375 , n59376 , n59377 , n59378 , n59379 , n59380 , n59381 , n59382 ,
     n59383 , n59384 , n59385 , n59386 , n59387 , n59388 , n59389 , n59390 , n59391 , n59392 ,
     n59393 , n59394 , n59395 , n59396 , n59397 , n59398 , n59399 , n59400 , n59401 , n59402 ,
     n59403 , n59404 , n59405 , n59406 , n59407 , n59408 , n59409 , n59410 , n59411 , n59412 ,
     n59413 , n59414 , n59415 , n59416 , n59417 , n59418 , n59419 , n59420 , n59421 , n59422 ,
     n59423 , n59424 , n59425 , n59426 , n59427 , n59428 , n59429 , n59430 , n59431 , n59432 ,
     n59433 , n59434 , n59435 , n59436 , n59437 , n59438 , n59439 , n59440 , n59441 , n59442 ,
     n59443 , n59444 , n59445 , n59446 , n59447 , n59448 , n59449 , n59450 , n59451 , n59452 ,
     n59453 , n59454 , n59455 , n59456 , n59457 , n59458 , n59459 , n59460 , n59461 , n59462 ,
     n59463 , n59464 , n59465 , n59466 , n59467 , n59468 , n59469 , n59470 , n59471 , n59472 ,
     n59473 , n59474 , n59475 , n59476 , n59477 , n59478 , n59479 , n59480 , n59481 , n59482 ,
     n59483 , n59484 , n59485 , n59486 , n59487 , n59488 , n59489 , n59490 , n59491 , n59492 ,
     n59493 , n59494 , n59495 , n59496 , n59497 , n59498 , n59499 , n59500 , n59501 , n59502 ,
     n59503 , n59504 , n59505 , n59506 , n59507 , n59508 , n59509 , n59510 , n59511 , n59512 ,
     n59513 , n59514 , n59515 , n59516 , n59517 , n59518 , n59519 , n59520 , n59521 , n59522 ,
     n59523 , n59524 , n59525 , n59526 , n59527 , n59528 , n59529 , n59530 , n59531 , n59532 ,
     n59533 , n59534 , n59535 , n59536 , n59537 , n59538 , n59539 , n59540 , n59541 , n59542 ,
     n59543 , n59544 , n59545 , n59546 , n59547 , n59548 , n59549 , n59550 , n59551 , n59552 ,
     n59553 , n59554 , n59555 , n59556 , n59557 , n59558 , n59559 , n59560 , n59561 , n59562 ,
     n59563 , n59564 , n59565 , n59566 , n59567 , n59568 , n59569 , n59570 , n59571 , n59572 ,
     n59573 , n59574 , n59575 , n59576 , n59577 , n59578 , n59579 , n59580 , n59581 , n59582 ,
     n59583 , n59584 , n59585 , n59586 , n59587 , n59588 , n59589 , n59590 , n59591 , n59592 ,
     n59593 , n59594 , n59595 , n59596 , n59597 , n59598 , n59599 , n59600 , n59601 , n59602 ,
     n59603 , n59604 , n59605 , n59606 , n59607 , n59608 , n59609 , n59610 , n59611 , n59612 ,
     n59613 , n59614 , n59615 , n59616 , n59617 , n59618 , n59619 , n59620 , n59621 , n59622 ,
     n59623 , n59624 , n59625 , n59626 , n59627 , n59628 , n59629 , n59630 , n59631 , n59632 ,
     n59633 , n59634 , n59635 , n59636 , n59637 , n59638 , n59639 , n59640 , n59641 , n59642 ,
     n59643 , n59644 , n59645 , n59646 , n59647 , n59648 , n59649 , n59650 , n59651 , n59652 ,
     n59653 , n59654 , n59655 , n59656 , n59657 , n59658 , n59659 , n59660 , n59661 , n59662 ,
     n59663 , n59664 , n59665 , n59666 , n59667 , n59668 , n59669 , n59670 , n59671 , n59672 ,
     n59673 , n59674 , n59675 , n59676 , n59677 , n59678 , n59679 , n59680 , n59681 , n59682 ,
     n59683 , n59684 , n59685 , n59686 , n59687 , n59688 , n59689 , n59690 , n59691 , n59692 ,
     n59693 , n59694 , n59695 , n59696 , n59697 , n59698 , n59699 , n59700 , n59701 , n59702 ,
     n59703 , n59704 , n59705 , n59706 , n59707 , n59708 , n59709 , n59710 , n59711 , n59712 ,
     n59713 , n59714 , n59715 , n59716 , n59717 , n59718 , n59719 , n59720 , n59721 , n59722 ,
     n59723 , n59724 , n59725 , n59726 , n59727 , n59728 , n59729 , n59730 , n59731 , n59732 ,
     n59733 , n59734 , n59735 , n59736 , n59737 , n59738 , n59739 , n59740 , n59741 , n59742 ,
     n59743 , n59744 , n59745 , n59746 , n59747 , n59748 , n59749 , n59750 , n59751 , n59752 ,
     n59753 , n59754 , n59755 , n59756 , n59757 , n59758 , n59759 , n59760 , n59761 , n59762 ,
     n59763 , n59764 , n59765 , n59766 , n59767 , n59768 , n59769 , n59770 , n59771 , n59772 ,
     n59773 , n59774 , n59775 , n59776 , n59777 , n59778 , n59779 , n59780 , n59781 , n59782 ,
     n59783 , n59784 , n59785 , n59786 , n59787 , n59788 , n59789 , n59790 , n59791 , n59792 ,
     n59793 , n59794 , n59795 , n59796 , n59797 , n59798 , n59799 , n59800 , n59801 , n59802 ,
     n59803 , n59804 , n59805 , n59806 , n59807 , n59808 , n59809 , n59810 , n59811 , n59812 ,
     n59813 , n59814 , n59815 , n59816 , n59817 , n59818 , n59819 , n59820 , n59821 , n59822 ,
     n59823 , n59824 , n59825 , n59826 , n59827 , n59828 , n59829 , n59830 , n59831 , n59832 ,
     n59833 , n59834 , n59835 , n59836 , n59837 , n59838 , n59839 , n59840 , n59841 , n59842 ,
     n59843 , n59844 , n59845 , n59846 , n59847 , n59848 , n59849 , n59850 , n59851 , n59852 ,
     n59853 , n59854 , n59855 , n59856 , n59857 , n59858 , n59859 , n59860 , n59861 , n59862 ,
     n59863 , n59864 , n59865 , n59866 , n59867 , n59868 , n59869 , n59870 , n59871 , n59872 ,
     n59873 , n59874 , n59875 , n59876 , n59877 , n59878 , n59879 , n59880 , n59881 , n59882 ,
     n59883 , n59884 , n59885 , n59886 , n59887 , n59888 , n59889 , n59890 , n59891 , n59892 ,
     n59893 , n59894 , n59895 , n59896 , n59897 , n59898 , n59899 , n59900 , n59901 , n59902 ,
     n59903 , n59904 , n59905 , n59906 , n59907 , n59908 , n59909 , n59910 , n59911 , n59912 ,
     n59913 , n59914 , n59915 , n59916 , n59917 , n59918 , n59919 , n59920 , n59921 , n59922 ,
     n59923 , n59924 , n59925 , n59926 , n59927 , n59928 , n59929 , n59930 , n59931 , n59932 ,
     n59933 , n59934 , n59935 , n59936 , n59937 , n59938 , n59939 , n59940 , n59941 , n59942 ,
     n59943 , n59944 , n59945 , n59946 , n59947 , n59948 , n59949 , n59950 , n59951 , n59952 ,
     n59953 , n59954 , n59955 , n59956 , n59957 , n59958 , n59959 , n59960 , n59961 , n59962 ,
     n59963 , n59964 , n59965 , n59966 , n59967 , n59968 , n59969 , n59970 , n59971 , n59972 ,
     n59973 , n59974 , n59975 , n59976 , n59977 , n59978 , n59979 , n59980 , n59981 , n59982 ,
     n59983 , n59984 , n59985 , n59986 , n59987 , n59988 , n59989 , n59990 , n59991 , n59992 ,
     n59993 , n59994 , n59995 , n59996 , n59997 , n59998 , n59999 , n60000 , n60001 , n60002 ,
     n60003 , n60004 , n60005 , n60006 , n60007 , n60008 , n60009 , n60010 , n60011 , n60012 ,
     n60013 , n60014 , n60015 , n60016 , n60017 , n60018 , n60019 , n60020 , n60021 , n60022 ,
     n60023 , n60024 , n60025 , n60026 , n60027 , n60028 , n60029 , n60030 , n60031 , n60032 ,
     n60033 , n60034 , n60035 , n60036 , n60037 , n60038 , n60039 , n60040 , n60041 , n60042 ,
     n60043 , n60044 , n60045 , n60046 , n60047 , n60048 , n60049 , n60050 , n60051 , n60052 ,
     n60053 , n60054 , n60055 , n60056 , n60057 , n60058 , n60059 , n60060 , n60061 , n60062 ,
     n60063 , n60064 , n60065 , n60066 , n60067 , n60068 , n60069 , n60070 , n60071 , n60072 ,
     n60073 , n60074 , n60075 , n60076 , n60077 , n60078 , n60079 , n60080 , n60081 , n60082 ,
     n60083 , n60084 , n60085 , n60086 , n60087 , n60088 , n60089 , n60090 , n60091 , n60092 ,
     n60093 , n60094 , n60095 , n60096 , n60097 , n60098 , n60099 , n60100 , n60101 , n60102 ,
     n60103 , n60104 , n60105 , n60106 , n60107 , n60108 , n60109 , n60110 , n60111 , n60112 ,
     n60113 , n60114 , n60115 , n60116 , n60117 , n60118 , n60119 , n60120 , n60121 , n60122 ,
     n60123 , n60124 , n60125 , n60126 , n60127 , n60128 , n60129 , n60130 , n60131 , n60132 ,
     n60133 , n60134 , n60135 , n60136 , n60137 , n60138 , n60139 , n60140 , n60141 , n60142 ,
     n60143 , n60144 , n60145 , n60146 , n60147 , n60148 , n60149 , n60150 , n60151 , n60152 ,
     n60153 , n60154 , n60155 , n60156 , n60157 , n60158 , n60159 , n60160 , n60161 , n60162 ,
     n60163 , n60164 , n60165 , n60166 , n60167 , n60168 , n60169 , n60170 , n60171 , n60172 ,
     n60173 , n60174 , n60175 , n60176 , n60177 , n60178 , n60179 , n60180 , n60181 , n60182 ,
     n60183 , n60184 , n60185 , n60186 , n60187 , n60188 , n60189 , n60190 , n60191 , n60192 ,
     n60193 , n60194 , n60195 , n60196 , n60197 , n60198 , n60199 , n60200 , n60201 , n60202 ,
     n60203 , n60204 , n60205 , n60206 , n60207 , n60208 , n60209 , n60210 , n60211 , n60212 ,
     n60213 , n60214 , n60215 , n60216 , n60217 , n60218 , n60219 , n60220 , n60221 , n60222 ,
     n60223 , n60224 , n60225 , n60226 , n60227 , n60228 , n60229 , n60230 , n60231 , n60232 ,
     n60233 , n60234 , n60235 , n60236 , n60237 , n60238 , n60239 , n60240 , n60241 , n60242 ,
     n60243 , n60244 , n60245 , n60246 , n60247 , n60248 , n60249 , n60250 , n60251 , n60252 ,
     n60253 , n60254 , n60255 , n60256 , n60257 , n60258 , n60259 , n60260 , n60261 , n60262 ,
     n60263 , n60264 , n60265 , n60266 , n60267 , n60268 , n60269 , n60270 , n60271 , n60272 ,
     n60273 , n60274 , n60275 , n60276 , n60277 , n60278 , n60279 , n60280 , n60281 , n60282 ,
     n60283 , n60284 , n60285 , n60286 , n60287 , n60288 , n60289 , n60290 , n60291 , n60292 ,
     n60293 , n60294 , n60295 , n60296 , n60297 , n60298 , n60299 , n60300 , n60301 , n60302 ,
     n60303 , n60304 , n60305 , n60306 , n60307 , n60308 , n60309 , n60310 , n60311 , n60312 ,
     n60313 , n60314 , n60315 , n60316 , n60317 , n60318 , n60319 , n60320 , n60321 , n60322 ,
     n60323 , n60324 , n60325 , n60326 , n60327 , n60328 , n60329 , n60330 , n60331 , n60332 ,
     n60333 , n60334 , n60335 , n60336 , n60337 , n60338 , n60339 , n60340 , n60341 , n60342 ,
     n60343 , n60344 , n60345 , n60346 , n60347 , n60348 , n60349 , n60350 , n60351 , n60352 ,
     n60353 , n60354 , n60355 , n60356 , n60357 , n60358 , n60359 , n60360 , n60361 , n60362 ,
     n60363 , n60364 , n60365 , n60366 , n60367 , n60368 , n60369 , n60370 , n60371 , n60372 ,
     n60373 , n60374 , n60375 , n60376 , n60377 , n60378 , n60379 , n60380 , n60381 , n60382 ,
     n60383 , n60384 , n60385 , n60386 , n60387 , n60388 , n60389 , n60390 , n60391 , n60392 ,
     n60393 , n60394 , n60395 , n60396 , n60397 , n60398 , n60399 , n60400 , n60401 , n60402 ,
     n60403 , n60404 , n60405 , n60406 , n60407 , n60408 , n60409 , n60410 , n60411 , n60412 ,
     n60413 , n60414 , n60415 , n60416 , n60417 , n60418 , n60419 , n60420 , n60421 , n60422 ,
     n60423 , n60424 , n60425 , n60426 , n60427 , n60428 , n60429 , n60430 , n60431 , n60432 ,
     n60433 , n60434 , n60435 , n60436 , n60437 , n60438 , n60439 , n60440 , n60441 , n60442 ,
     n60443 , n60444 , n60445 , n60446 , n60447 , n60448 , n60449 , n60450 , n60451 , n60452 ,
     n60453 , n60454 , n60455 , n60456 , n60457 , n60458 , n60459 , n60460 , n60461 , n60462 ,
     n60463 , n60464 , n60465 , n60466 , n60467 , n60468 , n60469 , n60470 , n60471 , n60472 ,
     n60473 , n60474 , n60475 , n60476 , n60477 , n60478 , n60479 , n60480 , n60481 , n60482 ,
     n60483 , n60484 , n60485 , n60486 , n60487 , n60488 , n60489 , n60490 , n60491 , n60492 ,
     n60493 , n60494 , n60495 , n60496 , n60497 , n60498 , n60499 , n60500 , n60501 , n60502 ,
     n60503 , n60504 , n60505 , n60506 , n60507 , n60508 , n60509 , n60510 , n60511 , n60512 ,
     n60513 , n60514 , n60515 , n60516 , n60517 , n60518 , n60519 , n60520 , n60521 , n60522 ,
     n60523 , n60524 , n60525 , n60526 , n60527 , n60528 , n60529 , n60530 , n60531 , n60532 ,
     n60533 , n60534 , n60535 , n60536 , n60537 , n60538 , n60539 , n60540 , n60541 , n60542 ,
     n60543 , n60544 , n60545 , n60546 , n60547 , n60548 , n60549 , n60550 , n60551 , n60552 ,
     n60553 , n60554 , n60555 , n60556 , n60557 , n60558 , n60559 , n60560 , n60561 , n60562 ,
     n60563 , n60564 , n60565 , n60566 , n60567 , n60568 , n60569 , n60570 , n60571 , n60572 ,
     n60573 , n60574 , n60575 , n60576 , n60577 , n60578 , n60579 , n60580 , n60581 , n60582 ,
     n60583 , n60584 , n60585 , n60586 , n60587 , n60588 , n60589 , n60590 , n60591 , n60592 ,
     n60593 , n60594 , n60595 , n60596 , n60597 , n60598 , n60599 , n60600 , n60601 , n60602 ,
     n60603 , n60604 , n60605 , n60606 , n60607 , n60608 , n60609 , n60610 , n60611 , n60612 ,
     n60613 , n60614 , n60615 , n60616 , n60617 , n60618 , n60619 , n60620 , n60621 , n60622 ,
     n60623 , n60624 , n60625 , n60626 , n60627 , n60628 , n60629 , n60630 , n60631 , n60632 ,
     n60633 , n60634 , n60635 , n60636 , n60637 , n60638 , n60639 , n60640 , n60641 , n60642 ,
     n60643 , n60644 , n60645 , n60646 , n60647 , n60648 , n60649 , n60650 , n60651 , n60652 ,
     n60653 , n60654 , n60655 , n60656 , n60657 , n60658 , n60659 , n60660 , n60661 , n60662 ,
     n60663 , n60664 , n60665 , n60666 , n60667 , n60668 , n60669 , n60670 , n60671 , n60672 ,
     n60673 , n60674 , n60675 , n60676 , n60677 , n60678 , n60679 , n60680 , n60681 , n60682 ,
     n60683 , n60684 , n60685 , n60686 , n60687 , n60688 , n60689 , n60690 , n60691 , n60692 ,
     n60693 , n60694 , n60695 , n60696 , n60697 , n60698 , n60699 , n60700 , n60701 , n60702 ,
     n60703 , n60704 , n60705 , n60706 , n60707 , n60708 , n60709 , n60710 , n60711 , n60712 ,
     n60713 , n60714 , n60715 , n60716 , n60717 , n60718 , n60719 , n60720 , n60721 , n60722 ,
     n60723 , n60724 , n60725 , n60726 , n60727 , n60728 , n60729 , n60730 , n60731 , n60732 ,
     n60733 , n60734 , n60735 , n60736 , n60737 , n60738 , n60739 , n60740 , n60741 , n60742 ,
     n60743 , n60744 , n60745 , n60746 , n60747 , n60748 , n60749 , n60750 , n60751 , n60752 ,
     n60753 , n60754 , n60755 , n60756 , n60757 , n60758 , n60759 , n60760 , n60761 , n60762 ,
     n60763 , n60764 , n60765 , n60766 , n60767 , n60768 , n60769 , n60770 , n60771 , n60772 ,
     n60773 , n60774 , n60775 , n60776 , n60777 , n60778 , n60779 , n60780 , n60781 , n60782 ,
     n60783 , n60784 , n60785 , n60786 , n60787 , n60788 , n60789 , n60790 , n60791 , n60792 ,
     n60793 , n60794 , n60795 , n60796 , n60797 , n60798 , n60799 , n60800 , n60801 , n60802 ,
     n60803 , n60804 , n60805 , n60806 , n60807 , n60808 , n60809 , n60810 , n60811 , n60812 ,
     n60813 , n60814 , n60815 , n60816 , n60817 , n60818 , n60819 , n60820 , n60821 , n60822 ,
     n60823 , n60824 , n60825 , n60826 , n60827 , n60828 , n60829 , n60830 , n60831 , n60832 ,
     n60833 , n60834 , n60835 , n60836 , n60837 , n60838 , n60839 , n60840 , n60841 , n60842 ,
     n60843 , n60844 , n60845 , n60846 , n60847 , n60848 , n60849 , n60850 , n60851 , n60852 ,
     n60853 , n60854 , n60855 , n60856 , n60857 , n60858 , n60859 , n60860 , n60861 , n60862 ,
     n60863 , n60864 , n60865 , n60866 , n60867 , n60868 , n60869 , n60870 , n60871 , n60872 ,
     n60873 , n60874 , n60875 , n60876 , n60877 , n60878 , n60879 , n60880 , n60881 , n60882 ,
     n60883 , n60884 , n60885 , n60886 , n60887 , n60888 , n60889 , n60890 , n60891 , n60892 ,
     n60893 , n60894 , n60895 , n60896 , n60897 , n60898 , n60899 , n60900 , n60901 , n60902 ,
     n60903 , n60904 , n60905 , n60906 , n60907 , n60908 , n60909 , n60910 , n60911 , n60912 ,
     n60913 , n60914 , n60915 , n60916 , n60917 , n60918 , n60919 , n60920 , n60921 , n60922 ,
     n60923 , n60924 , n60925 , n60926 , n60927 , n60928 , n60929 , n60930 , n60931 , n60932 ,
     n60933 , n60934 , n60935 , n60936 , n60937 , n60938 , n60939 , n60940 , n60941 , n60942 ,
     n60943 , n60944 , n60945 , n60946 , n60947 , n60948 , n60949 , n60950 , n60951 , n60952 ,
     n60953 , n60954 , n60955 , n60956 , n60957 , n60958 , n60959 , n60960 , n60961 , n60962 ,
     n60963 , n60964 , n60965 , n60966 , n60967 , n60968 , n60969 , n60970 , n60971 , n60972 ,
     n60973 , n60974 , n60975 , n60976 , n60977 , n60978 , n60979 , n60980 , n60981 , n60982 ,
     n60983 , n60984 , n60985 , n60986 , n60987 , n60988 , n60989 , n60990 , n60991 , n60992 ,
     n60993 , n60994 , n60995 , n60996 , n60997 , n60998 , n60999 , n61000 , n61001 , n61002 ,
     n61003 , n61004 , n61005 , n61006 , n61007 , n61008 , n61009 , n61010 , n61011 , n61012 ,
     n61013 , n61014 , n61015 , n61016 , n61017 , n61018 , n61019 , n61020 , n61021 , n61022 ,
     n61023 , n61024 , n61025 , n61026 , n61027 , n61028 , n61029 , n61030 , n61031 , n61032 ,
     n61033 , n61034 , n61035 , n61036 , n61037 , n61038 , n61039 , n61040 , n61041 , n61042 ,
     n61043 , n61044 , n61045 , n61046 , n61047 , n61048 , n61049 , n61050 , n61051 , n61052 ,
     n61053 , n61054 , n61055 , n61056 , n61057 , n61058 , n61059 , n61060 , n61061 , n61062 ,
     n61063 , n61064 , n61065 , n61066 , n61067 , n61068 , n61069 , n61070 , n61071 , n61072 ,
     n61073 , n61074 , n61075 , n61076 , n61077 , n61078 , n61079 , n61080 , n61081 , n61082 ,
     n61083 , n61084 , n61085 , n61086 , n61087 , n61088 , n61089 , n61090 , n61091 , n61092 ,
     n61093 , n61094 , n61095 , n61096 , n61097 , n61098 , n61099 , n61100 , n61101 , n61102 ,
     n61103 , n61104 , n61105 , n61106 , n61107 , n61108 , n61109 , n61110 , n61111 , n61112 ,
     n61113 , n61114 , n61115 , n61116 , n61117 , n61118 , n61119 , n61120 , n61121 , n61122 ,
     n61123 , n61124 , n61125 , n61126 , n61127 , n61128 , n61129 , n61130 , n61131 , n61132 ,
     n61133 , n61134 , n61135 , n61136 , n61137 , n61138 , n61139 , n61140 , n61141 , n61142 ,
     n61143 , n61144 , n61145 , n61146 , n61147 , n61148 , n61149 , n61150 , n61151 , n61152 ,
     n61153 , n61154 , n61155 , n61156 , n61157 , n61158 , n61159 , n61160 , n61161 , n61162 ,
     n61163 , n61164 , n61165 , n61166 , n61167 , n61168 , n61169 , n61170 , n61171 , n61172 ,
     n61173 , n61174 , n61175 , n61176 , n61177 , n61178 , n61179 , n61180 , n61181 , n61182 ,
     n61183 , n61184 , n61185 , n61186 , n61187 , n61188 , n61189 , n61190 , n61191 , n61192 ,
     n61193 , n61194 , n61195 , n61196 , n61197 , n61198 , n61199 , n61200 , n61201 , n61202 ,
     n61203 , n61204 , n61205 , n61206 , n61207 , n61208 , n61209 , n61210 , n61211 , n61212 ,
     n61213 , n61214 , n61215 , n61216 , n61217 , n61218 , n61219 , n61220 , n61221 , n61222 ,
     n61223 , n61224 , n61225 , n61226 , n61227 , n61228 , n61229 , n61230 , n61231 , n61232 ,
     n61233 , n61234 , n61235 , n61236 , n61237 , n61238 , n61239 , n61240 , n61241 , n61242 ,
     n61243 , n61244 , n61245 , n61246 , n61247 , n61248 , n61249 , n61250 , n61251 , n61252 ,
     n61253 , n61254 , n61255 , n61256 , n61257 , n61258 , n61259 , n61260 , n61261 , n61262 ,
     n61263 , n61264 , n61265 , n61266 , n61267 , n61268 , n61269 , n61270 , n61271 , n61272 ,
     n61273 , n61274 , n61275 , n61276 , n61277 , n61278 , n61279 , n61280 , n61281 , n61282 ,
     n61283 , n61284 , n61285 , n61286 , n61287 , n61288 , n61289 , n61290 , n61291 , n61292 ,
     n61293 , n61294 , n61295 , n61296 , n61297 , n61298 , n61299 , n61300 , n61301 , n61302 ,
     n61303 , n61304 , n61305 , n61306 , n61307 , n61308 , n61309 , n61310 , n61311 , n61312 ,
     n61313 , n61314 , n61315 , n61316 , n61317 , n61318 , n61319 , n61320 , n61321 , n61322 ,
     n61323 , n61324 , n61325 , n61326 , n61327 , n61328 , n61329 , n61330 , n61331 , n61332 ,
     n61333 , n61334 , n61335 , n61336 , n61337 , n61338 , n61339 , n61340 , n61341 , n61342 ,
     n61343 , n61344 , n61345 , n61346 , n61347 , n61348 , n61349 , n61350 , n61351 , n61352 ,
     n61353 , n61354 , n61355 , n61356 , n61357 , n61358 , n61359 , n61360 , n61361 , n61362 ,
     n61363 , n61364 , n61365 , n61366 , n61367 , n61368 , n61369 , n61370 , n61371 , n61372 ,
     n61373 , n61374 , n61375 , n61376 , n61377 , n61378 , n61379 , n61380 , n61381 , n61382 ,
     n61383 , n61384 , n61385 , n61386 , n61387 , n61388 , n61389 , n61390 , n61391 , n61392 ,
     n61393 , n61394 , n61395 , n61396 , n61397 , n61398 , n61399 , n61400 , n61401 , n61402 ,
     n61403 , n61404 , n61405 , n61406 , n61407 , n61408 , n61409 , n61410 , n61411 , n61412 ,
     n61413 , n61414 , n61415 , n61416 , n61417 , n61418 , n61419 , n61420 , n61421 , n61422 ,
     n61423 , n61424 , n61425 , n61426 , n61427 , n61428 , n61429 , n61430 , n61431 , n61432 ,
     n61433 , n61434 , n61435 , n61436 , n61437 , n61438 , n61439 , n61440 , n61441 , n61442 ,
     n61443 , n61444 , n61445 , n61446 , n61447 , n61448 , n61449 , n61450 , n61451 , n61452 ,
     n61453 , n61454 , n61455 , n61456 , n61457 , n61458 , n61459 , n61460 , n61461 , n61462 ,
     n61463 , n61464 , n61465 , n61466 , n61467 , n61468 , n61469 , n61470 , n61471 , n61472 ,
     n61473 , n61474 , n61475 , n61476 , n61477 , n61478 , n61479 , n61480 , n61481 , n61482 ,
     n61483 , n61484 , n61485 , n61486 , n61487 , n61488 , n61489 , n61490 , n61491 , n61492 ,
     n61493 , n61494 , n61495 , n61496 , n61497 , n61498 , n61499 , n61500 , n61501 , n61502 ,
     n61503 , n61504 , n61505 , n61506 , n61507 , n61508 , n61509 , n61510 , n61511 , n61512 ,
     n61513 , n61514 , n61515 , n61516 , n61517 , n61518 , n61519 , n61520 , n61521 , n61522 ,
     n61523 , n61524 , n61525 , n61526 , n61527 , n61528 , n61529 , n61530 , n61531 , n61532 ,
     n61533 , n61534 , n61535 , n61536 , n61537 , n61538 , n61539 , n61540 , n61541 , n61542 ,
     n61543 , n61544 , n61545 , n61546 , n61547 , n61548 , n61549 , n61550 , n61551 , n61552 ,
     n61553 , n61554 , n61555 , n61556 , n61557 , n61558 , n61559 , n61560 , n61561 , n61562 ,
     n61563 , n61564 , n61565 , n61566 , n61567 , n61568 , n61569 , n61570 , n61571 , n61572 ,
     n61573 , n61574 , n61575 , n61576 , n61577 , n61578 , n61579 , n61580 , n61581 , n61582 ,
     n61583 , n61584 , n61585 , n61586 , n61587 , n61588 , n61589 , n61590 , n61591 , n61592 ,
     n61593 , n61594 , n61595 , n61596 , n61597 , n61598 , n61599 , n61600 , n61601 , n61602 ,
     n61603 , n61604 , n61605 , n61606 , n61607 , n61608 , n61609 , n61610 , n61611 , n61612 ,
     n61613 , n61614 , n61615 , n61616 , n61617 , n61618 , n61619 , n61620 , n61621 , n61622 ,
     n61623 , n61624 , n61625 , n61626 , n61627 , n61628 , n61629 , n61630 , n61631 , n61632 ,
     n61633 , n61634 , n61635 , n61636 , n61637 , n61638 , n61639 , n61640 , n61641 , n61642 ,
     n61643 , n61644 , n61645 , n61646 , n61647 , n61648 , n61649 , n61650 , n61651 , n61652 ,
     n61653 , n61654 , n61655 , n61656 , n61657 , n61658 , n61659 , n61660 , n61661 , n61662 ,
     n61663 , n61664 , n61665 , n61666 , n61667 , n61668 , n61669 , n61670 , n61671 , n61672 ,
     n61673 , n61674 , n61675 , n61676 , n61677 , n61678 , n61679 , n61680 , n61681 , n61682 ,
     n61683 , n61684 , n61685 , n61686 , n61687 , n61688 , n61689 , n61690 , n61691 , n61692 ,
     n61693 , n61694 , n61695 , n61696 , n61697 , n61698 , n61699 , n61700 , n61701 , n61702 ,
     n61703 , n61704 , n61705 , n61706 , n61707 , n61708 , n61709 , n61710 , n61711 , n61712 ,
     n61713 , n61714 , n61715 , n61716 , n61717 , n61718 , n61719 , n61720 , n61721 , n61722 ,
     n61723 , n61724 , n61725 , n61726 , n61727 , n61728 , n61729 , n61730 , n61731 , n61732 ,
     n61733 , n61734 , n61735 , n61736 , n61737 , n61738 , n61739 , n61740 , n61741 , n61742 ,
     n61743 , n61744 , n61745 , n61746 , n61747 , n61748 , n61749 , n61750 , n61751 , n61752 ,
     n61753 , n61754 , n61755 , n61756 , n61757 , n61758 , n61759 , n61760 , n61761 , n61762 ,
     n61763 , n61764 , n61765 , n61766 , n61767 , n61768 , n61769 , n61770 , n61771 , n61772 ,
     n61773 , n61774 , n61775 , n61776 , n61777 , n61778 , n61779 , n61780 , n61781 , n61782 ,
     n61783 , n61784 , n61785 , n61786 , n61787 , n61788 , n61789 , n61790 , n61791 , n61792 ,
     n61793 , n61794 , n61795 , n61796 , n61797 , n61798 , n61799 , n61800 , n61801 , n61802 ,
     n61803 , n61804 , n61805 , n61806 , n61807 , n61808 , n61809 , n61810 , n61811 , n61812 ,
     n61813 , n61814 , n61815 , n61816 , n61817 , n61818 , n61819 , n61820 , n61821 , n61822 ,
     n61823 , n61824 , n61825 , n61826 , n61827 , n61828 , n61829 , n61830 , n61831 , n61832 ,
     n61833 , n61834 , n61835 , n61836 , n61837 , n61838 , n61839 , n61840 , n61841 , n61842 ,
     n61843 , n61844 , n61845 , n61846 , n61847 , n61848 , n61849 , n61850 , n61851 , n61852 ,
     n61853 , n61854 , n61855 , n61856 , n61857 , n61858 , n61859 , n61860 , n61861 , n61862 ,
     n61863 , n61864 , n61865 , n61866 , n61867 , n61868 , n61869 , n61870 , n61871 , n61872 ,
     n61873 , n61874 , n61875 , n61876 , n61877 , n61878 , n61879 , n61880 , n61881 , n61882 ,
     n61883 , n61884 , n61885 , n61886 , n61887 , n61888 , n61889 , n61890 , n61891 , n61892 ,
     n61893 , n61894 , n61895 , n61896 , n61897 , n61898 , n61899 , n61900 , n61901 , n61902 ,
     n61903 , n61904 , n61905 , n61906 , n61907 , n61908 , n61909 , n61910 , n61911 , n61912 ,
     n61913 , n61914 , n61915 , n61916 , n61917 , n61918 , n61919 , n61920 , n61921 , n61922 ,
     n61923 , n61924 , n61925 , n61926 , n61927 , n61928 , n61929 , n61930 , n61931 , n61932 ,
     n61933 , n61934 , n61935 , n61936 , n61937 , n61938 , n61939 , n61940 , n61941 , n61942 ,
     n61943 , n61944 , n61945 , n61946 , n61947 , n61948 , n61949 , n61950 , n61951 , n61952 ,
     n61953 , n61954 , n61955 , n61956 , n61957 , n61958 , n61959 , n61960 , n61961 , n61962 ,
     n61963 , n61964 , n61965 , n61966 , n61967 , n61968 , n61969 , n61970 , n61971 , n61972 ,
     n61973 , n61974 , n61975 , n61976 , n61977 , n61978 , n61979 , n61980 , n61981 , n61982 ,
     n61983 , n61984 , n61985 , n61986 , n61987 , n61988 , n61989 , n61990 , n61991 , n61992 ,
     n61993 , n61994 , n61995 , n61996 , n61997 , n61998 , n61999 , n62000 , n62001 , n62002 ,
     n62003 , n62004 , n62005 , n62006 , n62007 , n62008 , n62009 , n62010 , n62011 , n62012 ,
     n62013 , n62014 , n62015 , n62016 , n62017 , n62018 , n62019 , n62020 , n62021 , n62022 ,
     n62023 , n62024 , n62025 , n62026 , n62027 , n62028 , n62029 , n62030 , n62031 , n62032 ,
     n62033 , n62034 , n62035 , n62036 , n62037 , n62038 , n62039 , n62040 , n62041 , n62042 ,
     n62043 , n62044 , n62045 , n62046 , n62047 , n62048 , n62049 , n62050 , n62051 , n62052 ,
     n62053 , n62054 , n62055 , n62056 , n62057 , n62058 , n62059 , n62060 , n62061 , n62062 ,
     n62063 , n62064 , n62065 , n62066 , n62067 , n62068 , n62069 , n62070 , n62071 , n62072 ,
     n62073 , n62074 , n62075 , n62076 , n62077 , n62078 , n62079 , n62080 , n62081 , n62082 ,
     n62083 , n62084 , n62085 , n62086 , n62087 , n62088 , n62089 , n62090 , n62091 , n62092 ,
     n62093 , n62094 , n62095 , n62096 , n62097 , n62098 , n62099 , n62100 , n62101 , n62102 ,
     n62103 , n62104 , n62105 , n62106 , n62107 , n62108 , n62109 , n62110 , n62111 , n62112 ,
     n62113 , n62114 , n62115 , n62116 , n62117 , n62118 , n62119 , n62120 , n62121 , n62122 ,
     n62123 , n62124 , n62125 , n62126 , n62127 , n62128 , n62129 , n62130 , n62131 , n62132 ,
     n62133 , n62134 , n62135 , n62136 , n62137 , n62138 , n62139 , n62140 , n62141 , n62142 ,
     n62143 , n62144 , n62145 , n62146 , n62147 , n62148 , n62149 , n62150 , n62151 , n62152 ,
     n62153 , n62154 , n62155 , n62156 , n62157 , n62158 , n62159 , n62160 , n62161 , n62162 ,
     n62163 , n62164 , n62165 , n62166 , n62167 , n62168 , n62169 , n62170 , n62171 , n62172 ,
     n62173 , n62174 , n62175 , n62176 , n62177 , n62178 , n62179 , n62180 , n62181 , n62182 ,
     n62183 , n62184 , n62185 , n62186 , n62187 , n62188 , n62189 , n62190 , n62191 , n62192 ,
     n62193 , n62194 , n62195 , n62196 , n62197 , n62198 , n62199 , n62200 , n62201 , n62202 ,
     n62203 , n62204 , n62205 , n62206 , n62207 , n62208 , n62209 , n62210 , n62211 , n62212 ,
     n62213 , n62214 , n62215 , n62216 , n62217 , n62218 , n62219 , n62220 , n62221 , n62222 ,
     n62223 , n62224 , n62225 , n62226 , n62227 , n62228 , n62229 , n62230 , n62231 , n62232 ,
     n62233 , n62234 , n62235 , n62236 , n62237 , n62238 , n62239 , n62240 , n62241 , n62242 ,
     n62243 , n62244 , n62245 , n62246 , n62247 , n62248 , n62249 , n62250 , n62251 , n62252 ,
     n62253 , n62254 , n62255 , n62256 , n62257 , n62258 , n62259 , n62260 , n62261 , n62262 ,
     n62263 , n62264 , n62265 , n62266 , n62267 , n62268 , n62269 , n62270 , n62271 , n62272 ,
     n62273 , n62274 , n62275 , n62276 , n62277 , n62278 , n62279 , n62280 , n62281 , n62282 ,
     n62283 , n62284 , n62285 , n62286 , n62287 , n62288 , n62289 , n62290 , n62291 , n62292 ,
     n62293 , n62294 , n62295 , n62296 , n62297 , n62298 , n62299 , n62300 , n62301 , n62302 ,
     n62303 , n62304 , n62305 , n62306 , n62307 , n62308 , n62309 , n62310 , n62311 , n62312 ,
     n62313 , n62314 , n62315 , n62316 , n62317 , n62318 , n62319 , n62320 , n62321 , n62322 ,
     n62323 , n62324 , n62325 , n62326 , n62327 , n62328 , n62329 , n62330 , n62331 , n62332 ,
     n62333 , n62334 , n62335 , n62336 , n62337 , n62338 , n62339 , n62340 , n62341 , n62342 ,
     n62343 , n62344 , n62345 , n62346 , n62347 , n62348 , n62349 , n62350 , n62351 , n62352 ,
     n62353 , n62354 , n62355 , n62356 , n62357 , n62358 , n62359 , n62360 , n62361 , n62362 ,
     n62363 , n62364 , n62365 , n62366 , n62367 , n62368 , n62369 , n62370 , n62371 , n62372 ,
     n62373 , n62374 , n62375 , n62376 , n62377 , n62378 , n62379 , n62380 , n62381 , n62382 ,
     n62383 , n62384 , n62385 , n62386 , n62387 , n62388 , n62389 , n62390 , n62391 , n62392 ,
     n62393 , n62394 , n62395 , n62396 , n62397 , n62398 , n62399 , n62400 , n62401 , n62402 ,
     n62403 , n62404 , n62405 , n62406 , n62407 , n62408 , n62409 , n62410 , n62411 , n62412 ,
     n62413 , n62414 , n62415 , n62416 , n62417 , n62418 , n62419 , n62420 , n62421 , n62422 ,
     n62423 , n62424 , n62425 , n62426 , n62427 , n62428 , n62429 , n62430 , n62431 , n62432 ,
     n62433 , n62434 , n62435 , n62436 , n62437 , n62438 , n62439 , n62440 , n62441 , n62442 ,
     n62443 , n62444 , n62445 , n62446 , n62447 , n62448 , n62449 , n62450 , n62451 , n62452 ,
     n62453 , n62454 , n62455 , n62456 , n62457 , n62458 , n62459 , n62460 , n62461 , n62462 ,
     n62463 , n62464 , n62465 , n62466 , n62467 , n62468 , n62469 , n62470 , n62471 , n62472 ,
     n62473 , n62474 , n62475 , n62476 , n62477 , n62478 , n62479 , n62480 , n62481 , n62482 ,
     n62483 , n62484 , n62485 , n62486 , n62487 , n62488 , n62489 , n62490 , n62491 , n62492 ,
     n62493 , n62494 , n62495 , n62496 , n62497 , n62498 , n62499 , n62500 , n62501 , n62502 ,
     n62503 , n62504 , n62505 , n62506 , n62507 , n62508 , n62509 , n62510 , n62511 , n62512 ,
     n62513 , n62514 , n62515 , n62516 , n62517 , n62518 , n62519 , n62520 , n62521 , n62522 ,
     n62523 , n62524 , n62525 , n62526 , n62527 , n62528 , n62529 , n62530 , n62531 , n62532 ,
     n62533 , n62534 , n62535 , n62536 , n62537 , n62538 , n62539 , n62540 , n62541 , n62542 ,
     n62543 , n62544 , n62545 , n62546 , n62547 , n62548 , n62549 , n62550 , n62551 , n62552 ,
     n62553 , n62554 , n62555 , n62556 , n62557 , n62558 , n62559 , n62560 , n62561 , n62562 ,
     n62563 , n62564 , n62565 , n62566 , n62567 , n62568 , n62569 , n62570 , n62571 , n62572 ,
     n62573 , n62574 , n62575 , n62576 , n62577 , n62578 , n62579 , n62580 , n62581 , n62582 ,
     n62583 , n62584 , n62585 , n62586 , n62587 , n62588 , n62589 , n62590 , n62591 , n62592 ,
     n62593 , n62594 , n62595 , n62596 , n62597 , n62598 , n62599 , n62600 , n62601 , n62602 ,
     n62603 , n62604 , n62605 , n62606 , n62607 , n62608 , n62609 , n62610 , n62611 , n62612 ,
     n62613 , n62614 , n62615 , n62616 , n62617 , n62618 , n62619 , n62620 , n62621 , n62622 ,
     n62623 , n62624 , n62625 , n62626 , n62627 , n62628 , n62629 , n62630 , n62631 , n62632 ,
     n62633 , n62634 , n62635 , n62636 , n62637 , n62638 , n62639 , n62640 , n62641 , n62642 ,
     n62643 , n62644 , n62645 , n62646 , n62647 , n62648 , n62649 , n62650 , n62651 , n62652 ,
     n62653 , n62654 , n62655 , n62656 , n62657 , n62658 , n62659 , n62660 , n62661 , n62662 ,
     n62663 , n62664 , n62665 , n62666 , n62667 , n62668 , n62669 , n62670 , n62671 , n62672 ,
     n62673 , n62674 , n62675 , n62676 , n62677 , n62678 , n62679 , n62680 , n62681 , n62682 ,
     n62683 , n62684 , n62685 , n62686 , n62687 , n62688 , n62689 , n62690 , n62691 , n62692 ,
     n62693 , n62694 , n62695 , n62696 , n62697 , n62698 , n62699 , n62700 , n62701 , n62702 ,
     n62703 , n62704 , n62705 , n62706 , n62707 , n62708 , n62709 , n62710 , n62711 , n62712 ,
     n62713 , n62714 , n62715 , n62716 , n62717 , n62718 , n62719 , n62720 , n62721 , n62722 ,
     n62723 , n62724 , n62725 , n62726 , n62727 , n62728 , n62729 , n62730 , n62731 , n62732 ,
     n62733 , n62734 , n62735 , n62736 , n62737 , n62738 , n62739 , n62740 , n62741 , n62742 ,
     n62743 , n62744 , n62745 , n62746 , n62747 , n62748 , n62749 , n62750 , n62751 , n62752 ,
     n62753 , n62754 , n62755 , n62756 , n62757 , n62758 , n62759 , n62760 , n62761 , n62762 ,
     n62763 , n62764 , n62765 , n62766 , n62767 , n62768 , n62769 , n62770 , n62771 , n62772 ,
     n62773 , n62774 , n62775 , n62776 , n62777 , n62778 , n62779 , n62780 , n62781 , n62782 ,
     n62783 , n62784 , n62785 , n62786 , n62787 , n62788 , n62789 , n62790 , n62791 , n62792 ,
     n62793 , n62794 , n62795 , n62796 , n62797 , n62798 , n62799 , n62800 , n62801 , n62802 ,
     n62803 , n62804 , n62805 , n62806 , n62807 , n62808 , n62809 , n62810 , n62811 , n62812 ,
     n62813 , n62814 , n62815 , n62816 , n62817 , n62818 , n62819 , n62820 , n62821 , n62822 ,
     n62823 , n62824 , n62825 , n62826 , n62827 , n62828 , n62829 , n62830 , n62831 , n62832 ,
     n62833 , n62834 , n62835 , n62836 , n62837 , n62838 , n62839 , n62840 , n62841 , n62842 ,
     n62843 , n62844 , n62845 , n62846 , n62847 , n62848 , n62849 , n62850 , n62851 , n62852 ,
     n62853 , n62854 , n62855 , n62856 , n62857 , n62858 , n62859 , n62860 , n62861 , n62862 ,
     n62863 , n62864 , n62865 , n62866 , n62867 , n62868 , n62869 , n62870 , n62871 , n62872 ,
     n62873 , n62874 , n62875 , n62876 , n62877 , n62878 , n62879 , n62880 , n62881 , n62882 ,
     n62883 , n62884 , n62885 , n62886 , n62887 , n62888 , n62889 , n62890 , n62891 , n62892 ,
     n62893 , n62894 , n62895 , n62896 , n62897 , n62898 , n62899 , n62900 , n62901 , n62902 ,
     n62903 , n62904 , n62905 , n62906 , n62907 , n62908 , n62909 , n62910 , n62911 , n62912 ,
     n62913 , n62914 , n62915 , n62916 , n62917 , n62918 , n62919 , n62920 , n62921 , n62922 ,
     n62923 , n62924 , n62925 , n62926 , n62927 , n62928 , n62929 , n62930 , n62931 , n62932 ,
     n62933 , n62934 , n62935 , n62936 , n62937 , n62938 , n62939 , n62940 , n62941 , n62942 ,
     n62943 , n62944 , n62945 , n62946 , n62947 , n62948 , n62949 , n62950 , n62951 , n62952 ,
     n62953 , n62954 , n62955 , n62956 , n62957 , n62958 , n62959 , n62960 , n62961 , n62962 ,
     n62963 , n62964 , n62965 , n62966 , n62967 , n62968 , n62969 , n62970 , n62971 , n62972 ,
     n62973 , n62974 , n62975 , n62976 , n62977 , n62978 , n62979 , n62980 , n62981 , n62982 ,
     n62983 , n62984 , n62985 , n62986 , n62987 , n62988 , n62989 , n62990 , n62991 , n62992 ,
     n62993 , n62994 , n62995 , n62996 , n62997 , n62998 , n62999 , n63000 , n63001 , n63002 ,
     n63003 , n63004 , n63005 , n63006 , n63007 , n63008 , n63009 , n63010 , n63011 , n63012 ,
     n63013 , n63014 , n63015 , n63016 , n63017 , n63018 , n63019 , n63020 , n63021 , n63022 ,
     n63023 , n63024 , n63025 , n63026 , n63027 , n63028 , n63029 , n63030 , n63031 , n63032 ,
     n63033 , n63034 , n63035 , n63036 , n63037 , n63038 , n63039 , n63040 , n63041 , n63042 ,
     n63043 , n63044 , n63045 , n63046 , n63047 , n63048 , n63049 , n63050 , n63051 , n63052 ,
     n63053 , n63054 , n63055 , n63056 , n63057 , n63058 , n63059 , n63060 , n63061 , n63062 ,
     n63063 , n63064 , n63065 , n63066 , n63067 , n63068 , n63069 , n63070 , n63071 , n63072 ,
     n63073 , n63074 , n63075 , n63076 , n63077 , n63078 , n63079 , n63080 , n63081 , n63082 ,
     n63083 , n63084 , n63085 , n63086 , n63087 , n63088 , n63089 , n63090 , n63091 , n63092 ,
     n63093 , n63094 , n63095 , n63096 , n63097 , n63098 , n63099 , n63100 , n63101 , n63102 ,
     n63103 , n63104 , n63105 , n63106 , n63107 , n63108 , n63109 , n63110 , n63111 , n63112 ,
     n63113 , n63114 , n63115 , n63116 , n63117 , n63118 , n63119 , n63120 , n63121 , n63122 ,
     n63123 , n63124 , n63125 , n63126 , n63127 , n63128 , n63129 , n63130 , n63131 , n63132 ,
     n63133 , n63134 , n63135 , n63136 , n63137 , n63138 , n63139 , n63140 , n63141 , n63142 ,
     n63143 , n63144 , n63145 , n63146 , n63147 , n63148 , n63149 , n63150 , n63151 , n63152 ,
     n63153 , n63154 , n63155 , n63156 , n63157 , n63158 , n63159 , n63160 , n63161 , n63162 ,
     n63163 , n63164 , n63165 , n63166 , n63167 , n63168 , n63169 , n63170 , n63171 , n63172 ,
     n63173 , n63174 , n63175 , n63176 , n63177 , n63178 , n63179 , n63180 , n63181 , n63182 ,
     n63183 , n63184 , n63185 , n63186 , n63187 , n63188 , n63189 , n63190 , n63191 , n63192 ,
     n63193 , n63194 , n63195 , n63196 , n63197 , n63198 , n63199 , n63200 , n63201 , n63202 ,
     n63203 , n63204 , n63205 , n63206 , n63207 , n63208 , n63209 , n63210 , n63211 , n63212 ,
     n63213 , n63214 , n63215 , n63216 , n63217 , n63218 , n63219 , n63220 , n63221 , n63222 ,
     n63223 , n63224 , n63225 , n63226 , n63227 , n63228 , n63229 , n63230 , n63231 , n63232 ,
     n63233 , n63234 , n63235 , n63236 , n63237 , n63238 , n63239 , n63240 , n63241 , n63242 ,
     n63243 , n63244 , n63245 , n63246 , n63247 , n63248 , n63249 , n63250 , n63251 , n63252 ,
     n63253 , n63254 , n63255 , n63256 , n63257 , n63258 , n63259 , n63260 , n63261 , n63262 ,
     n63263 , n63264 , n63265 , n63266 , n63267 , n63268 , n63269 , n63270 , n63271 , n63272 ,
     n63273 , n63274 , n63275 , n63276 , n63277 , n63278 , n63279 , n63280 , n63281 , n63282 ,
     n63283 , n63284 , n63285 , n63286 , n63287 , n63288 , n63289 , n63290 , n63291 , n63292 ,
     n63293 , n63294 , n63295 , n63296 , n63297 , n63298 , n63299 , n63300 , n63301 , n63302 ,
     n63303 , n63304 , n63305 , n63306 , n63307 , n63308 , n63309 , n63310 , n63311 , n63312 ,
     n63313 , n63314 , n63315 , n63316 , n63317 , n63318 , n63319 , n63320 , n63321 , n63322 ,
     n63323 , n63324 , n63325 , n63326 , n63327 , n63328 , n63329 , n63330 , n63331 , n63332 ,
     n63333 , n63334 , n63335 , n63336 , n63337 , n63338 , n63339 , n63340 , n63341 , n63342 ,
     n63343 , n63344 , n63345 , n63346 , n63347 , n63348 , n63349 , n63350 , n63351 , n63352 ,
     n63353 , n63354 , n63355 , n63356 , n63357 , n63358 , n63359 , n63360 , n63361 , n63362 ,
     n63363 , n63364 , n63365 , n63366 , n63367 , n63368 , n63369 , n63370 , n63371 , n63372 ,
     n63373 , n63374 , n63375 , n63376 , n63377 , n63378 , n63379 , n63380 , n63381 , n63382 ,
     n63383 , n63384 , n63385 , n63386 , n63387 , n63388 , n63389 , n63390 , n63391 , n63392 ,
     n63393 , n63394 , n63395 , n63396 , n63397 , n63398 , n63399 , n63400 , n63401 , n63402 ,
     n63403 , n63404 , n63405 , n63406 , n63407 , n63408 , n63409 , n63410 , n63411 , n63412 ,
     n63413 , n63414 , n63415 , n63416 , n63417 , n63418 , n63419 , n63420 , n63421 , n63422 ,
     n63423 , n63424 , n63425 , n63426 , n63427 , n63428 , n63429 , n63430 , n63431 , n63432 ,
     n63433 , n63434 , n63435 , n63436 , n63437 , n63438 , n63439 , n63440 , n63441 , n63442 ,
     n63443 , n63444 , n63445 , n63446 , n63447 , n63448 , n63449 , n63450 , n63451 , n63452 ,
     n63453 , n63454 , n63455 , n63456 , n63457 , n63458 , n63459 , n63460 , n63461 , n63462 ,
     n63463 , n63464 , n63465 , n63466 , n63467 , n63468 , n63469 , n63470 , n63471 , n63472 ,
     n63473 , n63474 , n63475 , n63476 , n63477 , n63478 , n63479 , n63480 , n63481 , n63482 ,
     n63483 , n63484 , n63485 , n63486 , n63487 , n63488 , n63489 , n63490 , n63491 , n63492 ,
     n63493 , n63494 , n63495 , n63496 , n63497 , n63498 , n63499 , n63500 , n63501 , n63502 ,
     n63503 , n63504 , n63505 , n63506 , n63507 , n63508 , n63509 , n63510 , n63511 , n63512 ,
     n63513 , n63514 , n63515 , n63516 , n63517 , n63518 , n63519 , n63520 , n63521 , n63522 ,
     n63523 , n63524 , n63525 , n63526 , n63527 , n63528 , n63529 , n63530 , n63531 , n63532 ,
     n63533 , n63534 , n63535 , n63536 , n63537 , n63538 , n63539 , n63540 , n63541 , n63542 ,
     n63543 , n63544 , n63545 , n63546 , n63547 , n63548 , n63549 , n63550 , n63551 , n63552 ,
     n63553 , n63554 , n63555 , n63556 , n63557 , n63558 , n63559 , n63560 , n63561 , n63562 ,
     n63563 , n63564 , n63565 , n63566 , n63567 , n63568 , n63569 , n63570 , n63571 , n63572 ,
     n63573 , n63574 , n63575 , n63576 , n63577 , n63578 , n63579 , n63580 , n63581 , n63582 ,
     n63583 , n63584 , n63585 , n63586 , n63587 , n63588 , n63589 , n63590 , n63591 , n63592 ,
     n63593 , n63594 , n63595 , n63596 , n63597 , n63598 , n63599 , n63600 , n63601 , n63602 ,
     n63603 , n63604 , n63605 , n63606 , n63607 , n63608 , n63609 , n63610 , n63611 , n63612 ,
     n63613 , n63614 , n63615 , n63616 , n63617 , n63618 , n63619 , n63620 , n63621 , n63622 ,
     n63623 , n63624 , n63625 , n63626 , n63627 , n63628 , n63629 , n63630 , n63631 , n63632 ,
     n63633 , n63634 , n63635 , n63636 , n63637 , n63638 , n63639 , n63640 , n63641 , n63642 ,
     n63643 , n63644 , n63645 , n63646 , n63647 , n63648 , n63649 , n63650 , n63651 , n63652 ,
     n63653 , n63654 , n63655 , n63656 , n63657 , n63658 , n63659 , n63660 , n63661 , n63662 ,
     n63663 , n63664 , n63665 , n63666 , n63667 , n63668 , n63669 , n63670 , n63671 , n63672 ,
     n63673 , n63674 , n63675 , n63676 , n63677 , n63678 , n63679 , n63680 , n63681 , n63682 ,
     n63683 , n63684 , n63685 , n63686 , n63687 , n63688 , n63689 , n63690 , n63691 , n63692 ,
     n63693 , n63694 , n63695 , n63696 , n63697 , n63698 , n63699 , n63700 , n63701 , n63702 ,
     n63703 , n63704 , n63705 , n63706 , n63707 , n63708 , n63709 , n63710 , n63711 , n63712 ,
     n63713 , n63714 , n63715 , n63716 , n63717 , n63718 , n63719 , n63720 , n63721 , n63722 ,
     n63723 , n63724 , n63725 , n63726 , n63727 , n63728 , n63729 , n63730 , n63731 , n63732 ,
     n63733 , n63734 , n63735 , n63736 , n63737 , n63738 , n63739 , n63740 , n63741 , n63742 ,
     n63743 , n63744 , n63745 , n63746 , n63747 , n63748 , n63749 , n63750 , n63751 , n63752 ,
     n63753 , n63754 , n63755 , n63756 , n63757 , n63758 , n63759 , n63760 , n63761 , n63762 ,
     n63763 , n63764 , n63765 , n63766 , n63767 , n63768 , n63769 , n63770 , n63771 , n63772 ,
     n63773 , n63774 , n63775 , n63776 , n63777 , n63778 , n63779 , n63780 , n63781 , n63782 ,
     n63783 , n63784 , n63785 , n63786 , n63787 , n63788 , n63789 , n63790 , n63791 , n63792 ,
     n63793 , n63794 , n63795 , n63796 , n63797 , n63798 , n63799 , n63800 , n63801 , n63802 ,
     n63803 , n63804 , n63805 , n63806 , n63807 , n63808 , n63809 , n63810 , n63811 , n63812 ,
     n63813 , n63814 , n63815 , n63816 , n63817 , n63818 , n63819 , n63820 , n63821 , n63822 ,
     n63823 , n63824 , n63825 , n63826 , n63827 , n63828 , n63829 , n63830 , n63831 , n63832 ,
     n63833 , n63834 , n63835 , n63836 , n63837 , n63838 , n63839 , n63840 , n63841 , n63842 ,
     n63843 , n63844 , n63845 , n63846 , n63847 , n63848 , n63849 , n63850 , n63851 , n63852 ,
     n63853 , n63854 , n63855 , n63856 , n63857 , n63858 , n63859 , n63860 , n63861 , n63862 ,
     n63863 , n63864 , n63865 , n63866 , n63867 , n63868 , n63869 , n63870 , n63871 , n63872 ,
     n63873 , n63874 , n63875 , n63876 , n63877 , n63878 , n63879 , n63880 , n63881 , n63882 ,
     n63883 , n63884 , n63885 , n63886 , n63887 , n63888 , n63889 , n63890 , n63891 , n63892 ,
     n63893 , n63894 , n63895 , n63896 , n63897 , n63898 , n63899 , n63900 , n63901 , n63902 ,
     n63903 , n63904 , n63905 , n63906 , n63907 , n63908 , n63909 , n63910 , n63911 , n63912 ,
     n63913 , n63914 , n63915 , n63916 , n63917 , n63918 , n63919 , n63920 , n63921 , n63922 ,
     n63923 , n63924 , n63925 , n63926 , n63927 , n63928 , n63929 , n63930 , n63931 , n63932 ,
     n63933 , n63934 , n63935 , n63936 , n63937 , n63938 , n63939 , n63940 , n63941 , n63942 ,
     n63943 , n63944 , n63945 , n63946 , n63947 , n63948 , n63949 , n63950 , n63951 , n63952 ,
     n63953 , n63954 , n63955 , n63956 , n63957 , n63958 , n63959 , n63960 , n63961 , n63962 ,
     n63963 , n63964 , n63965 , n63966 , n63967 , n63968 , n63969 , n63970 , n63971 , n63972 ,
     n63973 , n63974 , n63975 , n63976 , n63977 , n63978 , n63979 , n63980 , n63981 , n63982 ,
     n63983 , n63984 , n63985 , n63986 , n63987 , n63988 , n63989 , n63990 , n63991 , n63992 ,
     n63993 , n63994 , n63995 , n63996 , n63997 , n63998 , n63999 , n64000 , n64001 , n64002 ,
     n64003 , n64004 , n64005 , n64006 , n64007 , n64008 , n64009 , n64010 , n64011 , n64012 ,
     n64013 , n64014 , n64015 , n64016 , n64017 , n64018 , n64019 , n64020 , n64021 , n64022 ,
     n64023 , n64024 , n64025 , n64026 , n64027 , n64028 , n64029 , n64030 , n64031 , n64032 ,
     n64033 , n64034 , n64035 , n64036 , n64037 , n64038 , n64039 , n64040 , n64041 , n64042 ,
     n64043 , n64044 , n64045 , n64046 , n64047 , n64048 , n64049 , n64050 , n64051 , n64052 ,
     n64053 , n64054 , n64055 , n64056 , n64057 , n64058 , n64059 , n64060 , n64061 , n64062 ,
     n64063 , n64064 , n64065 , n64066 , n64067 , n64068 , n64069 , n64070 , n64071 , n64072 ,
     n64073 , n64074 , n64075 , n64076 , n64077 , n64078 , n64079 , n64080 , n64081 , n64082 ,
     n64083 , n64084 , n64085 , n64086 , n64087 , n64088 , n64089 , n64090 , n64091 , n64092 ,
     n64093 , n64094 , n64095 , n64096 , n64097 , n64098 , n64099 , n64100 , n64101 , n64102 ,
     n64103 , n64104 , n64105 , n64106 , n64107 , n64108 , n64109 , n64110 , n64111 , n64112 ,
     n64113 , n64114 , n64115 , n64116 , n64117 , n64118 , n64119 , n64120 , n64121 , n64122 ,
     n64123 , n64124 , n64125 , n64126 , n64127 , n64128 , n64129 , n64130 , n64131 , n64132 ,
     n64133 , n64134 , n64135 , n64136 , n64137 , n64138 , n64139 , n64140 , n64141 , n64142 ,
     n64143 , n64144 , n64145 , n64146 , n64147 , n64148 , n64149 , n64150 , n64151 , n64152 ,
     n64153 , n64154 , n64155 , n64156 , n64157 , n64158 , n64159 , n64160 , n64161 , n64162 ,
     n64163 , n64164 , n64165 , n64166 , n64167 , n64168 , n64169 , n64170 , n64171 , n64172 ,
     n64173 , n64174 , n64175 , n64176 , n64177 , n64178 , n64179 , n64180 , n64181 , n64182 ,
     n64183 , n64184 , n64185 , n64186 , n64187 , n64188 , n64189 , n64190 , n64191 , n64192 ,
     n64193 , n64194 , n64195 , n64196 , n64197 , n64198 , n64199 , n64200 , n64201 , n64202 ,
     n64203 , n64204 , n64205 , n64206 , n64207 , n64208 , n64209 , n64210 , n64211 , n64212 ,
     n64213 , n64214 , n64215 , n64216 , n64217 , n64218 , n64219 , n64220 , n64221 , n64222 ,
     n64223 , n64224 , n64225 , n64226 , n64227 , n64228 , n64229 , n64230 , n64231 , n64232 ,
     n64233 , n64234 , n64235 , n64236 , n64237 , n64238 , n64239 , n64240 , n64241 , n64242 ,
     n64243 , n64244 , n64245 , n64246 , n64247 , n64248 , n64249 , n64250 , n64251 , n64252 ,
     n64253 , n64254 , n64255 , n64256 , n64257 , n64258 , n64259 , n64260 , n64261 , n64262 ,
     n64263 , n64264 , n64265 , n64266 , n64267 , n64268 , n64269 , n64270 , n64271 , n64272 ,
     n64273 , n64274 , n64275 , n64276 , n64277 , n64278 , n64279 , n64280 , n64281 , n64282 ,
     n64283 , n64284 , n64285 , n64286 , n64287 , n64288 , n64289 , n64290 , n64291 , n64292 ,
     n64293 , n64294 , n64295 , n64296 , n64297 , n64298 , n64299 , n64300 , n64301 , n64302 ,
     n64303 , n64304 , n64305 , n64306 , n64307 , n64308 , n64309 , n64310 , n64311 , n64312 ,
     n64313 , n64314 , n64315 , n64316 , n64317 , n64318 , n64319 , n64320 , n64321 , n64322 ,
     n64323 , n64324 , n64325 , n64326 , n64327 , n64328 , n64329 , n64330 , n64331 , n64332 ,
     n64333 , n64334 , n64335 , n64336 , n64337 , n64338 , n64339 , n64340 , n64341 , n64342 ,
     n64343 , n64344 , n64345 , n64346 , n64347 , n64348 , n64349 , n64350 , n64351 , n64352 ,
     n64353 , n64354 , n64355 , n64356 , n64357 , n64358 , n64359 , n64360 , n64361 , n64362 ,
     n64363 , n64364 , n64365 , n64366 , n64367 , n64368 , n64369 , n64370 , n64371 , n64372 ,
     n64373 , n64374 , n64375 , n64376 , n64377 , n64378 , n64379 , n64380 , n64381 , n64382 ,
     n64383 , n64384 , n64385 , n64386 , n64387 , n64388 , n64389 , n64390 , n64391 , n64392 ,
     n64393 , n64394 , n64395 , n64396 , n64397 , n64398 , n64399 , n64400 , n64401 , n64402 ,
     n64403 , n64404 , n64405 , n64406 , n64407 , n64408 , n64409 , n64410 , n64411 , n64412 ,
     n64413 , n64414 , n64415 , n64416 , n64417 , n64418 , n64419 , n64420 , n64421 , n64422 ,
     n64423 , n64424 , n64425 , n64426 , n64427 , n64428 , n64429 , n64430 , n64431 , n64432 ,
     n64433 , n64434 , n64435 , n64436 , n64437 , n64438 , n64439 , n64440 , n64441 , n64442 ,
     n64443 , n64444 , n64445 , n64446 , n64447 , n64448 , n64449 , n64450 , n64451 , n64452 ,
     n64453 , n64454 , n64455 , n64456 , n64457 , n64458 , n64459 , n64460 , n64461 , n64462 ,
     n64463 , n64464 , n64465 , n64466 , n64467 , n64468 , n64469 , n64470 , n64471 , n64472 ,
     n64473 , n64474 , n64475 , n64476 , n64477 , n64478 , n64479 , n64480 , n64481 , n64482 ,
     n64483 , n64484 , n64485 , n64486 , n64487 , n64488 , n64489 , n64490 , n64491 , n64492 ,
     n64493 , n64494 , n64495 , n64496 , n64497 , n64498 , n64499 , n64500 , n64501 , n64502 ,
     n64503 , n64504 , n64505 , n64506 , n64507 , n64508 , n64509 , n64510 , n64511 , n64512 ,
     n64513 , n64514 , n64515 , n64516 , n64517 , n64518 , n64519 , n64520 , n64521 , n64522 ,
     n64523 , n64524 , n64525 , n64526 , n64527 , n64528 , n64529 , n64530 , n64531 , n64532 ,
     n64533 , n64534 , n64535 , n64536 , n64537 , n64538 , n64539 , n64540 , n64541 , n64542 ,
     n64543 , n64544 , n64545 , n64546 , n64547 , n64548 , n64549 , n64550 , n64551 , n64552 ,
     n64553 , n64554 , n64555 , n64556 , n64557 , n64558 , n64559 , n64560 , n64561 , n64562 ,
     n64563 , n64564 , n64565 , n64566 , n64567 , n64568 , n64569 , n64570 , n64571 , n64572 ,
     n64573 , n64574 , n64575 , n64576 , n64577 , n64578 , n64579 , n64580 , n64581 , n64582 ,
     n64583 , n64584 , n64585 , n64586 , n64587 , n64588 , n64589 , n64590 , n64591 , n64592 ,
     n64593 , n64594 , n64595 , n64596 , n64597 , n64598 , n64599 , n64600 , n64601 , n64602 ,
     n64603 , n64604 , n64605 , n64606 , n64607 , n64608 , n64609 , n64610 , n64611 , n64612 ,
     n64613 , n64614 , n64615 , n64616 , n64617 , n64618 , n64619 , n64620 , n64621 , n64622 ,
     n64623 , n64624 , n64625 , n64626 , n64627 , n64628 , n64629 , n64630 , n64631 , n64632 ,
     n64633 , n64634 , n64635 , n64636 , n64637 , n64638 , n64639 , n64640 , n64641 , n64642 ,
     n64643 , n64644 , n64645 , n64646 , n64647 , n64648 , n64649 , n64650 , n64651 , n64652 ,
     n64653 , n64654 , n64655 , n64656 , n64657 , n64658 , n64659 , n64660 , n64661 , n64662 ,
     n64663 , n64664 , n64665 , n64666 , n64667 , n64668 , n64669 , n64670 , n64671 , n64672 ,
     n64673 , n64674 , n64675 , n64676 , n64677 , n64678 , n64679 , n64680 , n64681 , n64682 ,
     n64683 , n64684 , n64685 , n64686 , n64687 , n64688 , n64689 , n64690 , n64691 , n64692 ,
     n64693 , n64694 , n64695 , n64696 , n64697 , n64698 , n64699 , n64700 , n64701 , n64702 ,
     n64703 , n64704 , n64705 , n64706 , n64707 , n64708 , n64709 , n64710 , n64711 , n64712 ,
     n64713 , n64714 , n64715 , n64716 , n64717 , n64718 , n64719 , n64720 , n64721 , n64722 ,
     n64723 , n64724 , n64725 , n64726 , n64727 , n64728 , n64729 , n64730 , n64731 , n64732 ,
     n64733 , n64734 , n64735 , n64736 , n64737 , n64738 , n64739 , n64740 , n64741 , n64742 ,
     n64743 , n64744 , n64745 , n64746 , n64747 , n64748 , n64749 , n64750 , n64751 , n64752 ,
     n64753 , n64754 , n64755 , n64756 , n64757 , n64758 , n64759 , n64760 , n64761 , n64762 ,
     n64763 , n64764 , n64765 , n64766 , n64767 , n64768 , n64769 , n64770 , n64771 , n64772 ,
     n64773 , n64774 , n64775 , n64776 , n64777 , n64778 , n64779 , n64780 , n64781 , n64782 ,
     n64783 , n64784 , n64785 , n64786 , n64787 , n64788 , n64789 , n64790 , n64791 , n64792 ,
     n64793 , n64794 , n64795 , n64796 , n64797 , n64798 , n64799 , n64800 , n64801 , n64802 ,
     n64803 , n64804 , n64805 , n64806 , n64807 , n64808 , n64809 , n64810 , n64811 , n64812 ,
     n64813 , n64814 , n64815 , n64816 , n64817 , n64818 , n64819 , n64820 , n64821 , n64822 ,
     n64823 , n64824 , n64825 , n64826 , n64827 , n64828 , n64829 , n64830 , n64831 , n64832 ,
     n64833 , n64834 , n64835 , n64836 , n64837 , n64838 , n64839 , n64840 , n64841 , n64842 ,
     n64843 , n64844 , n64845 , n64846 , n64847 , n64848 , n64849 , n64850 , n64851 , n64852 ,
     n64853 , n64854 , n64855 , n64856 , n64857 , n64858 , n64859 , n64860 , n64861 , n64862 ,
     n64863 , n64864 , n64865 , n64866 , n64867 , n64868 , n64869 , n64870 , n64871 , n64872 ,
     n64873 , n64874 , n64875 , n64876 , n64877 , n64878 , n64879 , n64880 , n64881 , n64882 ,
     n64883 , n64884 , n64885 , n64886 , n64887 , n64888 , n64889 , n64890 , n64891 , n64892 ,
     n64893 , n64894 , n64895 , n64896 , n64897 , n64898 , n64899 , n64900 , n64901 , n64902 ,
     n64903 , n64904 , n64905 , n64906 , n64907 , n64908 , n64909 , n64910 , n64911 , n64912 ,
     n64913 , n64914 , n64915 , n64916 , n64917 , n64918 , n64919 , n64920 , n64921 , n64922 ,
     n64923 , n64924 , n64925 , n64926 , n64927 , n64928 , n64929 , n64930 , n64931 , n64932 ,
     n64933 , n64934 , n64935 , n64936 , n64937 , n64938 , n64939 , n64940 , n64941 , n64942 ,
     n64943 , n64944 , n64945 , n64946 , n64947 , n64948 , n64949 , n64950 , n64951 , n64952 ,
     n64953 , n64954 , n64955 , n64956 , n64957 , n64958 , n64959 , n64960 , n64961 , n64962 ,
     n64963 , n64964 , n64965 , n64966 , n64967 , n64968 , n64969 , n64970 , n64971 , n64972 ,
     n64973 , n64974 , n64975 , n64976 , n64977 , n64978 , n64979 , n64980 , n64981 , n64982 ,
     n64983 , n64984 , n64985 , n64986 , n64987 , n64988 , n64989 , n64990 , n64991 , n64992 ,
     n64993 , n64994 , n64995 , n64996 , n64997 , n64998 , n64999 , n65000 , n65001 , n65002 ,
     n65003 , n65004 , n65005 , n65006 , n65007 , n65008 , n65009 , n65010 , n65011 , n65012 ,
     n65013 , n65014 , n65015 , n65016 , n65017 , n65018 , n65019 , n65020 , n65021 , n65022 ,
     n65023 , n65024 , n65025 , n65026 , n65027 , n65028 , n65029 , n65030 , n65031 , n65032 ,
     n65033 , n65034 , n65035 , n65036 , n65037 , n65038 , n65039 , n65040 , n65041 , n65042 ,
     n65043 , n65044 , n65045 , n65046 , n65047 , n65048 , n65049 , n65050 , n65051 , n65052 ,
     n65053 , n65054 , n65055 , n65056 , n65057 , n65058 , n65059 , n65060 , n65061 , n65062 ,
     n65063 , n65064 , n65065 , n65066 , n65067 , n65068 , n65069 , n65070 , n65071 , n65072 ,
     n65073 , n65074 , n65075 , n65076 , n65077 , n65078 , n65079 , n65080 , n65081 , n65082 ,
     n65083 , n65084 , n65085 , n65086 , n65087 , n65088 , n65089 , n65090 , n65091 , n65092 ,
     n65093 , n65094 , n65095 , n65096 , n65097 , n65098 , n65099 , n65100 , n65101 , n65102 ,
     n65103 , n65104 , n65105 , n65106 , n65107 , n65108 , n65109 , n65110 , n65111 , n65112 ,
     n65113 , n65114 , n65115 , n65116 , n65117 , n65118 , n65119 , n65120 , n65121 , n65122 ,
     n65123 , n65124 , n65125 , n65126 , n65127 , n65128 , n65129 , n65130 , n65131 , n65132 ,
     n65133 , n65134 , n65135 , n65136 , n65137 , n65138 , n65139 , n65140 , n65141 , n65142 ,
     n65143 , n65144 , n65145 , n65146 , n65147 , n65148 , n65149 , n65150 , n65151 , n65152 ,
     n65153 , n65154 , n65155 , n65156 , n65157 , n65158 , n65159 , n65160 , n65161 , n65162 ,
     n65163 , n65164 , n65165 , n65166 , n65167 , n65168 , n65169 , n65170 , n65171 , n65172 ,
     n65173 , n65174 , n65175 , n65176 , n65177 , n65178 , n65179 , n65180 , n65181 , n65182 ,
     n65183 , n65184 , n65185 , n65186 , n65187 , n65188 , n65189 , n65190 , n65191 , n65192 ,
     n65193 , n65194 , n65195 , n65196 , n65197 , n65198 , n65199 , n65200 , n65201 , n65202 ,
     n65203 , n65204 , n65205 , n65206 , n65207 , n65208 , n65209 , n65210 , n65211 , n65212 ,
     n65213 , n65214 , n65215 , n65216 , n65217 , n65218 , n65219 , n65220 , n65221 , n65222 ,
     n65223 , n65224 , n65225 , n65226 , n65227 , n65228 , n65229 , n65230 , n65231 , n65232 ,
     n65233 , n65234 , n65235 , n65236 , n65237 , n65238 , n65239 , n65240 , n65241 , n65242 ,
     n65243 , n65244 , n65245 , n65246 , n65247 , n65248 , n65249 , n65250 , n65251 , n65252 ,
     n65253 , n65254 , n65255 , n65256 , n65257 , n65258 , n65259 , n65260 , n65261 , n65262 ,
     n65263 , n65264 , n65265 , n65266 , n65267 , n65268 , n65269 , n65270 , n65271 , n65272 ,
     n65273 , n65274 , n65275 , n65276 , n65277 , n65278 , n65279 , n65280 , n65281 , n65282 ,
     n65283 , n65284 , n65285 , n65286 , n65287 , n65288 , n65289 , n65290 , n65291 , n65292 ,
     n65293 , n65294 , n65295 , n65296 , n65297 , n65298 , n65299 , n65300 , n65301 , n65302 ,
     n65303 , n65304 , n65305 , n65306 , n65307 , n65308 , n65309 , n65310 , n65311 , n65312 ,
     n65313 , n65314 , n65315 , n65316 , n65317 , n65318 , n65319 , n65320 , n65321 , n65322 ,
     n65323 , n65324 , n65325 , n65326 , n65327 , n65328 , n65329 , n65330 , n65331 , n65332 ,
     n65333 , n65334 , n65335 , n65336 , n65337 , n65338 , n65339 , n65340 , n65341 , n65342 ,
     n65343 , n65344 , n65345 , n65346 , n65347 , n65348 , n65349 , n65350 , n65351 , n65352 ,
     n65353 , n65354 , n65355 , n65356 , n65357 , n65358 , n65359 , n65360 , n65361 , n65362 ,
     n65363 , n65364 , n65365 , n65366 , n65367 , n65368 , n65369 , n65370 , n65371 , n65372 ,
     n65373 , n65374 , n65375 , n65376 , n65377 , n65378 , n65379 , n65380 , n65381 , n65382 ,
     n65383 , n65384 , n65385 , n65386 , n65387 , n65388 , n65389 , n65390 , n65391 , n65392 ,
     n65393 , n65394 , n65395 , n65396 , n65397 , n65398 , n65399 , n65400 , n65401 , n65402 ,
     n65403 , n65404 , n65405 , n65406 , n65407 , n65408 , n65409 , n65410 , n65411 , n65412 ,
     n65413 , n65414 , n65415 , n65416 , n65417 , n65418 , n65419 , n65420 , n65421 , n65422 ,
     n65423 , n65424 , n65425 , n65426 , n65427 , n65428 , n65429 , n65430 , n65431 , n65432 ,
     n65433 , n65434 , n65435 , n65436 , n65437 , n65438 , n65439 , n65440 , n65441 , n65442 ,
     n65443 , n65444 , n65445 , n65446 , n65447 , n65448 , n65449 , n65450 , n65451 , n65452 ,
     n65453 , n65454 , n65455 , n65456 , n65457 , n65458 , n65459 , n65460 , n65461 , n65462 ,
     n65463 , n65464 , n65465 , n65466 , n65467 , n65468 , n65469 , n65470 , n65471 , n65472 ,
     n65473 , n65474 , n65475 , n65476 , n65477 , n65478 , n65479 , n65480 , n65481 , n65482 ,
     n65483 , n65484 , n65485 , n65486 , n65487 , n65488 , n65489 , n65490 , n65491 , n65492 ,
     n65493 , n65494 , n65495 , n65496 , n65497 , n65498 , n65499 , n65500 , n65501 , n65502 ,
     n65503 , n65504 , n65505 , n65506 , n65507 , n65508 , n65509 , n65510 , n65511 , n65512 ,
     n65513 , n65514 , n65515 , n65516 , n65517 , n65518 , n65519 , n65520 , n65521 , n65522 ,
     n65523 , n65524 , n65525 , n65526 , n65527 , n65528 , n65529 , n65530 , n65531 , n65532 ,
     n65533 , n65534 , n65535 , n65536 , n65537 , n65538 , n65539 , n65540 , n65541 , n65542 ,
     n65543 , n65544 , n65545 , n65546 , n65547 , n65548 , n65549 , n65550 , n65551 , n65552 ,
     n65553 , n65554 , n65555 , n65556 , n65557 , n65558 , n65559 , n65560 , n65561 , n65562 ,
     n65563 , n65564 , n65565 , n65566 , n65567 , n65568 , n65569 , n65570 , n65571 , n65572 ,
     n65573 , n65574 , n65575 , n65576 , n65577 , n65578 , n65579 , n65580 , n65581 , n65582 ,
     n65583 , n65584 , n65585 , n65586 , n65587 , n65588 , n65589 , n65590 , n65591 , n65592 ,
     n65593 , n65594 , n65595 , n65596 , n65597 , n65598 , n65599 , n65600 , n65601 , n65602 ,
     n65603 , n65604 , n65605 , n65606 , n65607 , n65608 , n65609 , n65610 , n65611 , n65612 ,
     n65613 , n65614 , n65615 , n65616 , n65617 , n65618 , n65619 , n65620 , n65621 , n65622 ,
     n65623 , n65624 , n65625 , n65626 , n65627 , n65628 , n65629 , n65630 , n65631 , n65632 ,
     n65633 , n65634 , n65635 , n65636 , n65637 , n65638 , n65639 , n65640 , n65641 , n65642 ,
     n65643 , n65644 , n65645 , n65646 , n65647 , n65648 , n65649 , n65650 , n65651 , n65652 ,
     n65653 , n65654 , n65655 , n65656 , n65657 , n65658 , n65659 , n65660 , n65661 , n65662 ,
     n65663 , n65664 , n65665 , n65666 , n65667 , n65668 , n65669 , n65670 , n65671 , n65672 ,
     n65673 , n65674 , n65675 , n65676 , n65677 , n65678 , n65679 , n65680 , n65681 , n65682 ,
     n65683 , n65684 , n65685 , n65686 , n65687 , n65688 , n65689 , n65690 , n65691 , n65692 ,
     n65693 , n65694 , n65695 , n65696 , n65697 , n65698 , n65699 , n65700 , n65701 , n65702 ,
     n65703 , n65704 , n65705 , n65706 , n65707 , n65708 , n65709 , n65710 , n65711 , n65712 ,
     n65713 , n65714 , n65715 , n65716 , n65717 , n65718 , n65719 , n65720 , n65721 , n65722 ,
     n65723 , n65724 , n65725 , n65726 , n65727 , n65728 , n65729 , n65730 , n65731 , n65732 ,
     n65733 , n65734 , n65735 , n65736 , n65737 , n65738 , n65739 , n65740 , n65741 , n65742 ,
     n65743 , n65744 , n65745 , n65746 , n65747 , n65748 , n65749 , n65750 , n65751 , n65752 ,
     n65753 , n65754 , n65755 , n65756 , n65757 , n65758 , n65759 , n65760 , n65761 , n65762 ,
     n65763 , n65764 , n65765 , n65766 , n65767 , n65768 , n65769 , n65770 , n65771 , n65772 ,
     n65773 , n65774 , n65775 , n65776 , n65777 , n65778 , n65779 , n65780 , n65781 , n65782 ,
     n65783 , n65784 , n65785 , n65786 , n65787 , n65788 , n65789 , n65790 , n65791 , n65792 ,
     n65793 , n65794 , n65795 , n65796 , n65797 , n65798 , n65799 , n65800 , n65801 , n65802 ,
     n65803 , n65804 , n65805 , n65806 , n65807 , n65808 , n65809 , n65810 , n65811 , n65812 ,
     n65813 , n65814 , n65815 , n65816 , n65817 , n65818 , n65819 , n65820 , n65821 , n65822 ,
     n65823 , n65824 , n65825 , n65826 , n65827 , n65828 , n65829 , n65830 , n65831 , n65832 ,
     n65833 , n65834 , n65835 , n65836 , n65837 , n65838 , n65839 , n65840 , n65841 , n65842 ,
     n65843 , n65844 , n65845 , n65846 , n65847 , n65848 , n65849 , n65850 , n65851 , n65852 ,
     n65853 , n65854 , n65855 , n65856 , n65857 , n65858 , n65859 , n65860 , n65861 , n65862 ,
     n65863 , n65864 , n65865 , n65866 , n65867 , n65868 , n65869 , n65870 , n65871 , n65872 ,
     n65873 , n65874 , n65875 , n65876 , n65877 , n65878 , n65879 , n65880 , n65881 , n65882 ,
     n65883 , n65884 , n65885 , n65886 , n65887 , n65888 , n65889 , n65890 , n65891 , n65892 ,
     n65893 , n65894 , n65895 , n65896 , n65897 , n65898 , n65899 , n65900 , n65901 , n65902 ,
     n65903 , n65904 , n65905 , n65906 , n65907 , n65908 , n65909 , n65910 , n65911 , n65912 ,
     n65913 , n65914 , n65915 , n65916 , n65917 , n65918 , n65919 , n65920 , n65921 , n65922 ,
     n65923 , n65924 , n65925 , n65926 , n65927 , n65928 , n65929 , n65930 , n65931 , n65932 ,
     n65933 , n65934 , n65935 , n65936 , n65937 , n65938 , n65939 , n65940 , n65941 , n65942 ,
     n65943 , n65944 , n65945 , n65946 , n65947 , n65948 , n65949 , n65950 , n65951 , n65952 ,
     n65953 , n65954 , n65955 , n65956 , n65957 , n65958 , n65959 , n65960 , n65961 , n65962 ,
     n65963 , n65964 , n65965 , n65966 , n65967 , n65968 , n65969 , n65970 , n65971 , n65972 ,
     n65973 , n65974 , n65975 , n65976 , n65977 , n65978 , n65979 , n65980 , n65981 , n65982 ,
     n65983 , n65984 , n65985 , n65986 , n65987 , n65988 , n65989 , n65990 , n65991 , n65992 ,
     n65993 , n65994 , n65995 , n65996 , n65997 , n65998 , n65999 , n66000 , n66001 , n66002 ,
     n66003 , n66004 , n66005 , n66006 , n66007 , n66008 , n66009 , n66010 , n66011 , n66012 ,
     n66013 , n66014 , n66015 , n66016 , n66017 , n66018 , n66019 , n66020 , n66021 , n66022 ,
     n66023 , n66024 , n66025 , n66026 , n66027 , n66028 , n66029 , n66030 , n66031 , n66032 ,
     n66033 , n66034 , n66035 , n66036 , n66037 , n66038 , n66039 , n66040 , n66041 , n66042 ,
     n66043 , n66044 , n66045 , n66046 , n66047 , n66048 , n66049 , n66050 , n66051 , n66052 ,
     n66053 , n66054 , n66055 , n66056 , n66057 , n66058 , n66059 , n66060 , n66061 , n66062 ,
     n66063 , n66064 , n66065 , n66066 , n66067 , n66068 , n66069 , n66070 , n66071 , n66072 ,
     n66073 , n66074 , n66075 , n66076 , n66077 , n66078 , n66079 , n66080 , n66081 , n66082 ,
     n66083 , n66084 , n66085 , n66086 , n66087 , n66088 , n66089 , n66090 , n66091 , n66092 ,
     n66093 , n66094 , n66095 , n66096 , n66097 , n66098 , n66099 , n66100 , n66101 , n66102 ,
     n66103 , n66104 , n66105 , n66106 , n66107 , n66108 , n66109 , n66110 , n66111 , n66112 ,
     n66113 , n66114 , n66115 , n66116 , n66117 , n66118 , n66119 , n66120 , n66121 , n66122 ,
     n66123 , n66124 , n66125 , n66126 , n66127 , n66128 , n66129 , n66130 , n66131 , n66132 ,
     n66133 , n66134 , n66135 , n66136 , n66137 , n66138 , n66139 , n66140 , n66141 , n66142 ,
     n66143 , n66144 , n66145 , n66146 , n66147 , n66148 , n66149 , n66150 , n66151 , n66152 ,
     n66153 , n66154 , n66155 , n66156 , n66157 , n66158 , n66159 , n66160 , n66161 , n66162 ,
     n66163 , n66164 , n66165 , n66166 , n66167 , n66168 , n66169 , n66170 , n66171 , n66172 ,
     n66173 , n66174 , n66175 , n66176 , n66177 , n66178 , n66179 , n66180 , n66181 , n66182 ,
     n66183 , n66184 , n66185 , n66186 , n66187 , n66188 , n66189 , n66190 , n66191 , n66192 ,
     n66193 , n66194 , n66195 , n66196 , n66197 , n66198 , n66199 , n66200 , n66201 , n66202 ,
     n66203 , n66204 , n66205 , n66206 , n66207 , n66208 , n66209 , n66210 , n66211 , n66212 ,
     n66213 , n66214 , n66215 , n66216 , n66217 , n66218 , n66219 , n66220 , n66221 , n66222 ,
     n66223 , n66224 , n66225 , n66226 , n66227 , n66228 , n66229 , n66230 , n66231 , n66232 ,
     n66233 , n66234 , n66235 , n66236 , n66237 , n66238 , n66239 , n66240 , n66241 , n66242 ,
     n66243 , n66244 , n66245 , n66246 , n66247 , n66248 , n66249 , n66250 , n66251 , n66252 ,
     n66253 , n66254 , n66255 , n66256 , n66257 , n66258 , n66259 , n66260 , n66261 , n66262 ,
     n66263 , n66264 , n66265 , n66266 , n66267 , n66268 , n66269 , n66270 , n66271 , n66272 ,
     n66273 , n66274 , n66275 , n66276 , n66277 , n66278 , n66279 , n66280 , n66281 , n66282 ,
     n66283 , n66284 , n66285 , n66286 , n66287 , n66288 , n66289 , n66290 , n66291 , n66292 ,
     n66293 , n66294 , n66295 , n66296 , n66297 , n66298 , n66299 , n66300 , n66301 , n66302 ,
     n66303 , n66304 , n66305 , n66306 , n66307 , n66308 , n66309 , n66310 , n66311 , n66312 ,
     n66313 , n66314 , n66315 , n66316 , n66317 , n66318 , n66319 , n66320 , n66321 , n66322 ,
     n66323 , n66324 , n66325 , n66326 , n66327 , n66328 , n66329 , n66330 , n66331 , n66332 ,
     n66333 , n66334 , n66335 , n66336 , n66337 , n66338 , n66339 , n66340 , n66341 , n66342 ,
     n66343 , n66344 , n66345 , n66346 , n66347 , n66348 , n66349 , n66350 , n66351 , n66352 ,
     n66353 , n66354 , n66355 , n66356 , n66357 , n66358 , n66359 , n66360 , n66361 , n66362 ,
     n66363 , n66364 , n66365 , n66366 , n66367 , n66368 , n66369 , n66370 , n66371 , n66372 ,
     n66373 , n66374 , n66375 , n66376 , n66377 , n66378 , n66379 , n66380 , n66381 , n66382 ,
     n66383 , n66384 , n66385 , n66386 , n66387 , n66388 , n66389 , n66390 , n66391 , n66392 ,
     n66393 , n66394 , n66395 , n66396 , n66397 , n66398 , n66399 , n66400 , n66401 , n66402 ,
     n66403 , n66404 , n66405 , n66406 , n66407 , n66408 , n66409 , n66410 , n66411 , n66412 ,
     n66413 , n66414 , n66415 , n66416 , n66417 , n66418 , n66419 , n66420 , n66421 , n66422 ,
     n66423 , n66424 , n66425 , n66426 , n66427 , n66428 , n66429 , n66430 , n66431 , n66432 ,
     n66433 , n66434 , n66435 , n66436 , n66437 , n66438 , n66439 , n66440 , n66441 , n66442 ,
     n66443 , n66444 , n66445 , n66446 , n66447 , n66448 , n66449 , n66450 , n66451 , n66452 ,
     n66453 , n66454 , n66455 , n66456 , n66457 , n66458 , n66459 , n66460 , n66461 , n66462 ,
     n66463 , n66464 , n66465 , n66466 , n66467 , n66468 , n66469 , n66470 , n66471 , n66472 ,
     n66473 , n66474 , n66475 , n66476 , n66477 , n66478 , n66479 , n66480 , n66481 , n66482 ,
     n66483 , n66484 , n66485 , n66486 , n66487 , n66488 , n66489 , n66490 , n66491 , n66492 ,
     n66493 , n66494 , n66495 , n66496 , n66497 , n66498 , n66499 , n66500 , n66501 , n66502 ,
     n66503 , n66504 , n66505 , n66506 , n66507 , n66508 , n66509 , n66510 , n66511 , n66512 ,
     n66513 , n66514 , n66515 , n66516 , n66517 , n66518 , n66519 , n66520 , n66521 , n66522 ,
     n66523 , n66524 , n66525 , n66526 , n66527 , n66528 , n66529 , n66530 , n66531 , n66532 ,
     n66533 , n66534 , n66535 , n66536 , n66537 , n66538 , n66539 , n66540 , n66541 , n66542 ,
     n66543 , n66544 , n66545 , n66546 , n66547 , n66548 , n66549 , n66550 , n66551 , n66552 ,
     n66553 , n66554 , n66555 , n66556 , n66557 , n66558 , n66559 , n66560 , n66561 , n66562 ,
     n66563 , n66564 , n66565 , n66566 , n66567 , n66568 , n66569 , n66570 , n66571 , n66572 ,
     n66573 , n66574 , n66575 , n66576 , n66577 , n66578 , n66579 , n66580 , n66581 , n66582 ,
     n66583 , n66584 , n66585 , n66586 , n66587 , n66588 , n66589 , n66590 , n66591 , n66592 ,
     n66593 , n66594 , n66595 , n66596 , n66597 , n66598 , n66599 , n66600 , n66601 , n66602 ,
     n66603 , n66604 , n66605 , n66606 , n66607 , n66608 , n66609 , n66610 , n66611 , n66612 ,
     n66613 , n66614 , n66615 , n66616 , n66617 , n66618 , n66619 , n66620 , n66621 , n66622 ,
     n66623 , n66624 , n66625 , n66626 , n66627 , n66628 , n66629 , n66630 , n66631 , n66632 ,
     n66633 , n66634 , n66635 , n66636 , n66637 , n66638 , n66639 , n66640 , n66641 , n66642 ,
     n66643 , n66644 , n66645 , n66646 , n66647 , n66648 , n66649 , n66650 , n66651 , n66652 ,
     n66653 , n66654 , n66655 , n66656 , n66657 , n66658 , n66659 , n66660 , n66661 , n66662 ,
     n66663 , n66664 , n66665 , n66666 , n66667 , n66668 , n66669 , n66670 , n66671 , n66672 ,
     n66673 , n66674 , n66675 , n66676 , n66677 , n66678 , n66679 , n66680 , n66681 , n66682 ,
     n66683 , n66684 , n66685 , n66686 , n66687 , n66688 , n66689 , n66690 , n66691 , n66692 ,
     n66693 , n66694 , n66695 , n66696 , n66697 , n66698 , n66699 , n66700 , n66701 , n66702 ,
     n66703 , n66704 , n66705 , n66706 , n66707 , n66708 , n66709 , n66710 , n66711 , n66712 ,
     n66713 , n66714 , n66715 , n66716 , n66717 , n66718 , n66719 , n66720 , n66721 , n66722 ,
     n66723 , n66724 , n66725 , n66726 , n66727 , n66728 , n66729 , n66730 , n66731 , n66732 ,
     n66733 , n66734 , n66735 , n66736 , n66737 , n66738 , n66739 , n66740 , n66741 , n66742 ,
     n66743 , n66744 , n66745 , n66746 , n66747 , n66748 , n66749 , n66750 , n66751 , n66752 ,
     n66753 , n66754 , n66755 , n66756 , n66757 , n66758 , n66759 , n66760 , n66761 , n66762 ,
     n66763 , n66764 , n66765 , n66766 , n66767 , n66768 , n66769 , n66770 , n66771 , n66772 ,
     n66773 , n66774 , n66775 , n66776 , n66777 , n66778 , n66779 , n66780 , n66781 , n66782 ,
     n66783 , n66784 , n66785 , n66786 , n66787 , n66788 , n66789 , n66790 , n66791 , n66792 ,
     n66793 , n66794 , n66795 , n66796 , n66797 , n66798 , n66799 , n66800 , n66801 , n66802 ,
     n66803 , n66804 , n66805 , n66806 , n66807 , n66808 , n66809 , n66810 , n66811 , n66812 ,
     n66813 , n66814 , n66815 , n66816 , n66817 , n66818 , n66819 , n66820 , n66821 , n66822 ,
     n66823 , n66824 , n66825 , n66826 , n66827 , n66828 , n66829 , n66830 , n66831 , n66832 ,
     n66833 , n66834 , n66835 , n66836 , n66837 , n66838 , n66839 , n66840 , n66841 , n66842 ,
     n66843 , n66844 , n66845 , n66846 , n66847 , n66848 , n66849 , n66850 , n66851 , n66852 ,
     n66853 , n66854 , n66855 , n66856 , n66857 , n66858 , n66859 , n66860 , n66861 , n66862 ,
     n66863 , n66864 , n66865 , n66866 , n66867 , n66868 , n66869 , n66870 , n66871 , n66872 ,
     n66873 , n66874 , n66875 , n66876 , n66877 , n66878 , n66879 , n66880 , n66881 , n66882 ,
     n66883 , n66884 , n66885 , n66886 , n66887 , n66888 , n66889 , n66890 , n66891 , n66892 ,
     n66893 , n66894 , n66895 , n66896 , n66897 , n66898 , n66899 , n66900 , n66901 , n66902 ,
     n66903 , n66904 , n66905 , n66906 , n66907 , n66908 , n66909 , n66910 , n66911 , n66912 ,
     n66913 , n66914 , n66915 , n66916 , n66917 , n66918 , n66919 , n66920 , n66921 , n66922 ,
     n66923 , n66924 , n66925 , n66926 , n66927 , n66928 , n66929 , n66930 , n66931 , n66932 ,
     n66933 , n66934 , n66935 , n66936 , n66937 , n66938 , n66939 , n66940 , n66941 , n66942 ,
     n66943 , n66944 , n66945 , n66946 , n66947 , n66948 , n66949 , n66950 , n66951 , n66952 ,
     n66953 , n66954 , n66955 , n66956 , n66957 , n66958 , n66959 , n66960 , n66961 , n66962 ,
     n66963 , n66964 , n66965 , n66966 , n66967 , n66968 , n66969 , n66970 , n66971 , n66972 ,
     n66973 , n66974 , n66975 , n66976 , n66977 , n66978 , n66979 , n66980 , n66981 , n66982 ,
     n66983 , n66984 , n66985 , n66986 , n66987 , n66988 , n66989 , n66990 , n66991 , n66992 ,
     n66993 , n66994 , n66995 , n66996 , n66997 , n66998 , n66999 , n67000 , n67001 , n67002 ,
     n67003 , n67004 , n67005 , n67006 , n67007 , n67008 , n67009 , n67010 , n67011 , n67012 ,
     n67013 , n67014 , n67015 , n67016 , n67017 , n67018 , n67019 , n67020 , n67021 , n67022 ,
     n67023 , n67024 , n67025 , n67026 , n67027 , n67028 , n67029 , n67030 , n67031 , n67032 ,
     n67033 , n67034 , n67035 , n67036 , n67037 , n67038 , n67039 , n67040 , n67041 , n67042 ,
     n67043 , n67044 , n67045 , n67046 , n67047 , n67048 , n67049 , n67050 , n67051 , n67052 ,
     n67053 , n67054 , n67055 , n67056 , n67057 , n67058 , n67059 , n67060 , n67061 , n67062 ,
     n67063 , n67064 , n67065 , n67066 , n67067 , n67068 , n67069 , n67070 , n67071 , n67072 ,
     n67073 , n67074 , n67075 , n67076 , n67077 , n67078 , n67079 , n67080 , n67081 , n67082 ,
     n67083 , n67084 , n67085 , n67086 , n67087 , n67088 , n67089 , n67090 , n67091 , n67092 ,
     n67093 , n67094 , n67095 , n67096 , n67097 , n67098 , n67099 , n67100 , n67101 , n67102 ,
     n67103 , n67104 , n67105 , n67106 , n67107 , n67108 , n67109 , n67110 , n67111 , n67112 ,
     n67113 , n67114 , n67115 , n67116 , n67117 , n67118 , n67119 , n67120 , n67121 , n67122 ,
     n67123 , n67124 , n67125 , n67126 , n67127 , n67128 , n67129 , n67130 , n67131 , n67132 ,
     n67133 , n67134 , n67135 , n67136 , n67137 , n67138 , n67139 , n67140 , n67141 , n67142 ,
     n67143 , n67144 , n67145 , n67146 , n67147 , n67148 , n67149 , n67150 , n67151 , n67152 ,
     n67153 , n67154 , n67155 , n67156 , n67157 , n67158 , n67159 , n67160 , n67161 , n67162 ,
     n67163 , n67164 , n67165 , n67166 , n67167 , n67168 , n67169 , n67170 , n67171 , n67172 ,
     n67173 , n67174 , n67175 , n67176 , n67177 , n67178 , n67179 , n67180 , n67181 , n67182 ,
     n67183 , n67184 , n67185 , n67186 , n67187 , n67188 , n67189 , n67190 , n67191 , n67192 ,
     n67193 , n67194 , n67195 , n67196 , n67197 , n67198 , n67199 , n67200 , n67201 , n67202 ,
     n67203 , n67204 , n67205 , n67206 , n67207 , n67208 , n67209 , n67210 , n67211 , n67212 ,
     n67213 , n67214 , n67215 , n67216 , n67217 , n67218 , n67219 , n67220 , n67221 , n67222 ,
     n67223 , n67224 , n67225 , n67226 , n67227 , n67228 , n67229 , n67230 , n67231 , n67232 ,
     n67233 , n67234 , n67235 , n67236 , n67237 , n67238 , n67239 , n67240 , n67241 , n67242 ,
     n67243 , n67244 , n67245 , n67246 , n67247 , n67248 , n67249 , n67250 , n67251 , n67252 ,
     n67253 , n67254 , n67255 , n67256 , n67257 , n67258 , n67259 , n67260 , n67261 , n67262 ,
     n67263 , n67264 , n67265 , n67266 , n67267 , n67268 , n67269 , n67270 , n67271 , n67272 ,
     n67273 , n67274 , n67275 , n67276 , n67277 , n67278 , n67279 , n67280 , n67281 , n67282 ,
     n67283 , n67284 , n67285 , n67286 , n67287 , n67288 , n67289 , n67290 , n67291 , n67292 ,
     n67293 , n67294 , n67295 , n67296 , n67297 , n67298 , n67299 , n67300 , n67301 , n67302 ,
     n67303 , n67304 , n67305 , n67306 , n67307 , n67308 , n67309 , n67310 , n67311 , n67312 ,
     n67313 , n67314 , n67315 , n67316 , n67317 , n67318 , n67319 , n67320 , n67321 , n67322 ,
     n67323 , n67324 , n67325 , n67326 , n67327 , n67328 , n67329 , n67330 , n67331 , n67332 ,
     n67333 , n67334 , n67335 , n67336 , n67337 , n67338 , n67339 , n67340 , n67341 , n67342 ,
     n67343 , n67344 , n67345 , n67346 , n67347 , n67348 , n67349 , n67350 , n67351 , n67352 ,
     n67353 , n67354 , n67355 , n67356 , n67357 , n67358 , n67359 , n67360 , n67361 , n67362 ,
     n67363 , n67364 , n67365 , n67366 , n67367 , n67368 , n67369 , n67370 , n67371 , n67372 ,
     n67373 , n67374 , n67375 , n67376 , n67377 , n67378 , n67379 , n67380 , n67381 , n67382 ,
     n67383 , n67384 , n67385 , n67386 , n67387 , n67388 , n67389 , n67390 , n67391 , n67392 ,
     n67393 , n67394 , n67395 , n67396 , n67397 , n67398 , n67399 , n67400 , n67401 , n67402 ,
     n67403 , n67404 , n67405 , n67406 , n67407 , n67408 , n67409 , n67410 , n67411 , n67412 ,
     n67413 , n67414 , n67415 , n67416 , n67417 , n67418 , n67419 , n67420 , n67421 , n67422 ,
     n67423 , n67424 , n67425 , n67426 , n67427 , n67428 , n67429 , n67430 , n67431 , n67432 ,
     n67433 , n67434 , n67435 , n67436 , n67437 , n67438 , n67439 , n67440 , n67441 , n67442 ,
     n67443 , n67444 , n67445 , n67446 , n67447 , n67448 , n67449 , n67450 , n67451 , n67452 ,
     n67453 , n67454 , n67455 , n67456 , n67457 , n67458 , n67459 , n67460 , n67461 , n67462 ,
     n67463 , n67464 , n67465 , n67466 , n67467 , n67468 , n67469 , n67470 , n67471 , n67472 ,
     n67473 , n67474 , n67475 , n67476 , n67477 , n67478 , n67479 , n67480 , n67481 , n67482 ,
     n67483 , n67484 , n67485 , n67486 , n67487 , n67488 , n67489 , n67490 , n67491 , n67492 ,
     n67493 , n67494 , n67495 , n67496 , n67497 , n67498 , n67499 , n67500 , n67501 , n67502 ,
     n67503 , n67504 , n67505 , n67506 , n67507 , n67508 , n67509 , n67510 , n67511 , n67512 ,
     n67513 , n67514 , n67515 , n67516 , n67517 , n67518 , n67519 , n67520 , n67521 , n67522 ,
     n67523 , n67524 , n67525 , n67526 , n67527 , n67528 , n67529 , n67530 , n67531 , n67532 ,
     n67533 , n67534 , n67535 , n67536 , n67537 , n67538 , n67539 , n67540 , n67541 , n67542 ,
     n67543 , n67544 , n67545 , n67546 , n67547 , n67548 , n67549 , n67550 , n67551 , n67552 ,
     n67553 , n67554 , n67555 , n67556 , n67557 , n67558 , n67559 , n67560 , n67561 , n67562 ,
     n67563 , n67564 , n67565 , n67566 , n67567 , n67568 , n67569 , n67570 , n67571 , n67572 ,
     n67573 , n67574 , n67575 , n67576 , n67577 , n67578 , n67579 , n67580 , n67581 , n67582 ,
     n67583 , n67584 , n67585 , n67586 , n67587 , n67588 , n67589 , n67590 , n67591 , n67592 ,
     n67593 , n67594 , n67595 , n67596 , n67597 , n67598 , n67599 , n67600 , n67601 , n67602 ,
     n67603 , n67604 , n67605 , n67606 , n67607 , n67608 , n67609 , n67610 , n67611 , n67612 ,
     n67613 , n67614 , n67615 , n67616 , n67617 , n67618 , n67619 , n67620 , n67621 , n67622 ,
     n67623 , n67624 , n67625 , n67626 , n67627 , n67628 , n67629 , n67630 , n67631 , n67632 ,
     n67633 , n67634 , n67635 , n67636 , n67637 , n67638 , n67639 , n67640 , n67641 , n67642 ,
     n67643 , n67644 , n67645 , n67646 , n67647 , n67648 , n67649 , n67650 , n67651 , n67652 ,
     n67653 , n67654 , n67655 , n67656 , n67657 , n67658 , n67659 , n67660 , n67661 , n67662 ,
     n67663 , n67664 , n67665 , n67666 , n67667 , n67668 , n67669 , n67670 , n67671 , n67672 ,
     n67673 , n67674 , n67675 , n67676 , n67677 , n67678 , n67679 , n67680 , n67681 , n67682 ,
     n67683 , n67684 , n67685 , n67686 , n67687 , n67688 , n67689 , n67690 , n67691 , n67692 ,
     n67693 , n67694 , n67695 , n67696 , n67697 , n67698 , n67699 , n67700 , n67701 , n67702 ,
     n67703 , n67704 , n67705 , n67706 , n67707 , n67708 , n67709 , n67710 , n67711 , n67712 ,
     n67713 , n67714 , n67715 , n67716 , n67717 , n67718 , n67719 , n67720 , n67721 , n67722 ,
     n67723 , n67724 , n67725 , n67726 , n67727 , n67728 , n67729 , n67730 , n67731 , n67732 ,
     n67733 , n67734 , n67735 , n67736 , n67737 , n67738 , n67739 , n67740 , n67741 , n67742 ,
     n67743 , n67744 , n67745 , n67746 , n67747 , n67748 , n67749 , n67750 , n67751 , n67752 ,
     n67753 , n67754 , n67755 , n67756 , n67757 , n67758 , n67759 , n67760 , n67761 , n67762 ,
     n67763 , n67764 , n67765 , n67766 , n67767 , n67768 , n67769 , n67770 , n67771 , n67772 ,
     n67773 , n67774 , n67775 , n67776 , n67777 , n67778 , n67779 , n67780 , n67781 , n67782 ,
     n67783 , n67784 , n67785 , n67786 , n67787 , n67788 , n67789 , n67790 , n67791 , n67792 ,
     n67793 , n67794 , n67795 , n67796 , n67797 , n67798 , n67799 , n67800 , n67801 , n67802 ,
     n67803 , n67804 , n67805 , n67806 , n67807 , n67808 , n67809 , n67810 , n67811 , n67812 ,
     n67813 , n67814 , n67815 , n67816 , n67817 , n67818 , n67819 , n67820 , n67821 , n67822 ,
     n67823 , n67824 , n67825 , n67826 , n67827 , n67828 , n67829 , n67830 , n67831 , n67832 ,
     n67833 , n67834 , n67835 , n67836 , n67837 , n67838 , n67839 , n67840 , n67841 , n67842 ,
     n67843 , n67844 , n67845 , n67846 , n67847 , n67848 , n67849 , n67850 , n67851 , n67852 ,
     n67853 , n67854 , n67855 , n67856 , n67857 , n67858 , n67859 , n67860 , n67861 , n67862 ,
     n67863 , n67864 , n67865 , n67866 , n67867 , n67868 , n67869 , n67870 , n67871 , n67872 ,
     n67873 , n67874 , n67875 , n67876 , n67877 , n67878 , n67879 , n67880 , n67881 , n67882 ,
     n67883 , n67884 , n67885 , n67886 , n67887 , n67888 , n67889 , n67890 , n67891 , n67892 ,
     n67893 , n67894 , n67895 , n67896 , n67897 , n67898 , n67899 , n67900 , n67901 , n67902 ,
     n67903 , n67904 , n67905 , n67906 , n67907 , n67908 , n67909 , n67910 , n67911 , n67912 ,
     n67913 , n67914 , n67915 , n67916 , n67917 , n67918 , n67919 , n67920 , n67921 , n67922 ,
     n67923 , n67924 , n67925 , n67926 , n67927 , n67928 , n67929 , n67930 , n67931 , n67932 ,
     n67933 , n67934 , n67935 , n67936 , n67937 , n67938 , n67939 , n67940 , n67941 , n67942 ,
     n67943 , n67944 , n67945 , n67946 , n67947 , n67948 , n67949 , n67950 , n67951 , n67952 ,
     n67953 , n67954 , n67955 , n67956 , n67957 , n67958 , n67959 , n67960 , n67961 , n67962 ,
     n67963 , n67964 , n67965 , n67966 , n67967 , n67968 , n67969 , n67970 , n67971 , n67972 ,
     n67973 , n67974 , n67975 , n67976 , n67977 , n67978 , n67979 , n67980 , n67981 , n67982 ,
     n67983 , n67984 , n67985 , n67986 , n67987 , n67988 , n67989 , n67990 , n67991 , n67992 ,
     n67993 , n67994 , n67995 , n67996 , n67997 , n67998 , n67999 , n68000 , n68001 , n68002 ,
     n68003 , n68004 , n68005 , n68006 , n68007 , n68008 , n68009 , n68010 , n68011 , n68012 ,
     n68013 , n68014 , n68015 , n68016 , n68017 , n68018 , n68019 , n68020 , n68021 , n68022 ,
     n68023 , n68024 , n68025 , n68026 , n68027 , n68028 , n68029 , n68030 , n68031 , n68032 ,
     n68033 , n68034 , n68035 , n68036 , n68037 , n68038 , n68039 , n68040 , n68041 , n68042 ,
     n68043 , n68044 , n68045 , n68046 , n68047 , n68048 , n68049 , n68050 , n68051 , n68052 ,
     n68053 , n68054 , n68055 , n68056 , n68057 , n68058 , n68059 , n68060 , n68061 , n68062 ,
     n68063 , n68064 , n68065 , n68066 , n68067 , n68068 , n68069 , n68070 , n68071 , n68072 ,
     n68073 , n68074 , n68075 , n68076 , n68077 , n68078 , n68079 , n68080 , n68081 , n68082 ,
     n68083 , n68084 , n68085 , n68086 , n68087 , n68088 , n68089 , n68090 , n68091 , n68092 ,
     n68093 , n68094 , n68095 , n68096 , n68097 , n68098 , n68099 , n68100 , n68101 , n68102 ,
     n68103 , n68104 , n68105 , n68106 , n68107 , n68108 , n68109 , n68110 , n68111 , n68112 ,
     n68113 , n68114 , n68115 , n68116 , n68117 , n68118 , n68119 , n68120 , n68121 , n68122 ,
     n68123 , n68124 , n68125 , n68126 , n68127 , n68128 , n68129 , n68130 , n68131 , n68132 ,
     n68133 , n68134 , n68135 , n68136 , n68137 , n68138 , n68139 , n68140 , n68141 , n68142 ,
     n68143 , n68144 , n68145 , n68146 , n68147 , n68148 , n68149 , n68150 , n68151 , n68152 ,
     n68153 , n68154 , n68155 , n68156 , n68157 , n68158 , n68159 , n68160 , n68161 , n68162 ,
     n68163 , n68164 , n68165 , n68166 , n68167 , n68168 , n68169 , n68170 , n68171 , n68172 ,
     n68173 , n68174 , n68175 , n68176 , n68177 , n68178 , n68179 , n68180 , n68181 , n68182 ,
     n68183 , n68184 , n68185 , n68186 , n68187 , n68188 , n68189 , n68190 , n68191 , n68192 ,
     n68193 , n68194 , n68195 , n68196 , n68197 , n68198 , n68199 , n68200 , n68201 , n68202 ,
     n68203 , n68204 , n68205 , n68206 , n68207 , n68208 , n68209 , n68210 , n68211 , n68212 ,
     n68213 , n68214 , n68215 , n68216 , n68217 , n68218 , n68219 , n68220 , n68221 , n68222 ,
     n68223 , n68224 , n68225 , n68226 , n68227 , n68228 , n68229 , n68230 , n68231 , n68232 ,
     n68233 , n68234 , n68235 , n68236 , n68237 , n68238 , n68239 , n68240 , n68241 , n68242 ,
     n68243 , n68244 , n68245 , n68246 , n68247 , n68248 , n68249 , n68250 , n68251 , n68252 ,
     n68253 , n68254 , n68255 , n68256 , n68257 , n68258 , n68259 , n68260 , n68261 , n68262 ,
     n68263 , n68264 , n68265 , n68266 , n68267 , n68268 , n68269 , n68270 , n68271 , n68272 ,
     n68273 , n68274 , n68275 , n68276 , n68277 , n68278 , n68279 , n68280 , n68281 , n68282 ,
     n68283 , n68284 , n68285 , n68286 , n68287 , n68288 , n68289 , n68290 , n68291 , n68292 ,
     n68293 , n68294 , n68295 , n68296 , n68297 , n68298 , n68299 , n68300 , n68301 , n68302 ,
     n68303 , n68304 , n68305 , n68306 , n68307 , n68308 , n68309 , n68310 , n68311 , n68312 ,
     n68313 , n68314 , n68315 , n68316 , n68317 , n68318 , n68319 , n68320 , n68321 , n68322 ,
     n68323 , n68324 , n68325 , n68326 , n68327 , n68328 , n68329 , n68330 , n68331 , n68332 ,
     n68333 , n68334 , n68335 , n68336 , n68337 , n68338 , n68339 , n68340 , n68341 , n68342 ,
     n68343 , n68344 , n68345 , n68346 , n68347 , n68348 , n68349 , n68350 , n68351 , n68352 ,
     n68353 , n68354 , n68355 , n68356 , n68357 , n68358 , n68359 , n68360 , n68361 , n68362 ,
     n68363 , n68364 , n68365 , n68366 , n68367 , n68368 , n68369 , n68370 , n68371 , n68372 ,
     n68373 , n68374 , n68375 , n68376 , n68377 , n68378 , n68379 , n68380 , n68381 , n68382 ,
     n68383 , n68384 , n68385 , n68386 , n68387 , n68388 , n68389 , n68390 , n68391 , n68392 ,
     n68393 , n68394 , n68395 , n68396 , n68397 , n68398 , n68399 , n68400 , n68401 , n68402 ,
     n68403 , n68404 , n68405 , n68406 , n68407 , n68408 , n68409 , n68410 , n68411 , n68412 ,
     n68413 , n68414 , n68415 , n68416 , n68417 , n68418 , n68419 , n68420 , n68421 , n68422 ,
     n68423 , n68424 , n68425 , n68426 , n68427 , n68428 , n68429 , n68430 , n68431 , n68432 ,
     n68433 , n68434 , n68435 , n68436 , n68437 , n68438 , n68439 , n68440 , n68441 , n68442 ,
     n68443 , n68444 , n68445 , n68446 , n68447 , n68448 , n68449 , n68450 , n68451 , n68452 ,
     n68453 , n68454 , n68455 , n68456 , n68457 , n68458 , n68459 , n68460 , n68461 , n68462 ,
     n68463 , n68464 , n68465 , n68466 , n68467 , n68468 , n68469 , n68470 , n68471 , n68472 ,
     n68473 , n68474 , n68475 , n68476 , n68477 , n68478 , n68479 , n68480 , n68481 , n68482 ,
     n68483 , n68484 , n68485 , n68486 , n68487 , n68488 , n68489 , n68490 , n68491 , n68492 ,
     n68493 , n68494 , n68495 , n68496 , n68497 , n68498 , n68499 , n68500 , n68501 , n68502 ,
     n68503 , n68504 , n68505 , n68506 , n68507 , n68508 , n68509 , n68510 , n68511 , n68512 ,
     n68513 , n68514 , n68515 , n68516 , n68517 , n68518 , n68519 , n68520 , n68521 , n68522 ,
     n68523 , n68524 , n68525 , n68526 , n68527 , n68528 , n68529 , n68530 , n68531 , n68532 ,
     n68533 , n68534 , n68535 , n68536 , n68537 , n68538 , n68539 , n68540 , n68541 , n68542 ,
     n68543 , n68544 , n68545 , n68546 , n68547 , n68548 , n68549 , n68550 , n68551 , n68552 ,
     n68553 , n68554 , n68555 , n68556 , n68557 , n68558 , n68559 , n68560 , n68561 , n68562 ,
     n68563 , n68564 , n68565 , n68566 , n68567 , n68568 , n68569 , n68570 , n68571 , n68572 ,
     n68573 , n68574 , n68575 , n68576 , n68577 , n68578 , n68579 , n68580 , n68581 , n68582 ,
     n68583 , n68584 , n68585 , n68586 , n68587 , n68588 , n68589 , n68590 , n68591 , n68592 ,
     n68593 , n68594 , n68595 , n68596 , n68597 , n68598 , n68599 , n68600 , n68601 , n68602 ,
     n68603 , n68604 , n68605 , n68606 , n68607 , n68608 , n68609 , n68610 , n68611 , n68612 ,
     n68613 , n68614 , n68615 , n68616 , n68617 , n68618 , n68619 , n68620 , n68621 , n68622 ,
     n68623 , n68624 , n68625 , n68626 , n68627 , n68628 , n68629 , n68630 , n68631 , n68632 ,
     n68633 , n68634 , n68635 , n68636 , n68637 , n68638 , n68639 , n68640 , n68641 , n68642 ,
     n68643 , n68644 , n68645 , n68646 , n68647 , n68648 , n68649 , n68650 , n68651 , n68652 ,
     n68653 , n68654 , n68655 , n68656 , n68657 , n68658 , n68659 , n68660 , n68661 , n68662 ,
     n68663 , n68664 , n68665 , n68666 , n68667 , n68668 , n68669 , n68670 , n68671 , n68672 ,
     n68673 , n68674 , n68675 , n68676 , n68677 , n68678 , n68679 , n68680 , n68681 , n68682 ,
     n68683 , n68684 , n68685 , n68686 , n68687 , n68688 , n68689 , n68690 , n68691 , n68692 ,
     n68693 , n68694 , n68695 , n68696 , n68697 , n68698 , n68699 , n68700 , n68701 , n68702 ,
     n68703 , n68704 , n68705 , n68706 , n68707 , n68708 , n68709 , n68710 , n68711 , n68712 ,
     n68713 , n68714 , n68715 , n68716 , n68717 , n68718 , n68719 , n68720 , n68721 , n68722 ,
     n68723 , n68724 , n68725 , n68726 , n68727 , n68728 , n68729 , n68730 , n68731 , n68732 ,
     n68733 , n68734 , n68735 , n68736 , n68737 , n68738 , n68739 , n68740 , n68741 , n68742 ,
     n68743 , n68744 , n68745 , n68746 , n68747 , n68748 , n68749 , n68750 , n68751 , n68752 ,
     n68753 , n68754 , n68755 , n68756 , n68757 , n68758 , n68759 , n68760 , n68761 , n68762 ,
     n68763 , n68764 , n68765 , n68766 , n68767 , n68768 , n68769 , n68770 , n68771 , n68772 ,
     n68773 , n68774 , n68775 , n68776 , n68777 , n68778 , n68779 , n68780 , n68781 , n68782 ,
     n68783 , n68784 , n68785 , n68786 , n68787 , n68788 , n68789 , n68790 , n68791 , n68792 ,
     n68793 , n68794 , n68795 , n68796 , n68797 , n68798 , n68799 , n68800 , n68801 , n68802 ,
     n68803 , n68804 , n68805 , n68806 , n68807 , n68808 , n68809 , n68810 , n68811 , n68812 ,
     n68813 , n68814 , n68815 , n68816 , n68817 , n68818 , n68819 , n68820 , n68821 , n68822 ,
     n68823 , n68824 , n68825 , n68826 , n68827 , n68828 , n68829 , n68830 , n68831 , n68832 ,
     n68833 , n68834 , n68835 , n68836 , n68837 , n68838 , n68839 , n68840 , n68841 , n68842 ,
     n68843 , n68844 , n68845 , n68846 , n68847 , n68848 , n68849 , n68850 , n68851 , n68852 ,
     n68853 , n68854 , n68855 , n68856 , n68857 , n68858 , n68859 , n68860 , n68861 , n68862 ,
     n68863 , n68864 , n68865 , n68866 , n68867 , n68868 , n68869 , n68870 , n68871 , n68872 ,
     n68873 , n68874 , n68875 , n68876 , n68877 , n68878 , n68879 , n68880 , n68881 , n68882 ,
     n68883 , n68884 , n68885 , n68886 , n68887 , n68888 , n68889 , n68890 , n68891 , n68892 ,
     n68893 , n68894 , n68895 , n68896 , n68897 , n68898 , n68899 , n68900 , n68901 , n68902 ,
     n68903 , n68904 , n68905 , n68906 , n68907 , n68908 , n68909 , n68910 , n68911 , n68912 ,
     n68913 , n68914 , n68915 , n68916 , n68917 , n68918 , n68919 , n68920 , n68921 , n68922 ,
     n68923 , n68924 , n68925 , n68926 , n68927 , n68928 , n68929 , n68930 , n68931 , n68932 ,
     n68933 , n68934 , n68935 , n68936 , n68937 , n68938 , n68939 , n68940 , n68941 , n68942 ,
     n68943 , n68944 , n68945 , n68946 , n68947 , n68948 , n68949 , n68950 , n68951 , n68952 ,
     n68953 , n68954 , n68955 , n68956 , n68957 , n68958 , n68959 , n68960 , n68961 , n68962 ,
     n68963 , n68964 , n68965 , n68966 , n68967 , n68968 , n68969 , n68970 , n68971 , n68972 ,
     n68973 , n68974 , n68975 , n68976 , n68977 , n68978 , n68979 , n68980 , n68981 , n68982 ,
     n68983 , n68984 , n68985 , n68986 , n68987 , n68988 , n68989 , n68990 , n68991 , n68992 ,
     n68993 , n68994 , n68995 , n68996 , n68997 , n68998 , n68999 , n69000 , n69001 , n69002 ,
     n69003 , n69004 , n69005 , n69006 , n69007 , n69008 , n69009 , n69010 , n69011 , n69012 ,
     n69013 , n69014 , n69015 , n69016 , n69017 , n69018 , n69019 , n69020 , n69021 , n69022 ,
     n69023 , n69024 , n69025 , n69026 , n69027 , n69028 , n69029 , n69030 , n69031 , n69032 ,
     n69033 , n69034 , n69035 , n69036 , n69037 , n69038 , n69039 , n69040 , n69041 , n69042 ,
     n69043 , n69044 , n69045 , n69046 , n69047 , n69048 , n69049 , n69050 , n69051 , n69052 ,
     n69053 , n69054 , n69055 , n69056 , n69057 , n69058 , n69059 , n69060 , n69061 , n69062 ,
     n69063 , n69064 , n69065 , n69066 , n69067 , n69068 , n69069 , n69070 , n69071 , n69072 ,
     n69073 , n69074 , n69075 , n69076 , n69077 , n69078 , n69079 , n69080 , n69081 , n69082 ,
     n69083 , n69084 , n69085 , n69086 , n69087 , n69088 , n69089 , n69090 , n69091 , n69092 ,
     n69093 , n69094 , n69095 , n69096 , n69097 , n69098 , n69099 , n69100 , n69101 , n69102 ,
     n69103 , n69104 , n69105 , n69106 , n69107 , n69108 , n69109 , n69110 , n69111 , n69112 ,
     n69113 , n69114 , n69115 , n69116 , n69117 , n69118 , n69119 , n69120 , n69121 , n69122 ,
     n69123 , n69124 , n69125 , n69126 , n69127 , n69128 , n69129 , n69130 , n69131 , n69132 ,
     n69133 , n69134 , n69135 , n69136 , n69137 , n69138 , n69139 , n69140 , n69141 , n69142 ,
     n69143 , n69144 , n69145 , n69146 , n69147 , n69148 , n69149 , n69150 , n69151 , n69152 ,
     n69153 , n69154 , n69155 , n69156 , n69157 , n69158 , n69159 , n69160 , n69161 , n69162 ,
     n69163 , n69164 , n69165 , n69166 , n69167 , n69168 , n69169 , n69170 , n69171 , n69172 ,
     n69173 , n69174 , n69175 , n69176 , n69177 , n69178 , n69179 , n69180 , n69181 , n69182 ,
     n69183 , n69184 , n69185 , n69186 , n69187 , n69188 , n69189 , n69190 , n69191 , n69192 ,
     n69193 , n69194 , n69195 , n69196 , n69197 , n69198 , n69199 , n69200 , n69201 , n69202 ,
     n69203 , n69204 , n69205 , n69206 , n69207 , n69208 , n69209 , n69210 , n69211 , n69212 ,
     n69213 , n69214 , n69215 , n69216 , n69217 , n69218 , n69219 , n69220 , n69221 , n69222 ,
     n69223 , n69224 , n69225 , n69226 , n69227 , n69228 , n69229 , n69230 , n69231 , n69232 ,
     n69233 , n69234 , n69235 , n69236 , n69237 , n69238 , n69239 , n69240 , n69241 , n69242 ,
     n69243 , n69244 , n69245 , n69246 , n69247 , n69248 , n69249 , n69250 , n69251 , n69252 ,
     n69253 , n69254 , n69255 , n69256 , n69257 , n69258 , n69259 , n69260 , n69261 , n69262 ,
     n69263 , n69264 , n69265 , n69266 , n69267 , n69268 , n69269 , n69270 , n69271 , n69272 ,
     n69273 , n69274 , n69275 , n69276 , n69277 , n69278 , n69279 , n69280 , n69281 , n69282 ,
     n69283 , n69284 , n69285 , n69286 , n69287 , n69288 , n69289 , n69290 , n69291 , n69292 ,
     n69293 , n69294 , n69295 , n69296 , n69297 , n69298 , n69299 , n69300 , n69301 , n69302 ,
     n69303 , n69304 , n69305 , n69306 , n69307 , n69308 , n69309 , n69310 , n69311 , n69312 ,
     n69313 , n69314 , n69315 , n69316 , n69317 , n69318 , n69319 , n69320 , n69321 , n69322 ,
     n69323 , n69324 , n69325 , n69326 , n69327 , n69328 , n69329 , n69330 , n69331 , n69332 ,
     n69333 , n69334 , n69335 , n69336 , n69337 , n69338 , n69339 , n69340 , n69341 , n69342 ,
     n69343 , n69344 , n69345 , n69346 , n69347 , n69348 , n69349 , n69350 , n69351 , n69352 ,
     n69353 , n69354 , n69355 , n69356 , n69357 , n69358 , n69359 , n69360 , n69361 , n69362 ,
     n69363 , n69364 , n69365 , n69366 , n69367 , n69368 , n69369 , n69370 , n69371 , n69372 ,
     n69373 , n69374 , n69375 , n69376 , n69377 , n69378 , n69379 , n69380 , n69381 , n69382 ,
     n69383 , n69384 , n69385 , n69386 , n69387 , n69388 , n69389 , n69390 , n69391 , n69392 ,
     n69393 , n69394 , n69395 , n69396 , n69397 , n69398 , n69399 , n69400 , n69401 , n69402 ,
     n69403 , n69404 , n69405 , n69406 , n69407 , n69408 , n69409 , n69410 , n69411 , n69412 ,
     n69413 , n69414 , n69415 , n69416 , n69417 , n69418 , n69419 , n69420 , n69421 , n69422 ,
     n69423 , n69424 , n69425 , n69426 , n69427 , n69428 , n69429 , n69430 , n69431 , n69432 ,
     n69433 , n69434 , n69435 , n69436 , n69437 , n69438 , n69439 , n69440 , n69441 , n69442 ,
     n69443 , n69444 , n69445 , n69446 , n69447 , n69448 , n69449 , n69450 , n69451 , n69452 ,
     n69453 , n69454 , n69455 , n69456 , n69457 , n69458 , n69459 , n69460 , n69461 , n69462 ,
     n69463 , n69464 , n69465 , n69466 , n69467 , n69468 , n69469 , n69470 , n69471 , n69472 ,
     n69473 , n69474 , n69475 , n69476 , n69477 , n69478 , n69479 , n69480 , n69481 , n69482 ,
     n69483 , n69484 , n69485 , n69486 , n69487 , n69488 , n69489 , n69490 , n69491 , n69492 ,
     n69493 , n69494 , n69495 , n69496 , n69497 , n69498 , n69499 , n69500 , n69501 , n69502 ,
     n69503 , n69504 , n69505 , n69506 , n69507 , n69508 , n69509 , n69510 , n69511 , n69512 ,
     n69513 , n69514 , n69515 , n69516 , n69517 , n69518 , n69519 , n69520 , n69521 , n69522 ,
     n69523 , n69524 , n69525 , n69526 , n69527 , n69528 , n69529 , n69530 , n69531 , n69532 ,
     n69533 , n69534 , n69535 , n69536 , n69537 , n69538 , n69539 , n69540 , n69541 , n69542 ,
     n69543 , n69544 , n69545 , n69546 , n69547 , n69548 , n69549 , n69550 , n69551 , n69552 ,
     n69553 , n69554 , n69555 , n69556 , n69557 , n69558 , n69559 , n69560 , n69561 , n69562 ,
     n69563 , n69564 , n69565 , n69566 , n69567 , n69568 , n69569 , n69570 , n69571 , n69572 ,
     n69573 , n69574 , n69575 , n69576 , n69577 , n69578 , n69579 , n69580 , n69581 , n69582 ,
     n69583 , n69584 , n69585 , n69586 , n69587 , n69588 , n69589 , n69590 , n69591 , n69592 ,
     n69593 , n69594 , n69595 , n69596 , n69597 , n69598 , n69599 , n69600 , n69601 , n69602 ,
     n69603 , n69604 , n69605 , n69606 , n69607 , n69608 , n69609 , n69610 , n69611 , n69612 ,
     n69613 , n69614 , n69615 , n69616 , n69617 , n69618 , n69619 , n69620 , n69621 , n69622 ,
     n69623 , n69624 , n69625 , n69626 , n69627 , n69628 , n69629 , n69630 , n69631 , n69632 ,
     n69633 , n69634 , n69635 , n69636 , n69637 , n69638 , n69639 , n69640 , n69641 , n69642 ,
     n69643 , n69644 , n69645 , n69646 , n69647 , n69648 , n69649 , n69650 , n69651 , n69652 ,
     n69653 , n69654 , n69655 , n69656 , n69657 , n69658 , n69659 , n69660 , n69661 , n69662 ,
     n69663 , n69664 , n69665 , n69666 , n69667 , n69668 , n69669 , n69670 , n69671 , n69672 ,
     n69673 , n69674 , n69675 , n69676 , n69677 , n69678 , n69679 , n69680 , n69681 , n69682 ,
     n69683 , n69684 , n69685 , n69686 , n69687 , n69688 , n69689 , n69690 , n69691 , n69692 ,
     n69693 , n69694 , n69695 , n69696 , n69697 , n69698 , n69699 , n69700 , n69701 , n69702 ,
     n69703 , n69704 , n69705 , n69706 , n69707 , n69708 , n69709 , n69710 , n69711 , n69712 ,
     n69713 , n69714 , n69715 , n69716 , n69717 , n69718 , n69719 , n69720 , n69721 , n69722 ,
     n69723 , n69724 , n69725 , n69726 , n69727 , n69728 , n69729 , n69730 , n69731 , n69732 ,
     n69733 , n69734 , n69735 , n69736 , n69737 , n69738 , n69739 , n69740 , n69741 , n69742 ,
     n69743 , n69744 , n69745 , n69746 , n69747 , n69748 , n69749 , n69750 , n69751 , n69752 ,
     n69753 , n69754 , n69755 , n69756 , n69757 , n69758 , n69759 , n69760 , n69761 , n69762 ,
     n69763 , n69764 , n69765 , n69766 , n69767 , n69768 , n69769 , n69770 , n69771 , n69772 ,
     n69773 , n69774 , n69775 , n69776 , n69777 , n69778 , n69779 , n69780 , n69781 , n69782 ,
     n69783 , n69784 , n69785 , n69786 , n69787 , n69788 , n69789 , n69790 , n69791 , n69792 ,
     n69793 , n69794 , n69795 , n69796 , n69797 , n69798 , n69799 , n69800 , n69801 , n69802 ,
     n69803 , n69804 , n69805 , n69806 , n69807 , n69808 , n69809 , n69810 , n69811 , n69812 ,
     n69813 , n69814 , n69815 , n69816 , n69817 , n69818 , n69819 , n69820 , n69821 , n69822 ,
     n69823 , n69824 , n69825 , n69826 , n69827 , n69828 , n69829 , n69830 , n69831 , n69832 ,
     n69833 , n69834 , n69835 , n69836 , n69837 , n69838 , n69839 , n69840 , n69841 , n69842 ,
     n69843 , n69844 , n69845 , n69846 , n69847 , n69848 , n69849 , n69850 , n69851 , n69852 ,
     n69853 , n69854 , n69855 , n69856 , n69857 , n69858 , n69859 , n69860 , n69861 , n69862 ,
     n69863 , n69864 , n69865 , n69866 , n69867 , n69868 , n69869 , n69870 , n69871 , n69872 ,
     n69873 , n69874 , n69875 , n69876 , n69877 , n69878 , n69879 , n69880 , n69881 , n69882 ,
     n69883 , n69884 , n69885 , n69886 , n69887 , n69888 , n69889 , n69890 , n69891 , n69892 ,
     n69893 , n69894 , n69895 , n69896 , n69897 , n69898 , n69899 , n69900 , n69901 , n69902 ,
     n69903 , n69904 , n69905 , n69906 , n69907 , n69908 , n69909 , n69910 , n69911 , n69912 ,
     n69913 , n69914 , n69915 , n69916 , n69917 , n69918 , n69919 , n69920 , n69921 , n69922 ,
     n69923 , n69924 , n69925 , n69926 , n69927 , n69928 , n69929 , n69930 , n69931 , n69932 ,
     n69933 , n69934 , n69935 , n69936 , n69937 , n69938 , n69939 , n69940 , n69941 , n69942 ,
     n69943 , n69944 , n69945 , n69946 , n69947 , n69948 , n69949 , n69950 , n69951 , n69952 ,
     n69953 , n69954 , n69955 , n69956 , n69957 , n69958 , n69959 , n69960 , n69961 , n69962 ,
     n69963 , n69964 , n69965 , n69966 , n69967 , n69968 , n69969 , n69970 , n69971 , n69972 ,
     n69973 , n69974 , n69975 , n69976 , n69977 , n69978 , n69979 , n69980 , n69981 , n69982 ,
     n69983 , n69984 , n69985 , n69986 , n69987 , n69988 , n69989 , n69990 , n69991 , n69992 ,
     n69993 , n69994 , n69995 , n69996 , n69997 , n69998 , n69999 , n70000 , n70001 , n70002 ,
     n70003 , n70004 , n70005 , n70006 , n70007 , n70008 , n70009 , n70010 , n70011 , n70012 ,
     n70013 , n70014 , n70015 , n70016 , n70017 , n70018 , n70019 , n70020 , n70021 , n70022 ,
     n70023 , n70024 , n70025 , n70026 , n70027 , n70028 , n70029 , n70030 , n70031 , n70032 ,
     n70033 , n70034 , n70035 , n70036 , n70037 , n70038 , n70039 , n70040 , n70041 , n70042 ,
     n70043 , n70044 , n70045 , n70046 , n70047 , n70048 , n70049 , n70050 , n70051 , n70052 ,
     n70053 , n70054 , n70055 , n70056 , n70057 , n70058 , n70059 , n70060 , n70061 , n70062 ,
     n70063 , n70064 , n70065 , n70066 , n70067 , n70068 , n70069 , n70070 , n70071 , n70072 ,
     n70073 , n70074 , n70075 , n70076 , n70077 , n70078 , n70079 , n70080 , n70081 , n70082 ,
     n70083 , n70084 , n70085 , n70086 , n70087 , n70088 , n70089 , n70090 , n70091 , n70092 ,
     n70093 , n70094 , n70095 , n70096 , n70097 , n70098 , n70099 , n70100 , n70101 , n70102 ,
     n70103 , n70104 , n70105 , n70106 , n70107 , n70108 , n70109 , n70110 , n70111 , n70112 ,
     n70113 , n70114 , n70115 , n70116 , n70117 , n70118 , n70119 , n70120 , n70121 , n70122 ,
     n70123 , n70124 , n70125 , n70126 , n70127 , n70128 , n70129 , n70130 , n70131 , n70132 ,
     n70133 , n70134 , n70135 , n70136 , n70137 , n70138 , n70139 , n70140 , n70141 , n70142 ,
     n70143 , n70144 , n70145 , n70146 , n70147 , n70148 , n70149 , n70150 , n70151 , n70152 ,
     n70153 , n70154 , n70155 , n70156 , n70157 , n70158 , n70159 , n70160 , n70161 , n70162 ,
     n70163 , n70164 , n70165 , n70166 , n70167 , n70168 , n70169 , n70170 , n70171 , n70172 ,
     n70173 , n70174 , n70175 , n70176 , n70177 , n70178 , n70179 , n70180 , n70181 , n70182 ,
     n70183 , n70184 , n70185 , n70186 , n70187 , n70188 , n70189 , n70190 , n70191 , n70192 ,
     n70193 , n70194 , n70195 , n70196 , n70197 , n70198 , n70199 , n70200 , n70201 , n70202 ,
     n70203 , n70204 , n70205 , n70206 , n70207 , n70208 , n70209 , n70210 , n70211 , n70212 ,
     n70213 , n70214 , n70215 , n70216 , n70217 , n70218 , n70219 , n70220 , n70221 , n70222 ,
     n70223 , n70224 , n70225 , n70226 , n70227 , n70228 , n70229 , n70230 , n70231 , n70232 ,
     n70233 , n70234 , n70235 , n70236 , n70237 , n70238 , n70239 , n70240 , n70241 , n70242 ,
     n70243 , n70244 , n70245 , n70246 , n70247 , n70248 , n70249 , n70250 , n70251 , n70252 ,
     n70253 , n70254 , n70255 , n70256 , n70257 , n70258 , n70259 , n70260 , n70261 , n70262 ,
     n70263 , n70264 , n70265 , n70266 , n70267 , n70268 , n70269 , n70270 , n70271 , n70272 ,
     n70273 , n70274 , n70275 , n70276 , n70277 , n70278 , n70279 , n70280 , n70281 , n70282 ,
     n70283 , n70284 , n70285 , n70286 , n70287 , n70288 , n70289 , n70290 , n70291 , n70292 ,
     n70293 , n70294 , n70295 , n70296 , n70297 , n70298 , n70299 , n70300 , n70301 , n70302 ,
     n70303 , n70304 , n70305 , n70306 , n70307 , n70308 , n70309 , n70310 , n70311 , n70312 ,
     n70313 , n70314 , n70315 , n70316 , n70317 , n70318 , n70319 , n70320 , n70321 , n70322 ,
     n70323 , n70324 , n70325 , n70326 , n70327 , n70328 , n70329 , n70330 , n70331 , n70332 ,
     n70333 , n70334 , n70335 , n70336 , n70337 , n70338 , n70339 , n70340 , n70341 , n70342 ,
     n70343 , n70344 , n70345 , n70346 , n70347 , n70348 , n70349 , n70350 , n70351 , n70352 ,
     n70353 , n70354 , n70355 , n70356 , n70357 , n70358 , n70359 , n70360 , n70361 , n70362 ,
     n70363 , n70364 , n70365 , n70366 , n70367 , n70368 , n70369 , n70370 , n70371 , n70372 ,
     n70373 , n70374 , n70375 , n70376 , n70377 , n70378 , n70379 , n70380 , n70381 , n70382 ,
     n70383 , n70384 , n70385 , n70386 , n70387 , n70388 , n70389 , n70390 , n70391 , n70392 ,
     n70393 , n70394 , n70395 , n70396 , n70397 , n70398 , n70399 , n70400 , n70401 , n70402 ,
     n70403 , n70404 , n70405 , n70406 , n70407 , n70408 , n70409 , n70410 , n70411 , n70412 ,
     n70413 , n70414 , n70415 , n70416 , n70417 , n70418 , n70419 , n70420 , n70421 , n70422 ,
     n70423 , n70424 , n70425 , n70426 , n70427 , n70428 , n70429 , n70430 , n70431 , n70432 ,
     n70433 , n70434 , n70435 , n70436 , n70437 , n70438 , n70439 , n70440 , n70441 , n70442 ,
     n70443 , n70444 , n70445 , n70446 , n70447 , n70448 , n70449 , n70450 , n70451 , n70452 ,
     n70453 , n70454 , n70455 , n70456 , n70457 , n70458 , n70459 , n70460 , n70461 , n70462 ,
     n70463 , n70464 , n70465 , n70466 , n70467 , n70468 , n70469 , n70470 , n70471 , n70472 ,
     n70473 , n70474 , n70475 , n70476 , n70477 , n70478 , n70479 , n70480 , n70481 , n70482 ,
     n70483 , n70484 , n70485 , n70486 , n70487 , n70488 , n70489 , n70490 , n70491 , n70492 ,
     n70493 , n70494 , n70495 , n70496 , n70497 , n70498 , n70499 , n70500 , n70501 , n70502 ,
     n70503 , n70504 , n70505 , n70506 , n70507 , n70508 , n70509 , n70510 , n70511 , n70512 ,
     n70513 , n70514 , n70515 , n70516 , n70517 , n70518 , n70519 , n70520 , n70521 , n70522 ,
     n70523 , n70524 , n70525 , n70526 , n70527 , n70528 , n70529 , n70530 , n70531 , n70532 ,
     n70533 , n70534 , n70535 , n70536 , n70537 , n70538 , n70539 , n70540 , n70541 , n70542 ,
     n70543 , n70544 , n70545 , n70546 , n70547 , n70548 , n70549 , n70550 , n70551 , n70552 ,
     n70553 , n70554 , n70555 , n70556 , n70557 , n70558 , n70559 , n70560 , n70561 , n70562 ,
     n70563 , n70564 , n70565 , n70566 , n70567 , n70568 , n70569 , n70570 , n70571 , n70572 ,
     n70573 , n70574 , n70575 , n70576 , n70577 , n70578 , n70579 , n70580 , n70581 , n70582 ,
     n70583 , n70584 , n70585 , n70586 , n70587 , n70588 , n70589 , n70590 , n70591 , n70592 ,
     n70593 , n70594 , n70595 , n70596 , n70597 , n70598 , n70599 , n70600 , n70601 , n70602 ,
     n70603 , n70604 , n70605 , n70606 , n70607 , n70608 , n70609 , n70610 , n70611 , n70612 ,
     n70613 , n70614 , n70615 , n70616 , n70617 , n70618 , n70619 , n70620 , n70621 , n70622 ,
     n70623 , n70624 , n70625 , n70626 , n70627 , n70628 , n70629 , n70630 , n70631 , n70632 ,
     n70633 , n70634 , n70635 , n70636 , n70637 , n70638 , n70639 , n70640 , n70641 , n70642 ,
     n70643 , n70644 , n70645 , n70646 , n70647 , n70648 , n70649 , n70650 , n70651 , n70652 ,
     n70653 , n70654 , n70655 , n70656 , n70657 , n70658 , n70659 , n70660 , n70661 , n70662 ,
     n70663 , n70664 , n70665 , n70666 , n70667 , n70668 , n70669 , n70670 , n70671 , n70672 ,
     n70673 , n70674 , n70675 , n70676 , n70677 , n70678 , n70679 , n70680 , n70681 , n70682 ,
     n70683 , n70684 , n70685 , n70686 , n70687 , n70688 , n70689 , n70690 , n70691 , n70692 ,
     n70693 , n70694 , n70695 , n70696 , n70697 , n70698 , n70699 , n70700 , n70701 , n70702 ,
     n70703 , n70704 , n70705 , n70706 , n70707 , n70708 , n70709 , n70710 , n70711 , n70712 ,
     n70713 , n70714 , n70715 , n70716 , n70717 , n70718 , n70719 , n70720 , n70721 , n70722 ,
     n70723 , n70724 , n70725 , n70726 , n70727 , n70728 , n70729 , n70730 , n70731 , n70732 ,
     n70733 , n70734 , n70735 , n70736 , n70737 , n70738 , n70739 , n70740 , n70741 , n70742 ,
     n70743 , n70744 , n70745 , n70746 , n70747 , n70748 , n70749 , n70750 , n70751 , n70752 ,
     n70753 , n70754 , n70755 , n70756 , n70757 , n70758 , n70759 , n70760 , n70761 , n70762 ,
     n70763 , n70764 , n70765 , n70766 , n70767 , n70768 , n70769 , n70770 , n70771 , n70772 ,
     n70773 , n70774 , n70775 , n70776 , n70777 , n70778 , n70779 , n70780 , n70781 , n70782 ,
     n70783 , n70784 , n70785 , n70786 , n70787 , n70788 , n70789 , n70790 , n70791 , n70792 ,
     n70793 , n70794 , n70795 , n70796 , n70797 , n70798 , n70799 , n70800 , n70801 , n70802 ,
     n70803 , n70804 , n70805 , n70806 , n70807 , n70808 , n70809 , n70810 , n70811 , n70812 ,
     n70813 , n70814 , n70815 , n70816 , n70817 , n70818 , n70819 , n70820 , n70821 , n70822 ,
     n70823 , n70824 , n70825 , n70826 , n70827 , n70828 , n70829 , n70830 , n70831 , n70832 ,
     n70833 , n70834 , n70835 , n70836 , n70837 , n70838 , n70839 , n70840 , n70841 , n70842 ,
     n70843 , n70844 , n70845 , n70846 , n70847 , n70848 , n70849 , n70850 , n70851 , n70852 ,
     n70853 , n70854 , n70855 , n70856 , n70857 , n70858 , n70859 , n70860 , n70861 , n70862 ,
     n70863 , n70864 , n70865 , n70866 , n70867 , n70868 , n70869 , n70870 , n70871 , n70872 ,
     n70873 , n70874 , n70875 , n70876 , n70877 , n70878 , n70879 , n70880 , n70881 , n70882 ,
     n70883 , n70884 , n70885 , n70886 , n70887 , n70888 , n70889 , n70890 , n70891 , n70892 ,
     n70893 , n70894 , n70895 , n70896 , n70897 , n70898 , n70899 , n70900 , n70901 , n70902 ,
     n70903 , n70904 , n70905 , n70906 , n70907 , n70908 , n70909 , n70910 , n70911 , n70912 ,
     n70913 , n70914 , n70915 , n70916 , n70917 , n70918 , n70919 , n70920 , n70921 , n70922 ,
     n70923 , n70924 , n70925 , n70926 , n70927 , n70928 , n70929 , n70930 , n70931 , n70932 ,
     n70933 , n70934 , n70935 , n70936 , n70937 , n70938 , n70939 , n70940 , n70941 , n70942 ,
     n70943 , n70944 , n70945 , n70946 , n70947 , n70948 , n70949 , n70950 , n70951 , n70952 ,
     n70953 , n70954 , n70955 , n70956 , n70957 , n70958 , n70959 , n70960 , n70961 , n70962 ,
     n70963 , n70964 , n70965 , n70966 , n70967 , n70968 , n70969 , n70970 , n70971 , n70972 ,
     n70973 , n70974 , n70975 , n70976 , n70977 , n70978 , n70979 , n70980 , n70981 , n70982 ,
     n70983 , n70984 , n70985 , n70986 , n70987 , n70988 , n70989 , n70990 , n70991 , n70992 ,
     n70993 , n70994 , n70995 , n70996 , n70997 , n70998 , n70999 , n71000 , n71001 , n71002 ,
     n71003 , n71004 , n71005 , n71006 , n71007 , n71008 , n71009 , n71010 , n71011 , n71012 ,
     n71013 , n71014 , n71015 , n71016 , n71017 , n71018 , n71019 , n71020 , n71021 , n71022 ,
     n71023 , n71024 , n71025 , n71026 , n71027 , n71028 , n71029 , n71030 , n71031 , n71032 ,
     n71033 , n71034 , n71035 , n71036 , n71037 , n71038 , n71039 , n71040 , n71041 , n71042 ,
     n71043 , n71044 , n71045 , n71046 , n71047 , n71048 , n71049 , n71050 , n71051 , n71052 ,
     n71053 , n71054 , n71055 , n71056 , n71057 , n71058 , n71059 , n71060 , n71061 , n71062 ,
     n71063 , n71064 , n71065 , n71066 , n71067 , n71068 , n71069 , n71070 , n71071 , n71072 ,
     n71073 , n71074 , n71075 , n71076 , n71077 , n71078 , n71079 , n71080 , n71081 , n71082 ,
     n71083 , n71084 , n71085 , n71086 , n71087 , n71088 , n71089 , n71090 , n71091 , n71092 ,
     n71093 , n71094 , n71095 , n71096 , n71097 , n71098 , n71099 , n71100 , n71101 , n71102 ,
     n71103 , n71104 , n71105 , n71106 , n71107 , n71108 , n71109 , n71110 , n71111 , n71112 ,
     n71113 , n71114 , n71115 , n71116 , n71117 , n71118 , n71119 , n71120 , n71121 , n71122 ,
     n71123 , n71124 , n71125 , n71126 , n71127 , n71128 , n71129 , n71130 , n71131 , n71132 ,
     n71133 , n71134 , n71135 , n71136 , n71137 , n71138 , n71139 , n71140 , n71141 , n71142 ,
     n71143 , n71144 , n71145 , n71146 , n71147 , n71148 , n71149 , n71150 , n71151 , n71152 ,
     n71153 , n71154 , n71155 , n71156 , n71157 , n71158 , n71159 , n71160 , n71161 , n71162 ,
     n71163 , n71164 , n71165 , n71166 , n71167 , n71168 , n71169 , n71170 , n71171 , n71172 ,
     n71173 , n71174 , n71175 , n71176 , n71177 , n71178 , n71179 , n71180 , n71181 , n71182 ,
     n71183 , n71184 , n71185 , n71186 , n71187 , n71188 , n71189 , n71190 , n71191 , n71192 ,
     n71193 , n71194 , n71195 , n71196 , n71197 , n71198 , n71199 , n71200 , n71201 , n71202 ,
     n71203 , n71204 , n71205 , n71206 , n71207 , n71208 , n71209 , n71210 , n71211 , n71212 ,
     n71213 , n71214 , n71215 , n71216 , n71217 , n71218 , n71219 , n71220 , n71221 , n71222 ,
     n71223 , n71224 , n71225 , n71226 , n71227 , n71228 , n71229 , n71230 , n71231 , n71232 ,
     n71233 , n71234 , n71235 , n71236 , n71237 , n71238 , n71239 , n71240 , n71241 , n71242 ,
     n71243 , n71244 , n71245 , n71246 , n71247 , n71248 , n71249 , n71250 , n71251 , n71252 ,
     n71253 , n71254 , n71255 , n71256 , n71257 , n71258 , n71259 , n71260 , n71261 , n71262 ,
     n71263 , n71264 , n71265 , n71266 , n71267 , n71268 , n71269 , n71270 , n71271 , n71272 ,
     n71273 , n71274 , n71275 , n71276 , n71277 , n71278 , n71279 , n71280 , n71281 , n71282 ,
     n71283 , n71284 , n71285 , n71286 , n71287 , n71288 , n71289 , n71290 , n71291 , n71292 ,
     n71293 , n71294 , n71295 , n71296 , n71297 , n71298 , n71299 , n71300 , n71301 , n71302 ,
     n71303 , n71304 , n71305 , n71306 , n71307 , n71308 , n71309 , n71310 , n71311 , n71312 ,
     n71313 , n71314 , n71315 , n71316 , n71317 , n71318 , n71319 , n71320 , n71321 , n71322 ,
     n71323 , n71324 , n71325 , n71326 , n71327 , n71328 , n71329 , n71330 , n71331 , n71332 ,
     n71333 , n71334 , n71335 , n71336 , n71337 , n71338 , n71339 , n71340 , n71341 , n71342 ,
     n71343 , n71344 , n71345 , n71346 , n71347 , n71348 , n71349 , n71350 , n71351 , n71352 ,
     n71353 , n71354 , n71355 , n71356 , n71357 , n71358 , n71359 , n71360 , n71361 , n71362 ,
     n71363 , n71364 , n71365 , n71366 , n71367 , n71368 , n71369 , n71370 , n71371 , n71372 ,
     n71373 , n71374 , n71375 , n71376 , n71377 , n71378 , n71379 , n71380 , n71381 , n71382 ,
     n71383 , n71384 , n71385 , n71386 , n71387 , n71388 , n71389 , n71390 , n71391 , n71392 ,
     n71393 , n71394 , n71395 , n71396 , n71397 , n71398 , n71399 , n71400 , n71401 , n71402 ,
     n71403 , n71404 , n71405 , n71406 , n71407 , n71408 , n71409 , n71410 , n71411 , n71412 ,
     n71413 , n71414 , n71415 , n71416 , n71417 , n71418 , n71419 , n71420 , n71421 , n71422 ,
     n71423 , n71424 , n71425 , n71426 , n71427 , n71428 , n71429 , n71430 , n71431 , n71432 ,
     n71433 , n71434 , n71435 , n71436 , n71437 , n71438 , n71439 , n71440 , n71441 , n71442 ,
     n71443 , n71444 , n71445 , n71446 , n71447 , n71448 , n71449 , n71450 , n71451 , n71452 ,
     n71453 , n71454 , n71455 , n71456 , n71457 , n71458 , n71459 , n71460 , n71461 , n71462 ,
     n71463 , n71464 , n71465 , n71466 , n71467 , n71468 , n71469 , n71470 , n71471 , n71472 ,
     n71473 , n71474 , n71475 , n71476 , n71477 , n71478 , n71479 , n71480 , n71481 , n71482 ,
     n71483 , n71484 , n71485 , n71486 , n71487 , n71488 , n71489 , n71490 , n71491 , n71492 ,
     n71493 , n71494 , n71495 , n71496 , n71497 , n71498 , n71499 , n71500 , n71501 , n71502 ,
     n71503 , n71504 , n71505 , n71506 , n71507 , n71508 , n71509 , n71510 , n71511 , n71512 ,
     n71513 , n71514 , n71515 , n71516 , n71517 , n71518 , n71519 , n71520 , n71521 , n71522 ,
     n71523 , n71524 , n71525 , n71526 , n71527 , n71528 , n71529 , n71530 , n71531 , n71532 ,
     n71533 , n71534 , n71535 , n71536 , n71537 , n71538 , n71539 , n71540 , n71541 , n71542 ,
     n71543 , n71544 , n71545 , n71546 , n71547 , n71548 , n71549 , n71550 , n71551 , n71552 ,
     n71553 , n71554 , n71555 , n71556 , n71557 , n71558 , n71559 , n71560 , n71561 , n71562 ,
     n71563 , n71564 , n71565 , n71566 , n71567 , n71568 , n71569 , n71570 , n71571 , n71572 ,
     n71573 , n71574 , n71575 , n71576 , n71577 , n71578 , n71579 , n71580 , n71581 , n71582 ,
     n71583 , n71584 , n71585 , n71586 , n71587 , n71588 , n71589 , n71590 , n71591 , n71592 ,
     n71593 , n71594 , n71595 , n71596 , n71597 , n71598 , n71599 , n71600 , n71601 , n71602 ,
     n71603 , n71604 , n71605 , n71606 , n71607 , n71608 , n71609 , n71610 , n71611 , n71612 ,
     n71613 , n71614 , n71615 , n71616 , n71617 , n71618 , n71619 , n71620 , n71621 , n71622 ,
     n71623 , n71624 , n71625 , n71626 , n71627 , n71628 , n71629 , n71630 , n71631 , n71632 ,
     n71633 , n71634 , n71635 , n71636 , n71637 , n71638 , n71639 , n71640 , n71641 , n71642 ,
     n71643 , n71644 , n71645 , n71646 , n71647 , n71648 , n71649 , n71650 , n71651 , n71652 ,
     n71653 , n71654 , n71655 , n71656 , n71657 , n71658 , n71659 , n71660 , n71661 , n71662 ,
     n71663 , n71664 , n71665 , n71666 , n71667 , n71668 , n71669 , n71670 , n71671 , n71672 ,
     n71673 , n71674 , n71675 , n71676 , n71677 , n71678 , n71679 , n71680 , n71681 , n71682 ,
     n71683 , n71684 , n71685 , n71686 , n71687 , n71688 , n71689 , n71690 , n71691 , n71692 ,
     n71693 , n71694 , n71695 , n71696 , n71697 , n71698 , n71699 , n71700 , n71701 , n71702 ,
     n71703 , n71704 , n71705 , n71706 , n71707 , n71708 , n71709 , n71710 , n71711 , n71712 ,
     n71713 , n71714 , n71715 , n71716 , n71717 , n71718 , n71719 , n71720 , n71721 , n71722 ,
     n71723 , n71724 , n71725 , n71726 , n71727 , n71728 , n71729 , n71730 , n71731 , n71732 ,
     n71733 , n71734 , n71735 , n71736 , n71737 , n71738 , n71739 , n71740 , n71741 , n71742 ,
     n71743 , n71744 , n71745 , n71746 , n71747 , n71748 , n71749 , n71750 , n71751 , n71752 ,
     n71753 , n71754 , n71755 , n71756 , n71757 , n71758 , n71759 , n71760 , n71761 , n71762 ,
     n71763 , n71764 , n71765 , n71766 , n71767 , n71768 , n71769 , n71770 , n71771 , n71772 ,
     n71773 , n71774 , n71775 , n71776 , n71777 , n71778 , n71779 , n71780 , n71781 , n71782 ,
     n71783 , n71784 , n71785 , n71786 , n71787 , n71788 , n71789 , n71790 , n71791 , n71792 ,
     n71793 , n71794 , n71795 , n71796 , n71797 , n71798 , n71799 , n71800 , n71801 , n71802 ,
     n71803 , n71804 , n71805 , n71806 , n71807 , n71808 , n71809 , n71810 , n71811 , n71812 ,
     n71813 , n71814 , n71815 , n71816 , n71817 , n71818 , n71819 , n71820 , n71821 , n71822 ,
     n71823 , n71824 , n71825 , n71826 , n71827 , n71828 , n71829 , n71830 , n71831 , n71832 ,
     n71833 , n71834 , n71835 , n71836 , n71837 , n71838 , n71839 , n71840 , n71841 , n71842 ,
     n71843 , n71844 , n71845 , n71846 , n71847 , n71848 , n71849 , n71850 , n71851 , n71852 ,
     n71853 , n71854 , n71855 , n71856 , n71857 , n71858 , n71859 , n71860 , n71861 , n71862 ,
     n71863 , n71864 , n71865 , n71866 , n71867 , n71868 , n71869 , n71870 , n71871 , n71872 ,
     n71873 , n71874 , n71875 , n71876 , n71877 , n71878 , n71879 , n71880 , n71881 , n71882 ,
     n71883 , n71884 , n71885 , n71886 , n71887 , n71888 , n71889 , n71890 , n71891 , n71892 ,
     n71893 , n71894 , n71895 , n71896 , n71897 , n71898 , n71899 , n71900 , n71901 , n71902 ,
     n71903 , n71904 , n71905 , n71906 , n71907 , n71908 , n71909 , n71910 , n71911 , n71912 ,
     n71913 , n71914 , n71915 , n71916 , n71917 , n71918 , n71919 , n71920 , n71921 , n71922 ,
     n71923 , n71924 , n71925 , n71926 , n71927 , n71928 , n71929 , n71930 , n71931 , n71932 ,
     n71933 , n71934 , n71935 , n71936 , n71937 , n71938 , n71939 , n71940 , n71941 , n71942 ,
     n71943 , n71944 , n71945 , n71946 , n71947 , n71948 , n71949 , n71950 , n71951 , n71952 ,
     n71953 , n71954 , n71955 , n71956 , n71957 , n71958 , n71959 , n71960 , n71961 , n71962 ,
     n71963 , n71964 , n71965 , n71966 , n71967 , n71968 , n71969 , n71970 , n71971 , n71972 ,
     n71973 , n71974 , n71975 , n71976 , n71977 , n71978 , n71979 , n71980 , n71981 , n71982 ,
     n71983 , n71984 , n71985 , n71986 , n71987 , n71988 , n71989 , n71990 , n71991 , n71992 ,
     n71993 , n71994 , n71995 , n71996 , n71997 , n71998 , n71999 , n72000 , n72001 , n72002 ,
     n72003 , n72004 , n72005 , n72006 , n72007 , n72008 , n72009 , n72010 , n72011 , n72012 ,
     n72013 , n72014 , n72015 , n72016 , n72017 , n72018 , n72019 , n72020 , n72021 , n72022 ,
     n72023 , n72024 , n72025 , n72026 , n72027 , n72028 , n72029 , n72030 , n72031 , n72032 ,
     n72033 , n72034 , n72035 , n72036 , n72037 , n72038 , n72039 , n72040 , n72041 , n72042 ,
     n72043 , n72044 , n72045 , n72046 , n72047 , n72048 , n72049 , n72050 , n72051 , n72052 ,
     n72053 , n72054 , n72055 , n72056 , n72057 , n72058 , n72059 , n72060 , n72061 , n72062 ,
     n72063 , n72064 , n72065 , n72066 , n72067 , n72068 , n72069 , n72070 , n72071 , n72072 ,
     n72073 , n72074 , n72075 , n72076 , n72077 , n72078 , n72079 , n72080 , n72081 , n72082 ,
     n72083 , n72084 , n72085 , n72086 , n72087 , n72088 , n72089 , n72090 , n72091 , n72092 ,
     n72093 , n72094 , n72095 , n72096 , n72097 , n72098 , n72099 , n72100 , n72101 , n72102 ,
     n72103 , n72104 , n72105 , n72106 , n72107 , n72108 , n72109 , n72110 , n72111 , n72112 ,
     n72113 , n72114 , n72115 , n72116 , n72117 , n72118 , n72119 , n72120 , n72121 , n72122 ,
     n72123 , n72124 , n72125 , n72126 , n72127 , n72128 , n72129 , n72130 , n72131 , n72132 ,
     n72133 , n72134 , n72135 , n72136 , n72137 , n72138 , n72139 , n72140 , n72141 , n72142 ,
     n72143 , n72144 , n72145 , n72146 , n72147 , n72148 , n72149 , n72150 , n72151 , n72152 ,
     n72153 , n72154 , n72155 , n72156 , n72157 , n72158 , n72159 , n72160 , n72161 , n72162 ,
     n72163 , n72164 , n72165 , n72166 , n72167 , n72168 , n72169 , n72170 , n72171 , n72172 ,
     n72173 , n72174 , n72175 , n72176 , n72177 , n72178 , n72179 , n72180 , n72181 , n72182 ,
     n72183 , n72184 , n72185 , n72186 , n72187 , n72188 , n72189 , n72190 , n72191 , n72192 ,
     n72193 , n72194 , n72195 , n72196 , n72197 , n72198 , n72199 , n72200 , n72201 , n72202 ,
     n72203 , n72204 , n72205 , n72206 , n72207 , n72208 , n72209 , n72210 , n72211 , n72212 ,
     n72213 , n72214 , n72215 , n72216 , n72217 , n72218 , n72219 , n72220 , n72221 , n72222 ,
     n72223 , n72224 , n72225 , n72226 , n72227 , n72228 , n72229 , n72230 , n72231 , n72232 ,
     n72233 , n72234 , n72235 , n72236 , n72237 , n72238 , n72239 , n72240 , n72241 , n72242 ,
     n72243 , n72244 , n72245 , n72246 , n72247 , n72248 , n72249 , n72250 , n72251 , n72252 ,
     n72253 , n72254 , n72255 , n72256 , n72257 , n72258 , n72259 , n72260 , n72261 , n72262 ,
     n72263 , n72264 , n72265 , n72266 , n72267 , n72268 , n72269 , n72270 , n72271 , n72272 ,
     n72273 , n72274 , n72275 , n72276 , n72277 , n72278 , n72279 , n72280 , n72281 , n72282 ,
     n72283 , n72284 , n72285 , n72286 , n72287 , n72288 , n72289 , n72290 , n72291 , n72292 ,
     n72293 , n72294 , n72295 , n72296 , n72297 , n72298 , n72299 , n72300 , n72301 , n72302 ,
     n72303 , n72304 , n72305 , n72306 , n72307 , n72308 , n72309 , n72310 , n72311 , n72312 ,
     n72313 , n72314 , n72315 , n72316 , n72317 , n72318 , n72319 , n72320 , n72321 , n72322 ,
     n72323 , n72324 , n72325 , n72326 , n72327 , n72328 , n72329 , n72330 , n72331 , n72332 ,
     n72333 , n72334 , n72335 , n72336 , n72337 , n72338 , n72339 , n72340 , n72341 , n72342 ,
     n72343 , n72344 , n72345 , n72346 , n72347 , n72348 , n72349 , n72350 , n72351 , n72352 ,
     n72353 , n72354 , n72355 , n72356 , n72357 , n72358 , n72359 , n72360 , n72361 , n72362 ,
     n72363 , n72364 , n72365 , n72366 , n72367 , n72368 , n72369 , n72370 , n72371 , n72372 ,
     n72373 , n72374 , n72375 , n72376 , n72377 , n72378 , n72379 , n72380 , n72381 , n72382 ,
     n72383 , n72384 , n72385 , n72386 , n72387 , n72388 , n72389 , n72390 , n72391 , n72392 ,
     n72393 , n72394 , n72395 , n72396 , n72397 , n72398 , n72399 , n72400 , n72401 , n72402 ,
     n72403 , n72404 , n72405 , n72406 , n72407 , n72408 , n72409 , n72410 , n72411 , n72412 ,
     n72413 , n72414 , n72415 , n72416 , n72417 , n72418 , n72419 , n72420 , n72421 , n72422 ,
     n72423 , n72424 , n72425 , n72426 , n72427 , n72428 , n72429 , n72430 , n72431 , n72432 ,
     n72433 , n72434 , n72435 , n72436 , n72437 , n72438 , n72439 , n72440 , n72441 , n72442 ,
     n72443 , n72444 , n72445 , n72446 , n72447 , n72448 , n72449 , n72450 , n72451 , n72452 ,
     n72453 , n72454 , n72455 , n72456 , n72457 , n72458 , n72459 , n72460 , n72461 , n72462 ,
     n72463 , n72464 , n72465 , n72466 , n72467 , n72468 , n72469 , n72470 , n72471 , n72472 ,
     n72473 , n72474 , n72475 , n72476 , n72477 , n72478 , n72479 , n72480 , n72481 , n72482 ,
     n72483 , n72484 , n72485 , n72486 , n72487 , n72488 , n72489 , n72490 , n72491 , n72492 ,
     n72493 , n72494 , n72495 , n72496 , n72497 , n72498 , n72499 , n72500 , n72501 , n72502 ,
     n72503 , n72504 , n72505 , n72506 , n72507 , n72508 , n72509 , n72510 , n72511 , n72512 ,
     n72513 , n72514 , n72515 , n72516 , n72517 , n72518 , n72519 , n72520 , n72521 , n72522 ,
     n72523 , n72524 , n72525 , n72526 , n72527 , n72528 , n72529 , n72530 , n72531 , n72532 ,
     n72533 , n72534 , n72535 , n72536 , n72537 , n72538 , n72539 , n72540 , n72541 , n72542 ,
     n72543 , n72544 , n72545 , n72546 , n72547 , n72548 , n72549 , n72550 , n72551 , n72552 ,
     n72553 , n72554 , n72555 , n72556 , n72557 , n72558 , n72559 , n72560 , n72561 , n72562 ,
     n72563 , n72564 , n72565 , n72566 , n72567 , n72568 , n72569 , n72570 , n72571 , n72572 ,
     n72573 , n72574 , n72575 , n72576 , n72577 , n72578 , n72579 , n72580 , n72581 , n72582 ,
     n72583 , n72584 , n72585 , n72586 , n72587 , n72588 , n72589 , n72590 , n72591 , n72592 ,
     n72593 , n72594 , n72595 , n72596 , n72597 , n72598 , n72599 , n72600 , n72601 , n72602 ,
     n72603 , n72604 , n72605 , n72606 , n72607 , n72608 , n72609 , n72610 , n72611 , n72612 ,
     n72613 , n72614 , n72615 , n72616 , n72617 , n72618 , n72619 , n72620 , n72621 , n72622 ,
     n72623 , n72624 , n72625 , n72626 , n72627 , n72628 , n72629 , n72630 , n72631 , n72632 ,
     n72633 , n72634 , n72635 , n72636 , n72637 , n72638 , n72639 , n72640 , n72641 , n72642 ,
     n72643 , n72644 , n72645 , n72646 , n72647 , n72648 , n72649 , n72650 , n72651 , n72652 ,
     n72653 , n72654 , n72655 , n72656 , n72657 , n72658 , n72659 , n72660 , n72661 , n72662 ,
     n72663 , n72664 , n72665 , n72666 , n72667 , n72668 , n72669 , n72670 , n72671 , n72672 ,
     n72673 , n72674 , n72675 , n72676 , n72677 , n72678 , n72679 , n72680 , n72681 , n72682 ,
     n72683 , n72684 , n72685 , n72686 , n72687 , n72688 , n72689 , n72690 , n72691 , n72692 ,
     n72693 , n72694 , n72695 , n72696 , n72697 , n72698 , n72699 , n72700 , n72701 , n72702 ,
     n72703 , n72704 , n72705 , n72706 , n72707 , n72708 , n72709 , n72710 , n72711 , n72712 ,
     n72713 , n72714 , n72715 , n72716 , n72717 , n72718 , n72719 , n72720 , n72721 , n72722 ,
     n72723 , n72724 , n72725 , n72726 , n72727 , n72728 , n72729 , n72730 , n72731 , n72732 ,
     n72733 , n72734 , n72735 , n72736 , n72737 , n72738 , n72739 , n72740 , n72741 , n72742 ,
     n72743 , n72744 , n72745 , n72746 , n72747 , n72748 , n72749 , n72750 , n72751 , n72752 ,
     n72753 , n72754 , n72755 , n72756 , n72757 , n72758 , n72759 , n72760 , n72761 , n72762 ,
     n72763 , n72764 , n72765 , n72766 , n72767 , n72768 , n72769 , n72770 , n72771 , n72772 ,
     n72773 , n72774 , n72775 , n72776 , n72777 , n72778 , n72779 , n72780 , n72781 , n72782 ,
     n72783 , n72784 , n72785 , n72786 , n72787 , n72788 , n72789 , n72790 , n72791 , n72792 ,
     n72793 , n72794 , n72795 , n72796 , n72797 , n72798 , n72799 , n72800 , n72801 , n72802 ,
     n72803 , n72804 , n72805 , n72806 , n72807 , n72808 , n72809 , n72810 , n72811 , n72812 ,
     n72813 , n72814 , n72815 , n72816 , n72817 , n72818 , n72819 , n72820 , n72821 , n72822 ,
     n72823 , n72824 , n72825 , n72826 , n72827 , n72828 , n72829 , n72830 , n72831 , n72832 ,
     n72833 , n72834 , n72835 , n72836 , n72837 , n72838 , n72839 , n72840 , n72841 , n72842 ,
     n72843 , n72844 , n72845 , n72846 , n72847 , n72848 , n72849 , n72850 , n72851 , n72852 ,
     n72853 , n72854 , n72855 , n72856 , n72857 , n72858 , n72859 , n72860 , n72861 , n72862 ,
     n72863 , n72864 , n72865 , n72866 , n72867 , n72868 , n72869 , n72870 , n72871 , n72872 ,
     n72873 , n72874 , n72875 , n72876 , n72877 , n72878 , n72879 , n72880 , n72881 , n72882 ,
     n72883 , n72884 , n72885 , n72886 , n72887 , n72888 , n72889 , n72890 , n72891 , n72892 ,
     n72893 , n72894 , n72895 , n72896 , n72897 , n72898 , n72899 , n72900 , n72901 , n72902 ,
     n72903 , n72904 , n72905 , n72906 , n72907 , n72908 , n72909 , n72910 , n72911 , n72912 ,
     n72913 , n72914 , n72915 , n72916 , n72917 , n72918 , n72919 , n72920 , n72921 , n72922 ,
     n72923 , n72924 , n72925 , n72926 , n72927 , n72928 , n72929 , n72930 , n72931 , n72932 ,
     n72933 , n72934 , n72935 , n72936 , n72937 , n72938 , n72939 , n72940 , n72941 , n72942 ,
     n72943 , n72944 , n72945 , n72946 , n72947 , n72948 , n72949 , n72950 , n72951 , n72952 ,
     n72953 , n72954 , n72955 , n72956 , n72957 , n72958 , n72959 , n72960 , n72961 , n72962 ,
     n72963 , n72964 , n72965 , n72966 , n72967 , n72968 , n72969 , n72970 , n72971 , n72972 ,
     n72973 , n72974 , n72975 , n72976 , n72977 , n72978 , n72979 , n72980 , n72981 , n72982 ,
     n72983 , n72984 , n72985 , n72986 , n72987 , n72988 , n72989 , n72990 , n72991 , n72992 ,
     n72993 , n72994 , n72995 , n72996 , n72997 , n72998 , n72999 , n73000 , n73001 , n73002 ,
     n73003 , n73004 , n73005 , n73006 , n73007 , n73008 , n73009 , n73010 , n73011 , n73012 ,
     n73013 , n73014 , n73015 , n73016 , n73017 , n73018 , n73019 , n73020 , n73021 , n73022 ,
     n73023 , n73024 , n73025 , n73026 , n73027 , n73028 , n73029 , n73030 , n73031 , n73032 ,
     n73033 , n73034 , n73035 , n73036 , n73037 , n73038 , n73039 , n73040 , n73041 , n73042 ,
     n73043 , n73044 , n73045 , n73046 , n73047 , n73048 , n73049 , n73050 , n73051 , n73052 ,
     n73053 , n73054 , n73055 , n73056 , n73057 , n73058 , n73059 , n73060 , n73061 , n73062 ,
     n73063 , n73064 , n73065 , n73066 , n73067 , n73068 , n73069 , n73070 , n73071 , n73072 ,
     n73073 , n73074 , n73075 , n73076 , n73077 , n73078 , n73079 , n73080 , n73081 , n73082 ,
     n73083 , n73084 , n73085 , n73086 , n73087 , n73088 , n73089 , n73090 , n73091 , n73092 ,
     n73093 , n73094 , n73095 , n73096 , n73097 , n73098 , n73099 , n73100 , n73101 , n73102 ,
     n73103 , n73104 , n73105 , n73106 , n73107 , n73108 , n73109 , n73110 , n73111 , n73112 ,
     n73113 , n73114 , n73115 , n73116 , n73117 , n73118 , n73119 , n73120 , n73121 , n73122 ,
     n73123 , n73124 , n73125 , n73126 , n73127 , n73128 , n73129 , n73130 , n73131 , n73132 ,
     n73133 , n73134 , n73135 , n73136 , n73137 , n73138 , n73139 , n73140 , n73141 , n73142 ,
     n73143 , n73144 , n73145 , n73146 , n73147 , n73148 , n73149 , n73150 , n73151 , n73152 ,
     n73153 , n73154 , n73155 , n73156 , n73157 , n73158 , n73159 , n73160 , n73161 , n73162 ,
     n73163 , n73164 , n73165 , n73166 , n73167 , n73168 , n73169 , n73170 , n73171 , n73172 ,
     n73173 , n73174 , n73175 , n73176 , n73177 , n73178 , n73179 , n73180 , n73181 , n73182 ,
     n73183 , n73184 , n73185 , n73186 , n73187 , n73188 , n73189 , n73190 , n73191 , n73192 ,
     n73193 , n73194 , n73195 , n73196 , n73197 , n73198 , n73199 , n73200 , n73201 , n73202 ,
     n73203 , n73204 , n73205 , n73206 , n73207 , n73208 , n73209 , n73210 , n73211 , n73212 ,
     n73213 , n73214 , n73215 , n73216 , n73217 , n73218 , n73219 , n73220 , n73221 , n73222 ,
     n73223 , n73224 , n73225 , n73226 , n73227 , n73228 , n73229 , n73230 , n73231 , n73232 ,
     n73233 , n73234 , n73235 , n73236 , n73237 , n73238 , n73239 , n73240 , n73241 , n73242 ,
     n73243 , n73244 , n73245 , n73246 , n73247 , n73248 , n73249 , n73250 , n73251 , n73252 ,
     n73253 , n73254 , n73255 , n73256 , n73257 , n73258 , n73259 , n73260 , n73261 , n73262 ,
     n73263 , n73264 , n73265 , n73266 , n73267 , n73268 , n73269 , n73270 , n73271 , n73272 ,
     n73273 , n73274 , n73275 , n73276 , n73277 , n73278 , n73279 , n73280 , n73281 , n73282 ,
     n73283 , n73284 , n73285 , n73286 , n73287 , n73288 , n73289 , n73290 , n73291 , n73292 ,
     n73293 , n73294 , n73295 , n73296 , n73297 , n73298 , n73299 , n73300 , n73301 , n73302 ,
     n73303 , n73304 , n73305 , n73306 , n73307 , n73308 , n73309 , n73310 , n73311 , n73312 ,
     n73313 , n73314 , n73315 , n73316 , n73317 , n73318 , n73319 , n73320 , n73321 , n73322 ,
     n73323 , n73324 , n73325 , n73326 , n73327 , n73328 , n73329 , n73330 , n73331 , n73332 ,
     n73333 , n73334 , n73335 , n73336 , n73337 , n73338 , n73339 , n73340 , n73341 , n73342 ,
     n73343 , n73344 , n73345 , n73346 , n73347 , n73348 , n73349 , n73350 , n73351 , n73352 ,
     n73353 , n73354 , n73355 , n73356 , n73357 , n73358 , n73359 , n73360 , n73361 , n73362 ,
     n73363 , n73364 , n73365 , n73366 , n73367 , n73368 , n73369 , n73370 , n73371 , n73372 ,
     n73373 , n73374 , n73375 , n73376 , n73377 , n73378 , n73379 , n73380 , n73381 , n73382 ,
     n73383 , n73384 , n73385 , n73386 , n73387 , n73388 , n73389 , n73390 , n73391 , n73392 ,
     n73393 , n73394 , n73395 , n73396 , n73397 , n73398 , n73399 , n73400 , n73401 , n73402 ,
     n73403 , n73404 , n73405 , n73406 , n73407 , n73408 , n73409 , n73410 , n73411 , n73412 ,
     n73413 , n73414 , n73415 , n73416 , n73417 , n73418 , n73419 , n73420 , n73421 , n73422 ,
     n73423 , n73424 , n73425 , n73426 , n73427 , n73428 , n73429 , n73430 , n73431 , n73432 ,
     n73433 , n73434 , n73435 , n73436 , n73437 , n73438 , n73439 , n73440 , n73441 , n73442 ,
     n73443 , n73444 , n73445 , n73446 , n73447 , n73448 , n73449 , n73450 , n73451 , n73452 ,
     n73453 , n73454 , n73455 , n73456 , n73457 , n73458 , n73459 , n73460 , n73461 , n73462 ,
     n73463 , n73464 , n73465 , n73466 , n73467 , n73468 , n73469 , n73470 , n73471 , n73472 ,
     n73473 , n73474 , n73475 , n73476 , n73477 , n73478 , n73479 , n73480 , n73481 , n73482 ,
     n73483 , n73484 , n73485 , n73486 , n73487 , n73488 , n73489 , n73490 , n73491 , n73492 ,
     n73493 , n73494 , n73495 , n73496 , n73497 , n73498 , n73499 , n73500 , n73501 , n73502 ,
     n73503 , n73504 , n73505 , n73506 , n73507 , n73508 , n73509 , n73510 , n73511 , n73512 ,
     n73513 , n73514 , n73515 , n73516 , n73517 , n73518 , n73519 , n73520 , n73521 , n73522 ,
     n73523 , n73524 , n73525 , n73526 , n73527 , n73528 , n73529 , n73530 , n73531 , n73532 ,
     n73533 , n73534 , n73535 , n73536 , n73537 , n73538 , n73539 , n73540 , n73541 , n73542 ,
     n73543 , n73544 , n73545 , n73546 , n73547 , n73548 , n73549 , n73550 , n73551 , n73552 ,
     n73553 , n73554 , n73555 , n73556 , n73557 , n73558 , n73559 , n73560 , n73561 , n73562 ,
     n73563 , n73564 , n73565 , n73566 , n73567 , n73568 , n73569 , n73570 , n73571 , n73572 ,
     n73573 , n73574 , n73575 , n73576 , n73577 , n73578 , n73579 , n73580 , n73581 , n73582 ,
     n73583 , n73584 , n73585 , n73586 , n73587 , n73588 , n73589 , n73590 , n73591 , n73592 ,
     n73593 , n73594 , n73595 , n73596 , n73597 , n73598 , n73599 , n73600 , n73601 , n73602 ,
     n73603 , n73604 , n73605 , n73606 , n73607 , n73608 , n73609 , n73610 , n73611 , n73612 ,
     n73613 , n73614 , n73615 , n73616 , n73617 , n73618 , n73619 , n73620 , n73621 , n73622 ,
     n73623 , n73624 , n73625 , n73626 , n73627 , n73628 , n73629 , n73630 , n73631 , n73632 ,
     n73633 , n73634 , n73635 , n73636 , n73637 , n73638 , n73639 , n73640 , n73641 , n73642 ,
     n73643 , n73644 , n73645 , n73646 , n73647 , n73648 , n73649 , n73650 , n73651 , n73652 ,
     n73653 , n73654 , n73655 , n73656 , n73657 , n73658 , n73659 , n73660 , n73661 , n73662 ,
     n73663 , n73664 , n73665 , n73666 , n73667 , n73668 , n73669 , n73670 , n73671 , n73672 ,
     n73673 , n73674 , n73675 , n73676 , n73677 , n73678 , n73679 , n73680 , n73681 , n73682 ,
     n73683 , n73684 , n73685 , n73686 , n73687 , n73688 , n73689 , n73690 , n73691 , n73692 ,
     n73693 , n73694 , n73695 , n73696 , n73697 , n73698 , n73699 , n73700 , n73701 , n73702 ,
     n73703 , n73704 , n73705 , n73706 , n73707 , n73708 , n73709 , n73710 , n73711 , n73712 ,
     n73713 , n73714 , n73715 , n73716 , n73717 , n73718 , n73719 , n73720 , n73721 , n73722 ,
     n73723 , n73724 , n73725 , n73726 , n73727 , n73728 , n73729 , n73730 , n73731 , n73732 ,
     n73733 , n73734 , n73735 , n73736 , n73737 , n73738 , n73739 , n73740 , n73741 , n73742 ,
     n73743 , n73744 , n73745 , n73746 , n73747 , n73748 , n73749 , n73750 , n73751 , n73752 ,
     n73753 , n73754 , n73755 , n73756 , n73757 , n73758 , n73759 , n73760 , n73761 , n73762 ,
     n73763 , n73764 , n73765 , n73766 , n73767 , n73768 , n73769 , n73770 , n73771 , n73772 ,
     n73773 , n73774 , n73775 , n73776 , n73777 , n73778 , n73779 , n73780 , n73781 , n73782 ,
     n73783 , n73784 , n73785 , n73786 , n73787 , n73788 , n73789 , n73790 , n73791 , n73792 ,
     n73793 , n73794 , n73795 , n73796 , n73797 , n73798 , n73799 , n73800 , n73801 , n73802 ,
     n73803 , n73804 , n73805 , n73806 , n73807 , n73808 , n73809 , n73810 , n73811 , n73812 ,
     n73813 , n73814 , n73815 , n73816 , n73817 , n73818 , n73819 , n73820 , n73821 , n73822 ,
     n73823 , n73824 , n73825 , n73826 , n73827 , n73828 , n73829 , n73830 , n73831 , n73832 ,
     n73833 , n73834 , n73835 , n73836 , n73837 , n73838 , n73839 , n73840 , n73841 , n73842 ,
     n73843 , n73844 , n73845 , n73846 , n73847 , n73848 , n73849 , n73850 , n73851 , n73852 ,
     n73853 , n73854 , n73855 , n73856 , n73857 , n73858 , n73859 , n73860 , n73861 , n73862 ,
     n73863 , n73864 , n73865 , n73866 , n73867 , n73868 , n73869 , n73870 , n73871 , n73872 ,
     n73873 , n73874 , n73875 , n73876 , n73877 , n73878 , n73879 , n73880 , n73881 , n73882 ,
     n73883 , n73884 , n73885 , n73886 , n73887 , n73888 , n73889 , n73890 , n73891 , n73892 ,
     n73893 , n73894 , n73895 , n73896 , n73897 , n73898 , n73899 , n73900 , n73901 , n73902 ,
     n73903 , n73904 , n73905 , n73906 , n73907 , n73908 , n73909 , n73910 , n73911 , n73912 ,
     n73913 , n73914 , n73915 , n73916 , n73917 , n73918 , n73919 , n73920 , n73921 , n73922 ,
     n73923 , n73924 , n73925 , n73926 , n73927 , n73928 , n73929 , n73930 , n73931 , n73932 ,
     n73933 , n73934 , n73935 , n73936 , n73937 , n73938 , n73939 , n73940 , n73941 , n73942 ,
     n73943 , n73944 , n73945 , n73946 , n73947 , n73948 , n73949 , n73950 , n73951 , n73952 ,
     n73953 , n73954 , n73955 , n73956 , n73957 , n73958 , n73959 , n73960 , n73961 , n73962 ,
     n73963 , n73964 , n73965 , n73966 , n73967 , n73968 , n73969 , n73970 , n73971 , n73972 ,
     n73973 , n73974 , n73975 , n73976 , n73977 , n73978 , n73979 , n73980 , n73981 , n73982 ,
     n73983 , n73984 , n73985 , n73986 , n73987 , n73988 , n73989 , n73990 , n73991 , n73992 ,
     n73993 , n73994 , n73995 , n73996 , n73997 , n73998 , n73999 , n74000 , n74001 , n74002 ,
     n74003 , n74004 , n74005 , n74006 , n74007 , n74008 , n74009 , n74010 , n74011 , n74012 ,
     n74013 , n74014 , n74015 , n74016 , n74017 , n74018 , n74019 , n74020 , n74021 , n74022 ,
     n74023 , n74024 , n74025 , n74026 , n74027 , n74028 , n74029 , n74030 , n74031 , n74032 ,
     n74033 , n74034 , n74035 , n74036 , n74037 , n74038 , n74039 , n74040 , n74041 , n74042 ,
     n74043 , n74044 , n74045 , n74046 , n74047 , n74048 , n74049 , n74050 , n74051 , n74052 ,
     n74053 , n74054 , n74055 , n74056 , n74057 , n74058 , n74059 , n74060 , n74061 , n74062 ,
     n74063 , n74064 , n74065 , n74066 , n74067 , n74068 , n74069 , n74070 , n74071 , n74072 ,
     n74073 , n74074 , n74075 , n74076 , n74077 , n74078 , n74079 , n74080 , n74081 , n74082 ,
     n74083 , n74084 , n74085 , n74086 , n74087 , n74088 , n74089 , n74090 , n74091 , n74092 ,
     n74093 , n74094 , n74095 , n74096 , n74097 , n74098 , n74099 , n74100 , n74101 , n74102 ,
     n74103 , n74104 , n74105 , n74106 , n74107 , n74108 , n74109 , n74110 , n74111 , n74112 ,
     n74113 , n74114 , n74115 , n74116 , n74117 , n74118 , n74119 , n74120 , n74121 , n74122 ,
     n74123 , n74124 , n74125 , n74126 , n74127 , n74128 , n74129 , n74130 , n74131 , n74132 ,
     n74133 , n74134 , n74135 , n74136 , n74137 , n74138 , n74139 , n74140 , n74141 , n74142 ,
     n74143 , n74144 , n74145 , n74146 , n74147 , n74148 , n74149 , n74150 , n74151 , n74152 ,
     n74153 , n74154 , n74155 , n74156 , n74157 , n74158 , n74159 , n74160 , n74161 , n74162 ,
     n74163 , n74164 , n74165 , n74166 , n74167 , n74168 , n74169 , n74170 , n74171 , n74172 ,
     n74173 , n74174 , n74175 , n74176 , n74177 , n74178 , n74179 , n74180 , n74181 , n74182 ,
     n74183 , n74184 , n74185 , n74186 , n74187 , n74188 , n74189 , n74190 , n74191 , n74192 ,
     n74193 , n74194 , n74195 , n74196 , n74197 , n74198 , n74199 , n74200 , n74201 , n74202 ,
     n74203 , n74204 , n74205 , n74206 , n74207 , n74208 , n74209 , n74210 , n74211 , n74212 ,
     n74213 , n74214 , n74215 , n74216 , n74217 , n74218 , n74219 , n74220 , n74221 , n74222 ,
     n74223 , n74224 , n74225 , n74226 , n74227 , n74228 , n74229 , n74230 , n74231 , n74232 ,
     n74233 , n74234 , n74235 , n74236 , n74237 , n74238 , n74239 , n74240 , n74241 , n74242 ,
     n74243 , n74244 , n74245 , n74246 , n74247 , n74248 , n74249 , n74250 , n74251 , n74252 ,
     n74253 , n74254 , n74255 , n74256 , n74257 , n74258 , n74259 , n74260 , n74261 , n74262 ,
     n74263 , n74264 , n74265 , n74266 , n74267 , n74268 , n74269 , n74270 , n74271 , n74272 ,
     n74273 , n74274 , n74275 , n74276 , n74277 , n74278 , n74279 , n74280 , n74281 , n74282 ,
     n74283 , n74284 , n74285 , n74286 , n74287 , n74288 , n74289 , n74290 , n74291 , n74292 ,
     n74293 , n74294 , n74295 , n74296 , n74297 , n74298 , n74299 , n74300 , n74301 , n74302 ,
     n74303 , n74304 , n74305 , n74306 , n74307 , n74308 , n74309 , n74310 , n74311 , n74312 ,
     n74313 , n74314 , n74315 , n74316 , n74317 , n74318 , n74319 , n74320 , n74321 , n74322 ,
     n74323 , n74324 , n74325 , n74326 , n74327 , n74328 , n74329 , n74330 , n74331 , n74332 ,
     n74333 , n74334 , n74335 , n74336 , n74337 , n74338 , n74339 , n74340 , n74341 , n74342 ,
     n74343 , n74344 , n74345 , n74346 , n74347 , n74348 , n74349 , n74350 , n74351 , n74352 ,
     n74353 , n74354 , n74355 , n74356 , n74357 , n74358 , n74359 , n74360 , n74361 , n74362 ,
     n74363 , n74364 , n74365 , n74366 , n74367 , n74368 , n74369 , n74370 , n74371 , n74372 ,
     n74373 , n74374 , n74375 , n74376 , n74377 , n74378 , n74379 , n74380 , n74381 , n74382 ,
     n74383 , n74384 , n74385 , n74386 , n74387 , n74388 , n74389 , n74390 , n74391 , n74392 ,
     n74393 , n74394 , n74395 , n74396 , n74397 , n74398 , n74399 , n74400 , n74401 , n74402 ,
     n74403 , n74404 , n74405 , n74406 , n74407 , n74408 , n74409 , n74410 , n74411 , n74412 ,
     n74413 , n74414 , n74415 , n74416 , n74417 , n74418 , n74419 , n74420 , n74421 , n74422 ,
     n74423 , n74424 , n74425 , n74426 , n74427 , n74428 , n74429 , n74430 , n74431 , n74432 ,
     n74433 , n74434 , n74435 , n74436 , n74437 , n74438 , n74439 , n74440 , n74441 , n74442 ,
     n74443 , n74444 , n74445 , n74446 , n74447 , n74448 , n74449 , n74450 , n74451 , n74452 ,
     n74453 , n74454 , n74455 , n74456 , n74457 , n74458 , n74459 , n74460 , n74461 , n74462 ,
     n74463 , n74464 , n74465 , n74466 , n74467 , n74468 , n74469 , n74470 , n74471 , n74472 ,
     n74473 , n74474 , n74475 , n74476 , n74477 , n74478 , n74479 , n74480 , n74481 , n74482 ,
     n74483 , n74484 , n74485 , n74486 , n74487 , n74488 , n74489 , n74490 , n74491 , n74492 ,
     n74493 , n74494 , n74495 , n74496 , n74497 , n74498 , n74499 , n74500 , n74501 , n74502 ,
     n74503 , n74504 , n74505 , n74506 , n74507 , n74508 , n74509 , n74510 , n74511 , n74512 ,
     n74513 , n74514 , n74515 , n74516 , n74517 , n74518 , n74519 , n74520 , n74521 , n74522 ,
     n74523 , n74524 , n74525 , n74526 , n74527 , n74528 , n74529 , n74530 , n74531 , n74532 ,
     n74533 , n74534 , n74535 , n74536 , n74537 , n74538 , n74539 , n74540 , n74541 , n74542 ,
     n74543 , n74544 , n74545 , n74546 , n74547 , n74548 , n74549 , n74550 , n74551 , n74552 ,
     n74553 , n74554 , n74555 , n74556 , n74557 , n74558 , n74559 , n74560 , n74561 , n74562 ,
     n74563 , n74564 , n74565 , n74566 , n74567 , n74568 , n74569 , n74570 , n74571 , n74572 ,
     n74573 , n74574 , n74575 , n74576 , n74577 , n74578 , n74579 , n74580 , n74581 , n74582 ,
     n74583 , n74584 , n74585 , n74586 , n74587 , n74588 , n74589 , n74590 , n74591 , n74592 ,
     n74593 , n74594 , n74595 , n74596 , n74597 , n74598 , n74599 , n74600 , n74601 , n74602 ,
     n74603 , n74604 , n74605 , n74606 , n74607 , n74608 , n74609 , n74610 , n74611 , n74612 ,
     n74613 , n74614 , n74615 , n74616 , n74617 , n74618 , n74619 , n74620 , n74621 , n74622 ,
     n74623 , n74624 , n74625 , n74626 , n74627 , n74628 , n74629 , n74630 , n74631 , n74632 ,
     n74633 , n74634 , n74635 , n74636 , n74637 , n74638 , n74639 , n74640 , n74641 , n74642 ,
     n74643 , n74644 , n74645 , n74646 , n74647 , n74648 , n74649 , n74650 , n74651 , n74652 ,
     n74653 , n74654 , n74655 , n74656 , n74657 , n74658 , n74659 , n74660 , n74661 , n74662 ,
     n74663 , n74664 , n74665 , n74666 , n74667 , n74668 , n74669 , n74670 , n74671 , n74672 ,
     n74673 , n74674 , n74675 , n74676 , n74677 , n74678 , n74679 , n74680 , n74681 , n74682 ,
     n74683 , n74684 , n74685 , n74686 , n74687 , n74688 , n74689 , n74690 , n74691 , n74692 ,
     n74693 , n74694 , n74695 , n74696 , n74697 , n74698 , n74699 , n74700 , n74701 , n74702 ,
     n74703 , n74704 , n74705 , n74706 , n74707 , n74708 , n74709 , n74710 , n74711 , n74712 ,
     n74713 , n74714 , n74715 , n74716 , n74717 , n74718 , n74719 , n74720 , n74721 , n74722 ,
     n74723 , n74724 , n74725 , n74726 , n74727 , n74728 , n74729 , n74730 , n74731 , n74732 ,
     n74733 , n74734 , n74735 , n74736 , n74737 , n74738 , n74739 , n74740 , n74741 , n74742 ,
     n74743 , n74744 , n74745 , n74746 , n74747 , n74748 , n74749 , n74750 , n74751 , n74752 ,
     n74753 , n74754 , n74755 , n74756 , n74757 , n74758 , n74759 , n74760 , n74761 , n74762 ,
     n74763 , n74764 , n74765 , n74766 , n74767 , n74768 , n74769 , n74770 , n74771 , n74772 ,
     n74773 , n74774 , n74775 , n74776 , n74777 , n74778 , n74779 , n74780 , n74781 , n74782 ,
     n74783 , n74784 , n74785 , n74786 , n74787 , n74788 , n74789 , n74790 , n74791 , n74792 ,
     n74793 , n74794 , n74795 , n74796 , n74797 , n74798 , n74799 , n74800 , n74801 , n74802 ,
     n74803 , n74804 , n74805 , n74806 , n74807 , n74808 , n74809 , n74810 , n74811 , n74812 ,
     n74813 , n74814 , n74815 , n74816 , n74817 , n74818 , n74819 , n74820 , n74821 , n74822 ,
     n74823 , n74824 , n74825 , n74826 , n74827 , n74828 , n74829 , n74830 , n74831 , n74832 ,
     n74833 , n74834 , n74835 , n74836 , n74837 , n74838 , n74839 , n74840 , n74841 , n74842 ,
     n74843 , n74844 , n74845 , n74846 , n74847 , n74848 , n74849 , n74850 , n74851 , n74852 ,
     n74853 , n74854 , n74855 , n74856 , n74857 , n74858 , n74859 , n74860 , n74861 , n74862 ,
     n74863 , n74864 , n74865 , n74866 , n74867 , n74868 , n74869 , n74870 , n74871 , n74872 ,
     n74873 , n74874 , n74875 , n74876 , n74877 , n74878 , n74879 , n74880 , n74881 , n74882 ,
     n74883 , n74884 , n74885 , n74886 , n74887 , n74888 , n74889 , n74890 , n74891 , n74892 ,
     n74893 , n74894 , n74895 , n74896 , n74897 , n74898 , n74899 , n74900 , n74901 , n74902 ,
     n74903 , n74904 , n74905 , n74906 , n74907 , n74908 , n74909 , n74910 , n74911 , n74912 ,
     n74913 , n74914 , n74915 , n74916 , n74917 , n74918 , n74919 , n74920 , n74921 , n74922 ,
     n74923 , n74924 , n74925 , n74926 , n74927 , n74928 , n74929 , n74930 , n74931 , n74932 ,
     n74933 , n74934 , n74935 , n74936 , n74937 , n74938 , n74939 , n74940 , n74941 , n74942 ,
     n74943 , n74944 , n74945 , n74946 , n74947 , n74948 , n74949 , n74950 , n74951 , n74952 ,
     n74953 , n74954 , n74955 , n74956 , n74957 , n74958 , n74959 , n74960 , n74961 , n74962 ,
     n74963 , n74964 , n74965 , n74966 , n74967 , n74968 , n74969 , n74970 , n74971 , n74972 ,
     n74973 , n74974 , n74975 , n74976 , n74977 , n74978 , n74979 , n74980 , n74981 , n74982 ,
     n74983 , n74984 , n74985 , n74986 , n74987 , n74988 , n74989 , n74990 , n74991 , n74992 ,
     n74993 , n74994 , n74995 , n74996 , n74997 , n74998 , n74999 , n75000 , n75001 , n75002 ,
     n75003 , n75004 , n75005 , n75006 , n75007 , n75008 , n75009 , n75010 , n75011 , n75012 ,
     n75013 , n75014 , n75015 , n75016 , n75017 , n75018 , n75019 , n75020 , n75021 , n75022 ,
     n75023 , n75024 , n75025 , n75026 , n75027 , n75028 , n75029 , n75030 , n75031 , n75032 ,
     n75033 , n75034 , n75035 , n75036 , n75037 , n75038 , n75039 , n75040 , n75041 , n75042 ,
     n75043 , n75044 , n75045 , n75046 , n75047 , n75048 , n75049 , n75050 , n75051 , n75052 ,
     n75053 , n75054 , n75055 , n75056 , n75057 , n75058 , n75059 , n75060 , n75061 , n75062 ,
     n75063 , n75064 , n75065 , n75066 , n75067 , n75068 , n75069 , n75070 , n75071 , n75072 ,
     n75073 , n75074 , n75075 , n75076 , n75077 , n75078 , n75079 , n75080 , n75081 , n75082 ,
     n75083 , n75084 , n75085 , n75086 , n75087 , n75088 , n75089 , n75090 , n75091 , n75092 ,
     n75093 , n75094 , n75095 , n75096 , n75097 , n75098 , n75099 , n75100 , n75101 , n75102 ,
     n75103 , n75104 , n75105 , n75106 , n75107 , n75108 , n75109 , n75110 , n75111 , n75112 ,
     n75113 , n75114 , n75115 , n75116 , n75117 , n75118 , n75119 , n75120 , n75121 , n75122 ,
     n75123 , n75124 , n75125 , n75126 , n75127 , n75128 , n75129 , n75130 , n75131 , n75132 ,
     n75133 , n75134 , n75135 , n75136 , n75137 , n75138 , n75139 , n75140 , n75141 , n75142 ,
     n75143 , n75144 , n75145 , n75146 , n75147 , n75148 , n75149 , n75150 , n75151 , n75152 ,
     n75153 , n75154 , n75155 , n75156 , n75157 , n75158 , n75159 , n75160 , n75161 , n75162 ,
     n75163 , n75164 , n75165 , n75166 , n75167 , n75168 , n75169 , n75170 , n75171 , n75172 ,
     n75173 , n75174 , n75175 , n75176 , n75177 , n75178 , n75179 , n75180 , n75181 , n75182 ,
     n75183 , n75184 , n75185 , n75186 , n75187 , n75188 , n75189 , n75190 , n75191 , n75192 ,
     n75193 , n75194 , n75195 , n75196 , n75197 , n75198 , n75199 , n75200 , n75201 , n75202 ,
     n75203 , n75204 , n75205 , n75206 , n75207 , n75208 , n75209 , n75210 , n75211 , n75212 ,
     n75213 , n75214 , n75215 , n75216 , n75217 , n75218 , n75219 , n75220 , n75221 , n75222 ,
     n75223 , n75224 , n75225 , n75226 , n75227 , n75228 , n75229 , n75230 , n75231 , n75232 ,
     n75233 , n75234 , n75235 , n75236 , n75237 , n75238 , n75239 , n75240 , n75241 , n75242 ,
     n75243 , n75244 , n75245 , n75246 , n75247 , n75248 , n75249 , n75250 , n75251 , n75252 ,
     n75253 , n75254 , n75255 , n75256 , n75257 , n75258 , n75259 , n75260 , n75261 , n75262 ,
     n75263 , n75264 , n75265 , n75266 , n75267 , n75268 , n75269 , n75270 , n75271 , n75272 ,
     n75273 , n75274 , n75275 , n75276 , n75277 , n75278 , n75279 , n75280 , n75281 , n75282 ,
     n75283 , n75284 , n75285 , n75286 , n75287 , n75288 , n75289 , n75290 , n75291 , n75292 ,
     n75293 , n75294 , n75295 , n75296 , n75297 , n75298 , n75299 , n75300 , n75301 , n75302 ,
     n75303 , n75304 , n75305 , n75306 , n75307 , n75308 , n75309 , n75310 , n75311 , n75312 ,
     n75313 , n75314 , n75315 , n75316 , n75317 , n75318 , n75319 , n75320 , n75321 , n75322 ,
     n75323 , n75324 , n75325 , n75326 , n75327 , n75328 , n75329 , n75330 , n75331 , n75332 ,
     n75333 , n75334 , n75335 , n75336 , n75337 , n75338 , n75339 , n75340 , n75341 , n75342 ,
     n75343 , n75344 , n75345 , n75346 , n75347 , n75348 , n75349 , n75350 , n75351 , n75352 ,
     n75353 , n75354 , n75355 , n75356 , n75357 , n75358 , n75359 , n75360 , n75361 , n75362 ,
     n75363 , n75364 , n75365 , n75366 , n75367 , n75368 , n75369 , n75370 , n75371 , n75372 ,
     n75373 , n75374 , n75375 , n75376 , n75377 , n75378 , n75379 , n75380 , n75381 , n75382 ,
     n75383 , n75384 , n75385 , n75386 , n75387 , n75388 , n75389 , n75390 , n75391 , n75392 ,
     n75393 , n75394 , n75395 , n75396 , n75397 , n75398 , n75399 , n75400 , n75401 , n75402 ,
     n75403 , n75404 , n75405 , n75406 , n75407 , n75408 , n75409 , n75410 , n75411 , n75412 ,
     n75413 , n75414 , n75415 , n75416 , n75417 , n75418 , n75419 , n75420 , n75421 , n75422 ,
     n75423 , n75424 , n75425 , n75426 , n75427 , n75428 , n75429 , n75430 , n75431 , n75432 ,
     n75433 , n75434 , n75435 , n75436 , n75437 , n75438 , n75439 , n75440 , n75441 , n75442 ,
     n75443 , n75444 , n75445 , n75446 , n75447 , n75448 , n75449 , n75450 , n75451 , n75452 ,
     n75453 , n75454 , n75455 , n75456 , n75457 , n75458 , n75459 , n75460 , n75461 , n75462 ,
     n75463 , n75464 , n75465 , n75466 , n75467 , n75468 , n75469 , n75470 , n75471 , n75472 ,
     n75473 , n75474 , n75475 , n75476 , n75477 , n75478 , n75479 , n75480 , n75481 , n75482 ,
     n75483 , n75484 , n75485 , n75486 , n75487 , n75488 , n75489 , n75490 , n75491 , n75492 ,
     n75493 , n75494 , n75495 , n75496 , n75497 , n75498 , n75499 , n75500 , n75501 , n75502 ,
     n75503 , n75504 , n75505 , n75506 , n75507 , n75508 , n75509 , n75510 , n75511 , n75512 ,
     n75513 , n75514 , n75515 , n75516 , n75517 , n75518 , n75519 , n75520 , n75521 , n75522 ,
     n75523 , n75524 , n75525 , n75526 , n75527 , n75528 , n75529 , n75530 , n75531 , n75532 ,
     n75533 , n75534 , n75535 , n75536 , n75537 , n75538 , n75539 , n75540 , n75541 , n75542 ,
     n75543 , n75544 , n75545 , n75546 , n75547 , n75548 , n75549 , n75550 , n75551 , n75552 ,
     n75553 , n75554 , n75555 , n75556 , n75557 , n75558 , n75559 , n75560 , n75561 , n75562 ,
     n75563 , n75564 , n75565 , n75566 , n75567 , n75568 , n75569 , n75570 , n75571 , n75572 ,
     n75573 , n75574 , n75575 , n75576 , n75577 , n75578 , n75579 , n75580 , n75581 , n75582 ,
     n75583 , n75584 , n75585 , n75586 , n75587 , n75588 , n75589 , n75590 , n75591 , n75592 ,
     n75593 , n75594 , n75595 , n75596 , n75597 , n75598 , n75599 , n75600 , n75601 , n75602 ,
     n75603 , n75604 , n75605 , n75606 , n75607 , n75608 , n75609 , n75610 , n75611 , n75612 ,
     n75613 , n75614 , n75615 , n75616 , n75617 , n75618 , n75619 , n75620 , n75621 , n75622 ,
     n75623 , n75624 , n75625 , n75626 , n75627 , n75628 , n75629 , n75630 , n75631 , n75632 ,
     n75633 , n75634 , n75635 , n75636 , n75637 , n75638 , n75639 , n75640 , n75641 , n75642 ,
     n75643 , n75644 , n75645 , n75646 , n75647 , n75648 , n75649 , n75650 , n75651 , n75652 ,
     n75653 , n75654 , n75655 , n75656 , n75657 , n75658 , n75659 , n75660 , n75661 , n75662 ,
     n75663 , n75664 , n75665 , n75666 , n75667 , n75668 , n75669 , n75670 , n75671 , n75672 ,
     n75673 , n75674 , n75675 , n75676 , n75677 , n75678 , n75679 , n75680 , n75681 , n75682 ,
     n75683 , n75684 , n75685 , n75686 , n75687 , n75688 , n75689 , n75690 , n75691 , n75692 ,
     n75693 , n75694 , n75695 , n75696 , n75697 , n75698 , n75699 , n75700 , n75701 , n75702 ,
     n75703 , n75704 , n75705 , n75706 , n75707 , n75708 , n75709 , n75710 , n75711 , n75712 ,
     n75713 , n75714 , n75715 , n75716 , n75717 , n75718 , n75719 , n75720 , n75721 , n75722 ,
     n75723 , n75724 , n75725 , n75726 , n75727 , n75728 , n75729 , n75730 , n75731 , n75732 ,
     n75733 , n75734 , n75735 , n75736 , n75737 , n75738 , n75739 , n75740 , n75741 , n75742 ,
     n75743 , n75744 , n75745 , n75746 , n75747 , n75748 , n75749 , n75750 , n75751 , n75752 ,
     n75753 , n75754 , n75755 , n75756 , n75757 , n75758 , n75759 , n75760 , n75761 , n75762 ,
     n75763 , n75764 , n75765 , n75766 , n75767 , n75768 , n75769 , n75770 , n75771 , n75772 ,
     n75773 , n75774 , n75775 , n75776 , n75777 , n75778 , n75779 , n75780 , n75781 , n75782 ,
     n75783 , n75784 , n75785 , n75786 , n75787 , n75788 , n75789 , n75790 , n75791 , n75792 ,
     n75793 , n75794 , n75795 , n75796 , n75797 , n75798 , n75799 , n75800 , n75801 , n75802 ,
     n75803 , n75804 , n75805 , n75806 , n75807 , n75808 , n75809 , n75810 , n75811 , n75812 ,
     n75813 , n75814 , n75815 , n75816 , n75817 , n75818 , n75819 , n75820 , n75821 , n75822 ,
     n75823 , n75824 , n75825 , n75826 , n75827 , n75828 , n75829 , n75830 , n75831 , n75832 ,
     n75833 , n75834 , n75835 , n75836 , n75837 , n75838 , n75839 , n75840 , n75841 , n75842 ,
     n75843 , n75844 , n75845 , n75846 , n75847 , n75848 , n75849 , n75850 , n75851 , n75852 ,
     n75853 , n75854 , n75855 , n75856 , n75857 , n75858 , n75859 , n75860 , n75861 , n75862 ,
     n75863 , n75864 , n75865 , n75866 , n75867 , n75868 , n75869 , n75870 , n75871 , n75872 ,
     n75873 , n75874 , n75875 , n75876 , n75877 , n75878 , n75879 , n75880 , n75881 , n75882 ,
     n75883 , n75884 , n75885 , n75886 , n75887 , n75888 , n75889 , n75890 , n75891 , n75892 ,
     n75893 , n75894 , n75895 , n75896 , n75897 , n75898 , n75899 , n75900 , n75901 , n75902 ,
     n75903 , n75904 , n75905 , n75906 , n75907 , n75908 , n75909 , n75910 , n75911 , n75912 ,
     n75913 , n75914 , n75915 , n75916 , n75917 , n75918 , n75919 , n75920 , n75921 , n75922 ,
     n75923 , n75924 , n75925 , n75926 , n75927 , n75928 , n75929 , n75930 , n75931 , n75932 ,
     n75933 , n75934 , n75935 , n75936 , n75937 , n75938 , n75939 , n75940 , n75941 , n75942 ,
     n75943 , n75944 , n75945 , n75946 , n75947 , n75948 , n75949 , n75950 , n75951 , n75952 ,
     n75953 , n75954 , n75955 , n75956 , n75957 , n75958 , n75959 , n75960 , n75961 , n75962 ,
     n75963 , n75964 , n75965 , n75966 , n75967 , n75968 , n75969 , n75970 , n75971 , n75972 ,
     n75973 , n75974 , n75975 , n75976 , n75977 , n75978 , n75979 , n75980 , n75981 , n75982 ,
     n75983 , n75984 , n75985 , n75986 , n75987 , n75988 , n75989 , n75990 , n75991 , n75992 ,
     n75993 , n75994 , n75995 , n75996 , n75997 , n75998 , n75999 , n76000 , n76001 , n76002 ,
     n76003 , n76004 , n76005 , n76006 , n76007 , n76008 , n76009 , n76010 , n76011 , n76012 ,
     n76013 , n76014 , n76015 , n76016 , n76017 , n76018 , n76019 , n76020 , n76021 , n76022 ,
     n76023 , n76024 , n76025 , n76026 , n76027 , n76028 , n76029 , n76030 , n76031 , n76032 ,
     n76033 , n76034 , n76035 , n76036 , n76037 , n76038 , n76039 , n76040 , n76041 , n76042 ,
     n76043 , n76044 , n76045 , n76046 , n76047 , n76048 , n76049 , n76050 , n76051 , n76052 ,
     n76053 , n76054 , n76055 , n76056 , n76057 , n76058 , n76059 , n76060 , n76061 , n76062 ,
     n76063 , n76064 , n76065 , n76066 , n76067 , n76068 , n76069 , n76070 , n76071 , n76072 ,
     n76073 , n76074 , n76075 , n76076 , n76077 , n76078 , n76079 , n76080 , n76081 , n76082 ,
     n76083 , n76084 , n76085 , n76086 , n76087 , n76088 , n76089 , n76090 , n76091 , n76092 ,
     n76093 , n76094 , n76095 , n76096 , n76097 , n76098 , n76099 , n76100 , n76101 , n76102 ,
     n76103 , n76104 , n76105 , n76106 , n76107 , n76108 , n76109 , n76110 , n76111 , n76112 ,
     n76113 , n76114 , n76115 , n76116 , n76117 , n76118 , n76119 , n76120 , n76121 , n76122 ,
     n76123 , n76124 , n76125 , n76126 , n76127 , n76128 , n76129 , n76130 , n76131 , n76132 ,
     n76133 , n76134 , n76135 , n76136 , n76137 , n76138 , n76139 , n76140 , n76141 , n76142 ,
     n76143 , n76144 , n76145 , n76146 , n76147 , n76148 , n76149 , n76150 , n76151 , n76152 ,
     n76153 , n76154 , n76155 , n76156 , n76157 , n76158 , n76159 , n76160 , n76161 , n76162 ,
     n76163 , n76164 , n76165 , n76166 , n76167 , n76168 , n76169 , n76170 , n76171 , n76172 ,
     n76173 , n76174 , n76175 , n76176 , n76177 , n76178 , n76179 , n76180 , n76181 , n76182 ,
     n76183 , n76184 , n76185 , n76186 , n76187 , n76188 , n76189 , n76190 , n76191 , n76192 ,
     n76193 , n76194 , n76195 , n76196 , n76197 , n76198 , n76199 , n76200 , n76201 , n76202 ,
     n76203 , n76204 , n76205 , n76206 , n76207 , n76208 , n76209 , n76210 , n76211 , n76212 ,
     n76213 , n76214 , n76215 , n76216 , n76217 , n76218 , n76219 , n76220 , n76221 , n76222 ,
     n76223 , n76224 , n76225 , n76226 , n76227 , n76228 , n76229 , n76230 , n76231 , n76232 ,
     n76233 , n76234 , n76235 , n76236 , n76237 , n76238 , n76239 , n76240 , n76241 , n76242 ,
     n76243 , n76244 , n76245 , n76246 , n76247 , n76248 , n76249 , n76250 , n76251 , n76252 ,
     n76253 , n76254 , n76255 , n76256 , n76257 , n76258 , n76259 , n76260 , n76261 , n76262 ,
     n76263 , n76264 , n76265 , n76266 , n76267 , n76268 , n76269 , n76270 , n76271 , n76272 ,
     n76273 , n76274 , n76275 , n76276 , n76277 , n76278 , n76279 , n76280 , n76281 , n76282 ,
     n76283 , n76284 , n76285 , n76286 , n76287 , n76288 , n76289 , n76290 , n76291 , n76292 ,
     n76293 , n76294 , n76295 , n76296 , n76297 , n76298 , n76299 , n76300 , n76301 , n76302 ,
     n76303 , n76304 , n76305 , n76306 , n76307 , n76308 , n76309 , n76310 , n76311 , n76312 ,
     n76313 , n76314 , n76315 , n76316 , n76317 , n76318 , n76319 , n76320 , n76321 , n76322 ,
     n76323 , n76324 , n76325 , n76326 , n76327 , n76328 , n76329 , n76330 , n76331 , n76332 ,
     n76333 , n76334 , n76335 , n76336 , n76337 , n76338 , n76339 , n76340 , n76341 , n76342 ,
     n76343 , n76344 , n76345 , n76346 , n76347 , n76348 , n76349 , n76350 , n76351 , n76352 ,
     n76353 , n76354 , n76355 , n76356 , n76357 , n76358 , n76359 , n76360 , n76361 , n76362 ,
     n76363 , n76364 , n76365 , n76366 , n76367 , n76368 , n76369 , n76370 , n76371 , n76372 ,
     n76373 , n76374 , n76375 , n76376 , n76377 , n76378 , n76379 , n76380 , n76381 , n76382 ,
     n76383 , n76384 , n76385 , n76386 , n76387 , n76388 , n76389 , n76390 , n76391 , n76392 ,
     n76393 , n76394 , n76395 , n76396 , n76397 , n76398 , n76399 , n76400 , n76401 , n76402 ,
     n76403 , n76404 , n76405 , n76406 , n76407 , n76408 , n76409 , n76410 , n76411 , n76412 ,
     n76413 , n76414 , n76415 , n76416 , n76417 , n76418 , n76419 , n76420 , n76421 , n76422 ,
     n76423 , n76424 , n76425 , n76426 , n76427 , n76428 , n76429 , n76430 , n76431 , n76432 ,
     n76433 , n76434 , n76435 , n76436 , n76437 , n76438 , n76439 , n76440 , n76441 , n76442 ,
     n76443 , n76444 , n76445 , n76446 , n76447 , n76448 , n76449 , n76450 , n76451 , n76452 ,
     n76453 , n76454 , n76455 , n76456 , n76457 , n76458 , n76459 , n76460 , n76461 , n76462 ,
     n76463 , n76464 , n76465 , n76466 , n76467 , n76468 , n76469 , n76470 , n76471 , n76472 ,
     n76473 , n76474 , n76475 , n76476 , n76477 , n76478 , n76479 , n76480 , n76481 , n76482 ,
     n76483 , n76484 , n76485 , n76486 , n76487 , n76488 , n76489 , n76490 , n76491 , n76492 ,
     n76493 , n76494 , n76495 , n76496 , n76497 , n76498 , n76499 , n76500 , n76501 , n76502 ,
     n76503 , n76504 , n76505 , n76506 , n76507 , n76508 , n76509 , n76510 , n76511 , n76512 ,
     n76513 , n76514 , n76515 , n76516 , n76517 , n76518 , n76519 , n76520 , n76521 , n76522 ,
     n76523 , n76524 , n76525 , n76526 , n76527 , n76528 , n76529 , n76530 , n76531 , n76532 ,
     n76533 , n76534 , n76535 , n76536 , n76537 , n76538 , n76539 , n76540 , n76541 , n76542 ,
     n76543 , n76544 , n76545 , n76546 , n76547 , n76548 , n76549 , n76550 , n76551 , n76552 ,
     n76553 , n76554 , n76555 , n76556 , n76557 , n76558 , n76559 , n76560 , n76561 , n76562 ,
     n76563 , n76564 , n76565 , n76566 , n76567 , n76568 , n76569 , n76570 , n76571 , n76572 ,
     n76573 , n76574 , n76575 , n76576 , n76577 , n76578 , n76579 , n76580 , n76581 , n76582 ,
     n76583 , n76584 , n76585 , n76586 , n76587 , n76588 , n76589 , n76590 , n76591 , n76592 ,
     n76593 , n76594 , n76595 , n76596 , n76597 , n76598 , n76599 , n76600 , n76601 , n76602 ,
     n76603 , n76604 , n76605 , n76606 , n76607 , n76608 , n76609 , n76610 , n76611 , n76612 ,
     n76613 , n76614 , n76615 , n76616 , n76617 , n76618 , n76619 , n76620 , n76621 , n76622 ,
     n76623 , n76624 , n76625 , n76626 , n76627 , n76628 , n76629 , n76630 , n76631 , n76632 ,
     n76633 , n76634 , n76635 , n76636 , n76637 , n76638 , n76639 , n76640 , n76641 , n76642 ,
     n76643 , n76644 , n76645 , n76646 , n76647 , n76648 , n76649 , n76650 , n76651 , n76652 ,
     n76653 , n76654 , n76655 , n76656 , n76657 , n76658 , n76659 , n76660 , n76661 , n76662 ,
     n76663 , n76664 , n76665 , n76666 , n76667 , n76668 , n76669 , n76670 , n76671 , n76672 ,
     n76673 , n76674 , n76675 , n76676 , n76677 , n76678 , n76679 , n76680 , n76681 , n76682 ,
     n76683 , n76684 , n76685 , n76686 , n76687 , n76688 , n76689 , n76690 , n76691 , n76692 ,
     n76693 , n76694 , n76695 , n76696 , n76697 , n76698 , n76699 , n76700 , n76701 , n76702 ,
     n76703 , n76704 , n76705 , n76706 , n76707 , n76708 , n76709 , n76710 , n76711 , n76712 ,
     n76713 , n76714 , n76715 , n76716 , n76717 , n76718 , n76719 , n76720 , n76721 , n76722 ,
     n76723 , n76724 , n76725 , n76726 , n76727 , n76728 , n76729 , n76730 , n76731 , n76732 ,
     n76733 , n76734 , n76735 , n76736 , n76737 , n76738 , n76739 , n76740 , n76741 , n76742 ,
     n76743 , n76744 , n76745 , n76746 , n76747 , n76748 , n76749 , n76750 , n76751 , n76752 ,
     n76753 , n76754 , n76755 , n76756 , n76757 , n76758 , n76759 , n76760 , n76761 , n76762 ,
     n76763 , n76764 , n76765 , n76766 , n76767 , n76768 , n76769 , n76770 , n76771 , n76772 ,
     n76773 , n76774 , n76775 , n76776 , n76777 , n76778 , n76779 , n76780 , n76781 , n76782 ,
     n76783 , n76784 , n76785 , n76786 , n76787 , n76788 , n76789 , n76790 , n76791 , n76792 ,
     n76793 , n76794 , n76795 , n76796 , n76797 , n76798 , n76799 , n76800 , n76801 , n76802 ,
     n76803 , n76804 , n76805 , n76806 , n76807 , n76808 , n76809 , n76810 , n76811 , n76812 ,
     n76813 , n76814 , n76815 , n76816 , n76817 , n76818 , n76819 , n76820 , n76821 , n76822 ,
     n76823 , n76824 , n76825 , n76826 , n76827 , n76828 , n76829 , n76830 , n76831 , n76832 ,
     n76833 , n76834 , n76835 , n76836 , n76837 , n76838 , n76839 , n76840 , n76841 , n76842 ,
     n76843 , n76844 , n76845 , n76846 , n76847 , n76848 , n76849 , n76850 , n76851 , n76852 ,
     n76853 , n76854 , n76855 , n76856 , n76857 , n76858 , n76859 , n76860 , n76861 , n76862 ,
     n76863 , n76864 , n76865 , n76866 , n76867 , n76868 , n76869 , n76870 , n76871 , n76872 ,
     n76873 , n76874 , n76875 , n76876 , n76877 , n76878 , n76879 , n76880 , n76881 , n76882 ,
     n76883 , n76884 , n76885 , n76886 , n76887 , n76888 , n76889 , n76890 , n76891 , n76892 ,
     n76893 , n76894 , n76895 , n76896 , n76897 , n76898 , n76899 , n76900 , n76901 , n76902 ,
     n76903 , n76904 , n76905 , n76906 , n76907 , n76908 , n76909 , n76910 , n76911 , n76912 ,
     n76913 , n76914 , n76915 , n76916 , n76917 , n76918 , n76919 , n76920 , n76921 , n76922 ,
     n76923 , n76924 , n76925 , n76926 , n76927 , n76928 , n76929 , n76930 , n76931 , n76932 ,
     n76933 , n76934 , n76935 , n76936 , n76937 , n76938 , n76939 , n76940 , n76941 , n76942 ,
     n76943 , n76944 , n76945 , n76946 , n76947 , n76948 , n76949 , n76950 , n76951 , n76952 ,
     n76953 , n76954 , n76955 , n76956 , n76957 , n76958 , n76959 , n76960 , n76961 , n76962 ,
     n76963 , n76964 , n76965 , n76966 , n76967 , n76968 , n76969 , n76970 , n76971 , n76972 ,
     n76973 , n76974 , n76975 , n76976 , n76977 , n76978 , n76979 , n76980 , n76981 , n76982 ,
     n76983 , n76984 , n76985 , n76986 , n76987 , n76988 , n76989 , n76990 , n76991 , n76992 ,
     n76993 , n76994 , n76995 , n76996 , n76997 , n76998 , n76999 , n77000 , n77001 , n77002 ,
     n77003 , n77004 , n77005 , n77006 , n77007 , n77008 , n77009 , n77010 , n77011 , n77012 ,
     n77013 , n77014 , n77015 , n77016 , n77017 , n77018 , n77019 , n77020 , n77021 , n77022 ,
     n77023 , n77024 , n77025 , n77026 , n77027 , n77028 , n77029 , n77030 , n77031 , n77032 ,
     n77033 , n77034 , n77035 , n77036 , n77037 , n77038 , n77039 , n77040 , n77041 , n77042 ,
     n77043 , n77044 , n77045 , n77046 , n77047 , n77048 , n77049 , n77050 , n77051 , n77052 ,
     n77053 , n77054 , n77055 , n77056 , n77057 , n77058 , n77059 , n77060 , n77061 , n77062 ,
     n77063 , n77064 , n77065 , n77066 , n77067 , n77068 , n77069 , n77070 , n77071 , n77072 ,
     n77073 , n77074 , n77075 , n77076 , n77077 , n77078 , n77079 , n77080 , n77081 , n77082 ,
     n77083 , n77084 , n77085 , n77086 , n77087 , n77088 , n77089 , n77090 , n77091 , n77092 ,
     n77093 , n77094 , n77095 , n77096 , n77097 , n77098 , n77099 , n77100 , n77101 , n77102 ,
     n77103 , n77104 , n77105 , n77106 , n77107 , n77108 , n77109 , n77110 , n77111 , n77112 ,
     n77113 , n77114 , n77115 , n77116 , n77117 , n77118 , n77119 , n77120 , n77121 , n77122 ,
     n77123 , n77124 , n77125 , n77126 , n77127 , n77128 , n77129 , n77130 , n77131 , n77132 ,
     n77133 , n77134 , n77135 , n77136 , n77137 , n77138 , n77139 , n77140 , n77141 , n77142 ,
     n77143 , n77144 , n77145 , n77146 , n77147 , n77148 , n77149 , n77150 , n77151 , n77152 ,
     n77153 , n77154 , n77155 , n77156 , n77157 , n77158 , n77159 , n77160 , n77161 , n77162 ,
     n77163 , n77164 , n77165 , n77166 , n77167 , n77168 , n77169 , n77170 , n77171 , n77172 ,
     n77173 , n77174 , n77175 , n77176 , n77177 , n77178 , n77179 , n77180 , n77181 , n77182 ,
     n77183 , n77184 , n77185 , n77186 , n77187 , n77188 , n77189 , n77190 , n77191 , n77192 ,
     n77193 , n77194 , n77195 , n77196 , n77197 , n77198 , n77199 , n77200 , n77201 , n77202 ,
     n77203 , n77204 , n77205 , n77206 , n77207 , n77208 , n77209 , n77210 , n77211 , n77212 ,
     n77213 , n77214 , n77215 , n77216 , n77217 , n77218 , n77219 , n77220 , n77221 , n77222 ,
     n77223 , n77224 , n77225 , n77226 , n77227 , n77228 , n77229 , n77230 , n77231 , n77232 ,
     n77233 , n77234 , n77235 , n77236 , n77237 , n77238 , n77239 , n77240 , n77241 , n77242 ,
     n77243 , n77244 , n77245 , n77246 , n77247 , n77248 , n77249 , n77250 , n77251 , n77252 ,
     n77253 , n77254 , n77255 , n77256 , n77257 , n77258 , n77259 , n77260 , n77261 , n77262 ,
     n77263 , n77264 , n77265 , n77266 , n77267 , n77268 , n77269 , n77270 , n77271 , n77272 ,
     n77273 , n77274 , n77275 , n77276 , n77277 , n77278 , n77279 , n77280 , n77281 , n77282 ,
     n77283 , n77284 , n77285 , n77286 , n77287 , n77288 , n77289 , n77290 , n77291 , n77292 ,
     n77293 , n77294 , n77295 , n77296 , n77297 , n77298 , n77299 , n77300 , n77301 , n77302 ,
     n77303 , n77304 , n77305 , n77306 , n77307 , n77308 , n77309 , n77310 , n77311 , n77312 ,
     n77313 , n77314 , n77315 , n77316 , n77317 , n77318 , n77319 , n77320 , n77321 , n77322 ,
     n77323 , n77324 , n77325 , n77326 , n77327 , n77328 , n77329 , n77330 , n77331 , n77332 ,
     n77333 , n77334 , n77335 , n77336 , n77337 , n77338 , n77339 , n77340 , n77341 , n77342 ,
     n77343 , n77344 , n77345 , n77346 , n77347 , n77348 , n77349 , n77350 , n77351 , n77352 ,
     n77353 , n77354 , n77355 , n77356 , n77357 , n77358 , n77359 , n77360 , n77361 , n77362 ,
     n77363 , n77364 , n77365 , n77366 , n77367 , n77368 , n77369 , n77370 , n77371 , n77372 ,
     n77373 , n77374 , n77375 , n77376 , n77377 , n77378 , n77379 , n77380 , n77381 , n77382 ,
     n77383 , n77384 , n77385 , n77386 , n77387 , n77388 , n77389 , n77390 , n77391 , n77392 ,
     n77393 , n77394 , n77395 , n77396 , n77397 , n77398 , n77399 , n77400 , n77401 , n77402 ,
     n77403 , n77404 , n77405 , n77406 , n77407 , n77408 , n77409 , n77410 , n77411 , n77412 ,
     n77413 , n77414 , n77415 , n77416 , n77417 , n77418 , n77419 , n77420 , n77421 , n77422 ,
     n77423 , n77424 , n77425 , n77426 , n77427 , n77428 , n77429 , n77430 , n77431 , n77432 ,
     n77433 , n77434 , n77435 , n77436 , n77437 , n77438 , n77439 , n77440 , n77441 , n77442 ,
     n77443 , n77444 , n77445 , n77446 , n77447 , n77448 , n77449 , n77450 , n77451 , n77452 ,
     n77453 , n77454 , n77455 , n77456 , n77457 , n77458 , n77459 , n77460 , n77461 , n77462 ,
     n77463 , n77464 , n77465 , n77466 , n77467 , n77468 , n77469 , n77470 , n77471 , n77472 ,
     n77473 , n77474 , n77475 , n77476 , n77477 , n77478 , n77479 , n77480 , n77481 , n77482 ,
     n77483 , n77484 , n77485 , n77486 , n77487 , n77488 , n77489 , n77490 , n77491 , n77492 ,
     n77493 , n77494 , n77495 , n77496 , n77497 , n77498 , n77499 , n77500 , n77501 , n77502 ,
     n77503 , n77504 , n77505 , n77506 , n77507 , n77508 , n77509 , n77510 , n77511 , n77512 ,
     n77513 , n77514 , n77515 , n77516 , n77517 , n77518 , n77519 , n77520 , n77521 , n77522 ,
     n77523 , n77524 , n77525 , n77526 , n77527 , n77528 , n77529 , n77530 , n77531 , n77532 ,
     n77533 , n77534 , n77535 , n77536 , n77537 , n77538 , n77539 , n77540 , n77541 , n77542 ,
     n77543 , n77544 , n77545 , n77546 , n77547 , n77548 , n77549 , n77550 , n77551 , n77552 ,
     n77553 , n77554 , n77555 , n77556 , n77557 , n77558 , n77559 , n77560 , n77561 , n77562 ,
     n77563 , n77564 , n77565 , n77566 , n77567 , n77568 , n77569 , n77570 , n77571 , n77572 ,
     n77573 , n77574 , n77575 , n77576 , n77577 , n77578 , n77579 , n77580 , n77581 , n77582 ,
     n77583 , n77584 , n77585 , n77586 , n77587 , n77588 , n77589 , n77590 , n77591 , n77592 ,
     n77593 , n77594 , n77595 , n77596 , n77597 , n77598 , n77599 , n77600 , n77601 , n77602 ,
     n77603 , n77604 , n77605 , n77606 , n77607 , n77608 , n77609 , n77610 , n77611 , n77612 ,
     n77613 , n77614 , n77615 , n77616 , n77617 , n77618 , n77619 , n77620 , n77621 , n77622 ,
     n77623 , n77624 , n77625 , n77626 , n77627 , n77628 , n77629 , n77630 , n77631 , n77632 ,
     n77633 , n77634 , n77635 , n77636 , n77637 , n77638 , n77639 , n77640 , n77641 , n77642 ,
     n77643 , n77644 , n77645 , n77646 , n77647 , n77648 , n77649 , n77650 , n77651 , n77652 ,
     n77653 , n77654 , n77655 , n77656 , n77657 , n77658 , n77659 , n77660 , n77661 , n77662 ,
     n77663 , n77664 , n77665 , n77666 , n77667 , n77668 , n77669 , n77670 , n77671 , n77672 ,
     n77673 , n77674 , n77675 , n77676 , n77677 , n77678 , n77679 , n77680 , n77681 , n77682 ,
     n77683 , n77684 , n77685 , n77686 , n77687 , n77688 , n77689 , n77690 , n77691 , n77692 ,
     n77693 , n77694 , n77695 , n77696 , n77697 , n77698 , n77699 , n77700 , n77701 , n77702 ,
     n77703 , n77704 , n77705 , n77706 , n77707 , n77708 , n77709 , n77710 , n77711 , n77712 ,
     n77713 , n77714 , n77715 , n77716 , n77717 , n77718 , n77719 , n77720 , n77721 , n77722 ,
     n77723 , n77724 , n77725 , n77726 , n77727 , n77728 , n77729 , n77730 , n77731 , n77732 ,
     n77733 , n77734 , n77735 , n77736 , n77737 , n77738 , n77739 , n77740 , n77741 , n77742 ,
     n77743 , n77744 , n77745 , n77746 , n77747 , n77748 , n77749 , n77750 , n77751 , n77752 ,
     n77753 , n77754 , n77755 , n77756 , n77757 , n77758 , n77759 , n77760 , n77761 , n77762 ,
     n77763 , n77764 , n77765 , n77766 , n77767 , n77768 , n77769 , n77770 , n77771 , n77772 ,
     n77773 , n77774 , n77775 , n77776 , n77777 , n77778 , n77779 , n77780 , n77781 , n77782 ,
     n77783 , n77784 , n77785 , n77786 , n77787 , n77788 , n77789 , n77790 , n77791 , n77792 ,
     n77793 , n77794 , n77795 , n77796 , n77797 , n77798 , n77799 , n77800 , n77801 , n77802 ,
     n77803 , n77804 , n77805 , n77806 , n77807 , n77808 , n77809 , n77810 , n77811 , n77812 ,
     n77813 , n77814 , n77815 , n77816 , n77817 , n77818 , n77819 , n77820 , n77821 , n77822 ,
     n77823 , n77824 ;
buf ( n201 , n77797 );
buf ( n197 , n77800 );
buf ( n195 , n77803 );
buf ( n200 , n77806 );
buf ( n192 , n77809 );
buf ( n193 , n77812 );
buf ( n194 , n77815 );
buf ( n198 , n77818 );
buf ( n199 , n77821 );
buf ( n196 , n77824 );
buf ( n407 , n61 );
buf ( n408 , n161 );
buf ( n409 , n60 );
buf ( n410 , n8 );
buf ( n411 , n103 );
buf ( n412 , n66 );
buf ( n413 , n152 );
buf ( n414 , n42 );
buf ( n415 , n77 );
buf ( n416 , n157 );
buf ( n417 , n116 );
buf ( n418 , n82 );
buf ( n419 , n105 );
buf ( n420 , n56 );
buf ( n421 , n148 );
buf ( n422 , n188 );
buf ( n423 , n160 );
buf ( n424 , n100 );
buf ( n425 , n130 );
buf ( n426 , n83 );
buf ( n427 , n59 );
buf ( n428 , n65 );
buf ( n429 , n120 );
buf ( n430 , n54 );
buf ( n431 , n87 );
buf ( n432 , n76 );
buf ( n433 , n113 );
buf ( n434 , n104 );
buf ( n435 , n3 );
buf ( n436 , n179 );
buf ( n437 , n131 );
buf ( n438 , n93 );
buf ( n439 , n36 );
buf ( n440 , n72 );
buf ( n441 , n151 );
buf ( n442 , n89 );
buf ( n443 , n164 );
buf ( n444 , n92 );
buf ( n445 , n122 );
buf ( n446 , n51 );
buf ( n447 , n125 );
buf ( n448 , n94 );
buf ( n449 , n169 );
buf ( n450 , n123 );
buf ( n451 , n84 );
buf ( n452 , n137 );
buf ( n453 , n13 );
buf ( n454 , n86 );
buf ( n455 , n0 );
buf ( n456 , n127 );
buf ( n457 , n27 );
buf ( n458 , n190 );
buf ( n459 , n35 );
buf ( n460 , n110 );
buf ( n461 , n142 );
buf ( n462 , n166 );
buf ( n463 , n165 );
buf ( n464 , n118 );
buf ( n465 , n12 );
buf ( n466 , n73 );
buf ( n467 , n150 );
buf ( n468 , n178 );
buf ( n469 , n144 );
buf ( n470 , n187 );
buf ( n471 , n162 );
buf ( n472 , n143 );
buf ( n473 , n22 );
buf ( n474 , n180 );
buf ( n475 , n159 );
buf ( n476 , n45 );
buf ( n477 , n106 );
buf ( n478 , n49 );
buf ( n479 , n7 );
buf ( n480 , n171 );
buf ( n481 , n147 );
buf ( n482 , n133 );
buf ( n483 , n74 );
buf ( n484 , n1 );
buf ( n485 , n19 );
buf ( n486 , n29 );
buf ( n487 , n114 );
buf ( n488 , n46 );
buf ( n489 , n31 );
buf ( n490 , n139 );
buf ( n491 , n20 );
buf ( n492 , n70 );
buf ( n493 , n121 );
buf ( n494 , n134 );
buf ( n495 , n40 );
buf ( n496 , n129 );
buf ( n497 , n71 );
buf ( n498 , n173 );
buf ( n499 , n146 );
buf ( n500 , n135 );
buf ( n501 , n176 );
buf ( n502 , n158 );
buf ( n503 , n2 );
buf ( n504 , n175 );
buf ( n505 , n140 );
buf ( n506 , n163 );
buf ( n507 , n52 );
buf ( n508 , n68 );
buf ( n509 , n21 );
buf ( n510 , n5 );
buf ( n511 , n155 );
buf ( n512 , n80 );
buf ( n513 , n167 );
buf ( n514 , n108 );
buf ( n515 , n153 );
buf ( n516 , n53 );
buf ( n517 , n58 );
buf ( n518 , n128 );
buf ( n519 , n10 );
buf ( n520 , n96 );
buf ( n521 , n26 );
buf ( n522 , n14 );
buf ( n523 , n136 );
buf ( n524 , n47 );
buf ( n525 , n41 );
buf ( n526 , n95 );
buf ( n527 , n99 );
buf ( n528 , n109 );
buf ( n529 , n112 );
buf ( n530 , n37 );
buf ( n531 , n88 );
buf ( n532 , n191 );
buf ( n533 , n43 );
buf ( n534 , n124 );
buf ( n535 , n174 );
buf ( n536 , n67 );
buf ( n537 , n38 );
buf ( n538 , n138 );
buf ( n539 , n91 );
buf ( n540 , n62 );
buf ( n541 , n81 );
buf ( n542 , n9 );
buf ( n543 , n181 );
buf ( n544 , n18 );
buf ( n545 , n28 );
buf ( n546 , n168 );
buf ( n547 , n39 );
buf ( n548 , n85 );
buf ( n549 , n55 );
buf ( n550 , n24 );
buf ( n551 , n111 );
buf ( n552 , n15 );
buf ( n553 , n11 );
buf ( n554 , n33 );
buf ( n555 , n25 );
buf ( n556 , n17 );
buf ( n557 , n69 );
buf ( n558 , n154 );
buf ( n559 , n170 );
buf ( n560 , n50 );
buf ( n561 , n183 );
buf ( n562 , n145 );
buf ( n563 , n4 );
buf ( n564 , n156 );
buf ( n565 , n189 );
buf ( n566 , n16 );
buf ( n567 , n177 );
buf ( n568 , n98 );
buf ( n569 , n141 );
buf ( n570 , n186 );
buf ( n571 , n185 );
buf ( n572 , n117 );
buf ( n573 , n172 );
buf ( n574 , n63 );
buf ( n575 , n78 );
buf ( n576 , n30 );
buf ( n577 , n126 );
buf ( n578 , n149 );
buf ( n579 , n132 );
buf ( n580 , n34 );
buf ( n581 , n182 );
buf ( n582 , n6 );
buf ( n583 , n44 );
buf ( n584 , n107 );
buf ( n585 , n119 );
buf ( n586 , n101 );
buf ( n587 , n23 );
buf ( n588 , n115 );
buf ( n589 , n75 );
buf ( n590 , n57 );
buf ( n591 , n64 );
buf ( n592 , n97 );
buf ( n593 , n102 );
buf ( n594 , n79 );
buf ( n595 , n90 );
buf ( n596 , n184 );
buf ( n597 , n48 );
buf ( n598 , n32 );
buf ( n599 , n470 );
buf ( n600 , n599 );
not ( n601 , n600 );
buf ( n602 , n498 );
not ( n603 , n602 );
nor ( n604 , n601 , n603 );
buf ( n605 , n604 );
buf ( n606 , n468 );
and ( n607 , n599 , n606 );
buf ( n608 , n469 );
buf ( n609 , n608 );
xor ( n610 , n607 , n609 );
buf ( n611 , n468 );
buf ( n612 , n470 );
and ( n613 , n611 , n612 );
xor ( n614 , n610 , n613 );
buf ( n615 , n469 );
and ( n616 , n599 , n615 );
and ( n617 , n608 , n612 );
and ( n618 , n616 , n617 );
xor ( n619 , n614 , n618 );
buf ( n620 , n619 );
buf ( n621 , n620 );
not ( n622 , n621 );
buf ( n623 , n500 );
not ( n624 , n623 );
nor ( n625 , n622 , n624 );
xor ( n626 , n605 , n625 );
buf ( n627 , n626 );
and ( n628 , n607 , n609 );
and ( n629 , n609 , n613 );
and ( n630 , n607 , n613 );
or ( n631 , n628 , n629 , n630 );
buf ( n632 , n467 );
and ( n633 , n632 , n612 );
xor ( n634 , n631 , n633 );
buf ( n635 , n467 );
and ( n636 , n599 , n635 );
and ( n637 , n608 , n606 );
xor ( n638 , n636 , n637 );
and ( n639 , n611 , n615 );
xor ( n640 , n638 , n639 );
xor ( n641 , n634 , n640 );
and ( n642 , n614 , n618 );
xor ( n643 , n641 , n642 );
buf ( n644 , n643 );
buf ( n645 , n644 );
not ( n646 , n645 );
buf ( n647 , n501 );
not ( n648 , n647 );
nor ( n649 , n646 , n648 );
xor ( n650 , n627 , n649 );
buf ( n651 , n499 );
not ( n652 , n651 );
nor ( n653 , n601 , n652 );
buf ( n654 , n653 );
nor ( n655 , n622 , n648 );
and ( n656 , n654 , n655 );
buf ( n657 , n656 );
xor ( n658 , n650 , n657 );
and ( n659 , n636 , n637 );
and ( n660 , n637 , n639 );
and ( n661 , n636 , n639 );
or ( n662 , n659 , n660 , n661 );
buf ( n663 , n466 );
and ( n664 , n599 , n663 );
and ( n665 , n608 , n635 );
xor ( n666 , n664 , n665 );
buf ( n667 , n611 );
xor ( n668 , n666 , n667 );
xor ( n669 , n662 , n668 );
and ( n670 , n632 , n615 );
buf ( n671 , n466 );
and ( n672 , n671 , n612 );
xor ( n673 , n670 , n672 );
xor ( n674 , n669 , n673 );
and ( n675 , n631 , n633 );
and ( n676 , n633 , n640 );
and ( n677 , n631 , n640 );
or ( n678 , n675 , n676 , n677 );
xor ( n679 , n674 , n678 );
and ( n680 , n641 , n642 );
xor ( n681 , n679 , n680 );
buf ( n682 , n681 );
buf ( n683 , n682 );
not ( n684 , n683 );
buf ( n685 , n502 );
not ( n686 , n685 );
nor ( n687 , n684 , n686 );
xor ( n688 , n658 , n687 );
xor ( n689 , n654 , n655 );
buf ( n690 , n689 );
nor ( n691 , n646 , n686 );
and ( n692 , n690 , n691 );
xor ( n693 , n690 , n691 );
nor ( n694 , n601 , n624 );
buf ( n695 , n694 );
nor ( n696 , n622 , n686 );
and ( n697 , n695 , n696 );
buf ( n698 , n697 );
and ( n699 , n693 , n698 );
or ( n700 , n692 , n699 );
xor ( n701 , n688 , n700 );
and ( n702 , n670 , n672 );
and ( n703 , n662 , n668 );
and ( n704 , n668 , n673 );
and ( n705 , n662 , n673 );
or ( n706 , n703 , n704 , n705 );
xor ( n707 , n702 , n706 );
and ( n708 , n664 , n665 );
and ( n709 , n665 , n667 );
and ( n710 , n664 , n667 );
or ( n711 , n708 , n709 , n710 );
and ( n712 , n632 , n606 );
and ( n713 , n671 , n615 );
xor ( n714 , n712 , n713 );
buf ( n715 , n465 );
and ( n716 , n715 , n612 );
xor ( n717 , n714 , n716 );
xor ( n718 , n711 , n717 );
buf ( n719 , n465 );
and ( n720 , n599 , n719 );
and ( n721 , n608 , n663 );
xor ( n722 , n720 , n721 );
and ( n723 , n611 , n635 );
xor ( n724 , n722 , n723 );
xor ( n725 , n718 , n724 );
xor ( n726 , n707 , n725 );
and ( n727 , n674 , n678 );
and ( n728 , n679 , n680 );
or ( n729 , n727 , n728 );
xor ( n730 , n726 , n729 );
buf ( n731 , n730 );
buf ( n732 , n731 );
not ( n733 , n732 );
buf ( n734 , n503 );
not ( n735 , n734 );
nor ( n736 , n733 , n735 );
xor ( n737 , n701 , n736 );
xor ( n738 , n693 , n698 );
nor ( n739 , n684 , n735 );
and ( n740 , n738 , n739 );
xor ( n741 , n738 , n739 );
xor ( n742 , n695 , n696 );
buf ( n743 , n742 );
nor ( n744 , n646 , n735 );
and ( n745 , n743 , n744 );
xor ( n746 , n743 , n744 );
nor ( n747 , n601 , n648 );
buf ( n748 , n747 );
nor ( n749 , n622 , n735 );
and ( n750 , n748 , n749 );
buf ( n751 , n750 );
and ( n752 , n746 , n751 );
or ( n753 , n745 , n752 );
and ( n754 , n741 , n753 );
or ( n755 , n740 , n754 );
xor ( n756 , n737 , n755 );
and ( n757 , n711 , n717 );
and ( n758 , n717 , n724 );
and ( n759 , n711 , n724 );
or ( n760 , n757 , n758 , n759 );
and ( n761 , n720 , n721 );
and ( n762 , n721 , n723 );
and ( n763 , n720 , n723 );
or ( n764 , n761 , n762 , n763 );
buf ( n765 , n632 );
and ( n766 , n671 , n606 );
xor ( n767 , n765 , n766 );
and ( n768 , n715 , n615 );
xor ( n769 , n767 , n768 );
xor ( n770 , n764 , n769 );
buf ( n771 , n464 );
and ( n772 , n599 , n771 );
and ( n773 , n608 , n719 );
xor ( n774 , n772 , n773 );
and ( n775 , n611 , n663 );
xor ( n776 , n774 , n775 );
xor ( n777 , n770 , n776 );
xor ( n778 , n760 , n777 );
and ( n779 , n712 , n713 );
and ( n780 , n713 , n716 );
and ( n781 , n712 , n716 );
or ( n782 , n779 , n780 , n781 );
buf ( n783 , n464 );
and ( n784 , n783 , n612 );
xor ( n785 , n782 , n784 );
xor ( n786 , n778 , n785 );
and ( n787 , n702 , n706 );
and ( n788 , n706 , n725 );
and ( n789 , n702 , n725 );
or ( n790 , n787 , n788 , n789 );
xor ( n791 , n786 , n790 );
and ( n792 , n726 , n729 );
xor ( n793 , n791 , n792 );
buf ( n794 , n793 );
buf ( n795 , n794 );
not ( n796 , n795 );
buf ( n797 , n504 );
not ( n798 , n797 );
nor ( n799 , n796 , n798 );
xor ( n800 , n756 , n799 );
xor ( n801 , n741 , n753 );
nor ( n802 , n733 , n798 );
and ( n803 , n801 , n802 );
xor ( n804 , n801 , n802 );
xor ( n805 , n746 , n751 );
nor ( n806 , n684 , n798 );
and ( n807 , n805 , n806 );
xor ( n808 , n805 , n806 );
xor ( n809 , n748 , n749 );
buf ( n810 , n809 );
nor ( n811 , n646 , n798 );
and ( n812 , n810 , n811 );
xor ( n813 , n810 , n811 );
nor ( n814 , n601 , n686 );
buf ( n815 , n814 );
nor ( n816 , n622 , n798 );
and ( n817 , n815 , n816 );
buf ( n818 , n817 );
and ( n819 , n813 , n818 );
or ( n820 , n812 , n819 );
and ( n821 , n808 , n820 );
or ( n822 , n807 , n821 );
and ( n823 , n804 , n822 );
or ( n824 , n803 , n823 );
xor ( n825 , n800 , n824 );
and ( n826 , n782 , n784 );
and ( n827 , n760 , n777 );
and ( n828 , n777 , n785 );
and ( n829 , n760 , n785 );
or ( n830 , n827 , n828 , n829 );
xor ( n831 , n826 , n830 );
and ( n832 , n764 , n769 );
and ( n833 , n769 , n776 );
and ( n834 , n764 , n776 );
or ( n835 , n832 , n833 , n834 );
and ( n836 , n772 , n773 );
and ( n837 , n773 , n775 );
and ( n838 , n772 , n775 );
or ( n839 , n836 , n837 , n838 );
buf ( n840 , n463 );
and ( n841 , n599 , n840 );
and ( n842 , n608 , n771 );
xor ( n843 , n841 , n842 );
and ( n844 , n611 , n719 );
xor ( n845 , n843 , n844 );
xor ( n846 , n839 , n845 );
and ( n847 , n715 , n606 );
buf ( n848 , n847 );
xor ( n849 , n846 , n848 );
xor ( n850 , n835 , n849 );
and ( n851 , n765 , n766 );
and ( n852 , n766 , n768 );
and ( n853 , n765 , n768 );
or ( n854 , n851 , n852 , n853 );
and ( n855 , n783 , n615 );
buf ( n856 , n463 );
and ( n857 , n856 , n612 );
xor ( n858 , n855 , n857 );
xor ( n859 , n854 , n858 );
xor ( n860 , n850 , n859 );
xor ( n861 , n831 , n860 );
and ( n862 , n786 , n790 );
and ( n863 , n791 , n792 );
or ( n864 , n862 , n863 );
xor ( n865 , n861 , n864 );
buf ( n866 , n865 );
buf ( n867 , n866 );
not ( n868 , n867 );
buf ( n869 , n505 );
not ( n870 , n869 );
nor ( n871 , n868 , n870 );
xor ( n872 , n825 , n871 );
xor ( n873 , n804 , n822 );
nor ( n874 , n796 , n870 );
and ( n875 , n873 , n874 );
xor ( n876 , n873 , n874 );
xor ( n877 , n808 , n820 );
nor ( n878 , n733 , n870 );
and ( n879 , n877 , n878 );
xor ( n880 , n877 , n878 );
xor ( n881 , n813 , n818 );
nor ( n882 , n684 , n870 );
and ( n883 , n881 , n882 );
xor ( n884 , n881 , n882 );
xor ( n885 , n815 , n816 );
buf ( n886 , n885 );
nor ( n887 , n646 , n870 );
and ( n888 , n886 , n887 );
xor ( n889 , n886 , n887 );
nor ( n890 , n601 , n735 );
buf ( n891 , n890 );
nor ( n892 , n622 , n870 );
and ( n893 , n891 , n892 );
buf ( n894 , n893 );
and ( n895 , n889 , n894 );
or ( n896 , n888 , n895 );
and ( n897 , n884 , n896 );
or ( n898 , n883 , n897 );
and ( n899 , n880 , n898 );
or ( n900 , n879 , n899 );
and ( n901 , n876 , n900 );
or ( n902 , n875 , n901 );
xor ( n903 , n872 , n902 );
and ( n904 , n854 , n858 );
and ( n905 , n835 , n849 );
and ( n906 , n849 , n859 );
and ( n907 , n835 , n859 );
or ( n908 , n905 , n906 , n907 );
xor ( n909 , n904 , n908 );
and ( n910 , n839 , n845 );
and ( n911 , n845 , n848 );
and ( n912 , n839 , n848 );
or ( n913 , n910 , n911 , n912 );
and ( n914 , n632 , n663 );
and ( n915 , n671 , n635 );
and ( n916 , n914 , n915 );
and ( n917 , n915 , n847 );
and ( n918 , n914 , n847 );
or ( n919 , n916 , n917 , n918 );
and ( n920 , n855 , n857 );
xor ( n921 , n919 , n920 );
and ( n922 , n783 , n606 );
and ( n923 , n856 , n615 );
xor ( n924 , n922 , n923 );
buf ( n925 , n462 );
and ( n926 , n925 , n612 );
xor ( n927 , n924 , n926 );
xor ( n928 , n921 , n927 );
xor ( n929 , n913 , n928 );
and ( n930 , n841 , n842 );
and ( n931 , n842 , n844 );
and ( n932 , n841 , n844 );
or ( n933 , n930 , n931 , n932 );
and ( n934 , n632 , n719 );
buf ( n935 , n671 );
xor ( n936 , n934 , n935 );
and ( n937 , n715 , n635 );
xor ( n938 , n936 , n937 );
xor ( n939 , n933 , n938 );
buf ( n940 , n462 );
and ( n941 , n599 , n940 );
and ( n942 , n608 , n840 );
xor ( n943 , n941 , n942 );
and ( n944 , n611 , n771 );
xor ( n945 , n943 , n944 );
xor ( n946 , n939 , n945 );
xor ( n947 , n929 , n946 );
xor ( n948 , n909 , n947 );
and ( n949 , n826 , n830 );
and ( n950 , n830 , n860 );
and ( n951 , n826 , n860 );
or ( n952 , n949 , n950 , n951 );
xor ( n953 , n948 , n952 );
and ( n954 , n861 , n864 );
xor ( n955 , n953 , n954 );
buf ( n956 , n955 );
buf ( n957 , n956 );
not ( n958 , n957 );
buf ( n959 , n506 );
not ( n960 , n959 );
nor ( n961 , n958 , n960 );
xor ( n962 , n903 , n961 );
xor ( n963 , n876 , n900 );
nor ( n964 , n868 , n960 );
and ( n965 , n963 , n964 );
xor ( n966 , n963 , n964 );
xor ( n967 , n880 , n898 );
nor ( n968 , n796 , n960 );
and ( n969 , n967 , n968 );
xor ( n970 , n967 , n968 );
xor ( n971 , n884 , n896 );
nor ( n972 , n733 , n960 );
and ( n973 , n971 , n972 );
xor ( n974 , n971 , n972 );
xor ( n975 , n889 , n894 );
nor ( n976 , n684 , n960 );
and ( n977 , n975 , n976 );
xor ( n978 , n975 , n976 );
xor ( n979 , n891 , n892 );
buf ( n980 , n979 );
nor ( n981 , n646 , n960 );
and ( n982 , n980 , n981 );
xor ( n983 , n980 , n981 );
nor ( n984 , n601 , n798 );
buf ( n985 , n984 );
nor ( n986 , n622 , n960 );
and ( n987 , n985 , n986 );
buf ( n988 , n987 );
and ( n989 , n983 , n988 );
or ( n990 , n982 , n989 );
and ( n991 , n978 , n990 );
or ( n992 , n977 , n991 );
and ( n993 , n974 , n992 );
or ( n994 , n973 , n993 );
and ( n995 , n970 , n994 );
or ( n996 , n969 , n995 );
and ( n997 , n966 , n996 );
or ( n998 , n965 , n997 );
xor ( n999 , n962 , n998 );
and ( n1000 , n913 , n928 );
and ( n1001 , n928 , n946 );
and ( n1002 , n913 , n946 );
or ( n1003 , n1000 , n1001 , n1002 );
and ( n1004 , n933 , n938 );
and ( n1005 , n938 , n945 );
and ( n1006 , n933 , n945 );
or ( n1007 , n1004 , n1005 , n1006 );
and ( n1008 , n922 , n923 );
and ( n1009 , n923 , n926 );
and ( n1010 , n922 , n926 );
or ( n1011 , n1008 , n1009 , n1010 );
and ( n1012 , n934 , n935 );
and ( n1013 , n935 , n937 );
and ( n1014 , n934 , n937 );
or ( n1015 , n1012 , n1013 , n1014 );
xor ( n1016 , n1011 , n1015 );
and ( n1017 , n783 , n635 );
and ( n1018 , n856 , n606 );
xor ( n1019 , n1017 , n1018 );
and ( n1020 , n925 , n615 );
xor ( n1021 , n1019 , n1020 );
xor ( n1022 , n1016 , n1021 );
xor ( n1023 , n1007 , n1022 );
and ( n1024 , n941 , n942 );
and ( n1025 , n942 , n944 );
and ( n1026 , n941 , n944 );
or ( n1027 , n1024 , n1025 , n1026 );
and ( n1028 , n632 , n771 );
and ( n1029 , n671 , n719 );
xor ( n1030 , n1028 , n1029 );
and ( n1031 , n715 , n663 );
xor ( n1032 , n1030 , n1031 );
xor ( n1033 , n1027 , n1032 );
buf ( n1034 , n461 );
and ( n1035 , n599 , n1034 );
and ( n1036 , n608 , n940 );
xor ( n1037 , n1035 , n1036 );
and ( n1038 , n611 , n840 );
xor ( n1039 , n1037 , n1038 );
xor ( n1040 , n1033 , n1039 );
xor ( n1041 , n1023 , n1040 );
xor ( n1042 , n1003 , n1041 );
and ( n1043 , n919 , n920 );
and ( n1044 , n920 , n927 );
and ( n1045 , n919 , n927 );
or ( n1046 , n1043 , n1044 , n1045 );
buf ( n1047 , n461 );
and ( n1048 , n1047 , n612 );
xor ( n1049 , n1046 , n1048 );
xor ( n1050 , n1042 , n1049 );
and ( n1051 , n904 , n908 );
and ( n1052 , n908 , n947 );
and ( n1053 , n904 , n947 );
or ( n1054 , n1051 , n1052 , n1053 );
xor ( n1055 , n1050 , n1054 );
and ( n1056 , n948 , n952 );
and ( n1057 , n953 , n954 );
or ( n1058 , n1056 , n1057 );
xor ( n1059 , n1055 , n1058 );
buf ( n1060 , n1059 );
buf ( n1061 , n1060 );
not ( n1062 , n1061 );
buf ( n1063 , n507 );
not ( n1064 , n1063 );
nor ( n1065 , n1062 , n1064 );
xor ( n1066 , n999 , n1065 );
xor ( n1067 , n966 , n996 );
nor ( n1068 , n958 , n1064 );
and ( n1069 , n1067 , n1068 );
xor ( n1070 , n1067 , n1068 );
xor ( n1071 , n970 , n994 );
nor ( n1072 , n868 , n1064 );
and ( n1073 , n1071 , n1072 );
xor ( n1074 , n1071 , n1072 );
xor ( n1075 , n974 , n992 );
nor ( n1076 , n796 , n1064 );
and ( n1077 , n1075 , n1076 );
xor ( n1078 , n1075 , n1076 );
xor ( n1079 , n978 , n990 );
nor ( n1080 , n733 , n1064 );
and ( n1081 , n1079 , n1080 );
xor ( n1082 , n1079 , n1080 );
xor ( n1083 , n983 , n988 );
nor ( n1084 , n684 , n1064 );
and ( n1085 , n1083 , n1084 );
xor ( n1086 , n1083 , n1084 );
xor ( n1087 , n985 , n986 );
buf ( n1088 , n1087 );
nor ( n1089 , n646 , n1064 );
and ( n1090 , n1088 , n1089 );
xor ( n1091 , n1088 , n1089 );
nor ( n1092 , n601 , n870 );
buf ( n1093 , n1092 );
nor ( n1094 , n622 , n1064 );
and ( n1095 , n1093 , n1094 );
buf ( n1096 , n1095 );
and ( n1097 , n1091 , n1096 );
or ( n1098 , n1090 , n1097 );
and ( n1099 , n1086 , n1098 );
or ( n1100 , n1085 , n1099 );
and ( n1101 , n1082 , n1100 );
or ( n1102 , n1081 , n1101 );
and ( n1103 , n1078 , n1102 );
or ( n1104 , n1077 , n1103 );
and ( n1105 , n1074 , n1104 );
or ( n1106 , n1073 , n1105 );
and ( n1107 , n1070 , n1106 );
or ( n1108 , n1069 , n1107 );
xor ( n1109 , n1066 , n1108 );
and ( n1110 , n1046 , n1048 );
and ( n1111 , n1003 , n1041 );
and ( n1112 , n1041 , n1049 );
and ( n1113 , n1003 , n1049 );
or ( n1114 , n1111 , n1112 , n1113 );
xor ( n1115 , n1110 , n1114 );
and ( n1116 , n1007 , n1022 );
and ( n1117 , n1022 , n1040 );
and ( n1118 , n1007 , n1040 );
or ( n1119 , n1116 , n1117 , n1118 );
and ( n1120 , n1027 , n1032 );
and ( n1121 , n1032 , n1039 );
and ( n1122 , n1027 , n1039 );
or ( n1123 , n1120 , n1121 , n1122 );
and ( n1124 , n1035 , n1036 );
and ( n1125 , n1036 , n1038 );
and ( n1126 , n1035 , n1038 );
or ( n1127 , n1124 , n1125 , n1126 );
and ( n1128 , n632 , n840 );
and ( n1129 , n671 , n771 );
xor ( n1130 , n1128 , n1129 );
buf ( n1131 , n715 );
xor ( n1132 , n1130 , n1131 );
xor ( n1133 , n1127 , n1132 );
buf ( n1134 , n460 );
and ( n1135 , n599 , n1134 );
and ( n1136 , n608 , n1034 );
xor ( n1137 , n1135 , n1136 );
and ( n1138 , n611 , n940 );
xor ( n1139 , n1137 , n1138 );
xor ( n1140 , n1133 , n1139 );
xor ( n1141 , n1123 , n1140 );
and ( n1142 , n1017 , n1018 );
and ( n1143 , n1018 , n1020 );
and ( n1144 , n1017 , n1020 );
or ( n1145 , n1142 , n1143 , n1144 );
and ( n1146 , n1028 , n1029 );
and ( n1147 , n1029 , n1031 );
and ( n1148 , n1028 , n1031 );
or ( n1149 , n1146 , n1147 , n1148 );
xor ( n1150 , n1145 , n1149 );
and ( n1151 , n783 , n663 );
and ( n1152 , n856 , n635 );
xor ( n1153 , n1151 , n1152 );
and ( n1154 , n925 , n606 );
xor ( n1155 , n1153 , n1154 );
xor ( n1156 , n1150 , n1155 );
xor ( n1157 , n1141 , n1156 );
xor ( n1158 , n1119 , n1157 );
and ( n1159 , n1011 , n1015 );
and ( n1160 , n1015 , n1021 );
and ( n1161 , n1011 , n1021 );
or ( n1162 , n1159 , n1160 , n1161 );
and ( n1163 , n1047 , n615 );
buf ( n1164 , n460 );
and ( n1165 , n1164 , n612 );
xor ( n1166 , n1163 , n1165 );
xor ( n1167 , n1162 , n1166 );
xor ( n1168 , n1158 , n1167 );
xor ( n1169 , n1115 , n1168 );
and ( n1170 , n1050 , n1054 );
and ( n1171 , n1055 , n1058 );
or ( n1172 , n1170 , n1171 );
xor ( n1173 , n1169 , n1172 );
buf ( n1174 , n1173 );
buf ( n1175 , n1174 );
not ( n1176 , n1175 );
buf ( n1177 , n508 );
not ( n1178 , n1177 );
nor ( n1179 , n1176 , n1178 );
xor ( n1180 , n1109 , n1179 );
xor ( n1181 , n1070 , n1106 );
nor ( n1182 , n1062 , n1178 );
and ( n1183 , n1181 , n1182 );
xor ( n1184 , n1181 , n1182 );
xor ( n1185 , n1074 , n1104 );
nor ( n1186 , n958 , n1178 );
and ( n1187 , n1185 , n1186 );
xor ( n1188 , n1185 , n1186 );
xor ( n1189 , n1078 , n1102 );
nor ( n1190 , n868 , n1178 );
and ( n1191 , n1189 , n1190 );
xor ( n1192 , n1189 , n1190 );
xor ( n1193 , n1082 , n1100 );
nor ( n1194 , n796 , n1178 );
and ( n1195 , n1193 , n1194 );
xor ( n1196 , n1193 , n1194 );
xor ( n1197 , n1086 , n1098 );
nor ( n1198 , n733 , n1178 );
and ( n1199 , n1197 , n1198 );
xor ( n1200 , n1197 , n1198 );
xor ( n1201 , n1091 , n1096 );
nor ( n1202 , n684 , n1178 );
and ( n1203 , n1201 , n1202 );
xor ( n1204 , n1201 , n1202 );
xor ( n1205 , n1093 , n1094 );
buf ( n1206 , n1205 );
nor ( n1207 , n646 , n1178 );
and ( n1208 , n1206 , n1207 );
xor ( n1209 , n1206 , n1207 );
nor ( n1210 , n601 , n960 );
buf ( n1211 , n1210 );
nor ( n1212 , n622 , n1178 );
and ( n1213 , n1211 , n1212 );
buf ( n1214 , n1213 );
and ( n1215 , n1209 , n1214 );
or ( n1216 , n1208 , n1215 );
and ( n1217 , n1204 , n1216 );
or ( n1218 , n1203 , n1217 );
and ( n1219 , n1200 , n1218 );
or ( n1220 , n1199 , n1219 );
and ( n1221 , n1196 , n1220 );
or ( n1222 , n1195 , n1221 );
and ( n1223 , n1192 , n1222 );
or ( n1224 , n1191 , n1223 );
and ( n1225 , n1188 , n1224 );
or ( n1226 , n1187 , n1225 );
and ( n1227 , n1184 , n1226 );
or ( n1228 , n1183 , n1227 );
xor ( n1229 , n1180 , n1228 );
and ( n1230 , n1162 , n1166 );
and ( n1231 , n1119 , n1157 );
and ( n1232 , n1157 , n1167 );
and ( n1233 , n1119 , n1167 );
or ( n1234 , n1231 , n1232 , n1233 );
xor ( n1235 , n1230 , n1234 );
and ( n1236 , n1123 , n1140 );
and ( n1237 , n1140 , n1156 );
and ( n1238 , n1123 , n1156 );
or ( n1239 , n1236 , n1237 , n1238 );
and ( n1240 , n1127 , n1132 );
and ( n1241 , n1132 , n1139 );
and ( n1242 , n1127 , n1139 );
or ( n1243 , n1240 , n1241 , n1242 );
and ( n1244 , n1135 , n1136 );
and ( n1245 , n1136 , n1138 );
and ( n1246 , n1135 , n1138 );
or ( n1247 , n1244 , n1245 , n1246 );
and ( n1248 , n632 , n940 );
and ( n1249 , n671 , n840 );
xor ( n1250 , n1248 , n1249 );
and ( n1251 , n715 , n771 );
xor ( n1252 , n1250 , n1251 );
xor ( n1253 , n1247 , n1252 );
buf ( n1254 , n459 );
and ( n1255 , n599 , n1254 );
and ( n1256 , n608 , n1134 );
xor ( n1257 , n1255 , n1256 );
and ( n1258 , n611 , n1034 );
xor ( n1259 , n1257 , n1258 );
xor ( n1260 , n1253 , n1259 );
xor ( n1261 , n1243 , n1260 );
and ( n1262 , n1128 , n1129 );
and ( n1263 , n1129 , n1131 );
and ( n1264 , n1128 , n1131 );
or ( n1265 , n1262 , n1263 , n1264 );
and ( n1266 , n1151 , n1152 );
and ( n1267 , n1152 , n1154 );
and ( n1268 , n1151 , n1154 );
or ( n1269 , n1266 , n1267 , n1268 );
xor ( n1270 , n1265 , n1269 );
and ( n1271 , n783 , n719 );
and ( n1272 , n856 , n663 );
xor ( n1273 , n1271 , n1272 );
and ( n1274 , n925 , n635 );
xor ( n1275 , n1273 , n1274 );
xor ( n1276 , n1270 , n1275 );
xor ( n1277 , n1261 , n1276 );
xor ( n1278 , n1239 , n1277 );
and ( n1279 , n1145 , n1149 );
and ( n1280 , n1149 , n1155 );
and ( n1281 , n1145 , n1155 );
or ( n1282 , n1279 , n1280 , n1281 );
and ( n1283 , n1163 , n1165 );
and ( n1284 , n1047 , n606 );
and ( n1285 , n1164 , n615 );
xor ( n1286 , n1284 , n1285 );
buf ( n1287 , n459 );
and ( n1288 , n1287 , n612 );
xor ( n1289 , n1286 , n1288 );
xor ( n1290 , n1283 , n1289 );
xor ( n1291 , n1282 , n1290 );
xor ( n1292 , n1278 , n1291 );
xor ( n1293 , n1235 , n1292 );
and ( n1294 , n1110 , n1114 );
and ( n1295 , n1114 , n1168 );
and ( n1296 , n1110 , n1168 );
or ( n1297 , n1294 , n1295 , n1296 );
xor ( n1298 , n1293 , n1297 );
and ( n1299 , n1169 , n1172 );
xor ( n1300 , n1298 , n1299 );
buf ( n1301 , n1300 );
buf ( n1302 , n1301 );
not ( n1303 , n1302 );
buf ( n1304 , n509 );
not ( n1305 , n1304 );
nor ( n1306 , n1303 , n1305 );
xor ( n1307 , n1229 , n1306 );
xor ( n1308 , n1184 , n1226 );
nor ( n1309 , n1176 , n1305 );
and ( n1310 , n1308 , n1309 );
xor ( n1311 , n1308 , n1309 );
xor ( n1312 , n1188 , n1224 );
nor ( n1313 , n1062 , n1305 );
and ( n1314 , n1312 , n1313 );
xor ( n1315 , n1312 , n1313 );
xor ( n1316 , n1192 , n1222 );
nor ( n1317 , n958 , n1305 );
and ( n1318 , n1316 , n1317 );
xor ( n1319 , n1316 , n1317 );
xor ( n1320 , n1196 , n1220 );
nor ( n1321 , n868 , n1305 );
and ( n1322 , n1320 , n1321 );
xor ( n1323 , n1320 , n1321 );
xor ( n1324 , n1200 , n1218 );
nor ( n1325 , n796 , n1305 );
and ( n1326 , n1324 , n1325 );
xor ( n1327 , n1324 , n1325 );
xor ( n1328 , n1204 , n1216 );
nor ( n1329 , n733 , n1305 );
and ( n1330 , n1328 , n1329 );
xor ( n1331 , n1328 , n1329 );
xor ( n1332 , n1209 , n1214 );
nor ( n1333 , n684 , n1305 );
and ( n1334 , n1332 , n1333 );
xor ( n1335 , n1332 , n1333 );
xor ( n1336 , n1211 , n1212 );
buf ( n1337 , n1336 );
nor ( n1338 , n646 , n1305 );
and ( n1339 , n1337 , n1338 );
xor ( n1340 , n1337 , n1338 );
nor ( n1341 , n601 , n1064 );
buf ( n1342 , n1341 );
nor ( n1343 , n622 , n1305 );
and ( n1344 , n1342 , n1343 );
buf ( n1345 , n1344 );
and ( n1346 , n1340 , n1345 );
or ( n1347 , n1339 , n1346 );
and ( n1348 , n1335 , n1347 );
or ( n1349 , n1334 , n1348 );
and ( n1350 , n1331 , n1349 );
or ( n1351 , n1330 , n1350 );
and ( n1352 , n1327 , n1351 );
or ( n1353 , n1326 , n1352 );
and ( n1354 , n1323 , n1353 );
or ( n1355 , n1322 , n1354 );
and ( n1356 , n1319 , n1355 );
or ( n1357 , n1318 , n1356 );
and ( n1358 , n1315 , n1357 );
or ( n1359 , n1314 , n1358 );
and ( n1360 , n1311 , n1359 );
or ( n1361 , n1310 , n1360 );
xor ( n1362 , n1307 , n1361 );
and ( n1363 , n1282 , n1290 );
and ( n1364 , n1239 , n1277 );
and ( n1365 , n1277 , n1291 );
and ( n1366 , n1239 , n1291 );
or ( n1367 , n1364 , n1365 , n1366 );
xor ( n1368 , n1363 , n1367 );
and ( n1369 , n1243 , n1260 );
and ( n1370 , n1260 , n1276 );
and ( n1371 , n1243 , n1276 );
or ( n1372 , n1369 , n1370 , n1371 );
and ( n1373 , n1265 , n1269 );
and ( n1374 , n1269 , n1275 );
and ( n1375 , n1265 , n1275 );
or ( n1376 , n1373 , n1374 , n1375 );
and ( n1377 , n1283 , n1289 );
xor ( n1378 , n1376 , n1377 );
and ( n1379 , n1284 , n1285 );
and ( n1380 , n1285 , n1288 );
and ( n1381 , n1284 , n1288 );
or ( n1382 , n1379 , n1380 , n1381 );
buf ( n1383 , n458 );
and ( n1384 , n1383 , n612 );
xor ( n1385 , n1382 , n1384 );
and ( n1386 , n1047 , n635 );
and ( n1387 , n1164 , n606 );
xor ( n1388 , n1386 , n1387 );
and ( n1389 , n1287 , n615 );
xor ( n1390 , n1388 , n1389 );
xor ( n1391 , n1385 , n1390 );
xor ( n1392 , n1378 , n1391 );
xor ( n1393 , n1372 , n1392 );
and ( n1394 , n1247 , n1252 );
and ( n1395 , n1252 , n1259 );
and ( n1396 , n1247 , n1259 );
or ( n1397 , n1394 , n1395 , n1396 );
and ( n1398 , n1271 , n1272 );
and ( n1399 , n1272 , n1274 );
and ( n1400 , n1271 , n1274 );
or ( n1401 , n1398 , n1399 , n1400 );
and ( n1402 , n1248 , n1249 );
and ( n1403 , n1249 , n1251 );
and ( n1404 , n1248 , n1251 );
or ( n1405 , n1402 , n1403 , n1404 );
xor ( n1406 , n1401 , n1405 );
buf ( n1407 , n783 );
and ( n1408 , n856 , n719 );
xor ( n1409 , n1407 , n1408 );
and ( n1410 , n925 , n663 );
xor ( n1411 , n1409 , n1410 );
xor ( n1412 , n1406 , n1411 );
xor ( n1413 , n1397 , n1412 );
and ( n1414 , n1255 , n1256 );
and ( n1415 , n1256 , n1258 );
and ( n1416 , n1255 , n1258 );
or ( n1417 , n1414 , n1415 , n1416 );
and ( n1418 , n632 , n1034 );
and ( n1419 , n671 , n940 );
xor ( n1420 , n1418 , n1419 );
and ( n1421 , n715 , n840 );
xor ( n1422 , n1420 , n1421 );
xor ( n1423 , n1417 , n1422 );
buf ( n1424 , n458 );
and ( n1425 , n599 , n1424 );
and ( n1426 , n608 , n1254 );
xor ( n1427 , n1425 , n1426 );
and ( n1428 , n611 , n1134 );
xor ( n1429 , n1427 , n1428 );
xor ( n1430 , n1423 , n1429 );
xor ( n1431 , n1413 , n1430 );
xor ( n1432 , n1393 , n1431 );
xor ( n1433 , n1368 , n1432 );
and ( n1434 , n1230 , n1234 );
and ( n1435 , n1234 , n1292 );
and ( n1436 , n1230 , n1292 );
or ( n1437 , n1434 , n1435 , n1436 );
xor ( n1438 , n1433 , n1437 );
and ( n1439 , n1293 , n1297 );
and ( n1440 , n1298 , n1299 );
or ( n1441 , n1439 , n1440 );
xor ( n1442 , n1438 , n1441 );
buf ( n1443 , n1442 );
buf ( n1444 , n1443 );
not ( n1445 , n1444 );
buf ( n1446 , n510 );
not ( n1447 , n1446 );
nor ( n1448 , n1445 , n1447 );
xor ( n1449 , n1362 , n1448 );
xor ( n1450 , n1311 , n1359 );
nor ( n1451 , n1303 , n1447 );
and ( n1452 , n1450 , n1451 );
xor ( n1453 , n1450 , n1451 );
xor ( n1454 , n1315 , n1357 );
nor ( n1455 , n1176 , n1447 );
and ( n1456 , n1454 , n1455 );
xor ( n1457 , n1454 , n1455 );
xor ( n1458 , n1319 , n1355 );
nor ( n1459 , n1062 , n1447 );
and ( n1460 , n1458 , n1459 );
xor ( n1461 , n1458 , n1459 );
xor ( n1462 , n1323 , n1353 );
nor ( n1463 , n958 , n1447 );
and ( n1464 , n1462 , n1463 );
xor ( n1465 , n1462 , n1463 );
xor ( n1466 , n1327 , n1351 );
nor ( n1467 , n868 , n1447 );
and ( n1468 , n1466 , n1467 );
xor ( n1469 , n1466 , n1467 );
xor ( n1470 , n1331 , n1349 );
nor ( n1471 , n796 , n1447 );
and ( n1472 , n1470 , n1471 );
xor ( n1473 , n1470 , n1471 );
xor ( n1474 , n1335 , n1347 );
nor ( n1475 , n733 , n1447 );
and ( n1476 , n1474 , n1475 );
xor ( n1477 , n1474 , n1475 );
xor ( n1478 , n1340 , n1345 );
nor ( n1479 , n684 , n1447 );
and ( n1480 , n1478 , n1479 );
xor ( n1481 , n1478 , n1479 );
xor ( n1482 , n1342 , n1343 );
buf ( n1483 , n1482 );
nor ( n1484 , n646 , n1447 );
and ( n1485 , n1483 , n1484 );
xor ( n1486 , n1483 , n1484 );
nor ( n1487 , n601 , n1178 );
buf ( n1488 , n1487 );
nor ( n1489 , n622 , n1447 );
and ( n1490 , n1488 , n1489 );
buf ( n1491 , n1490 );
and ( n1492 , n1486 , n1491 );
or ( n1493 , n1485 , n1492 );
and ( n1494 , n1481 , n1493 );
or ( n1495 , n1480 , n1494 );
and ( n1496 , n1477 , n1495 );
or ( n1497 , n1476 , n1496 );
and ( n1498 , n1473 , n1497 );
or ( n1499 , n1472 , n1498 );
and ( n1500 , n1469 , n1499 );
or ( n1501 , n1468 , n1500 );
and ( n1502 , n1465 , n1501 );
or ( n1503 , n1464 , n1502 );
and ( n1504 , n1461 , n1503 );
or ( n1505 , n1460 , n1504 );
and ( n1506 , n1457 , n1505 );
or ( n1507 , n1456 , n1506 );
and ( n1508 , n1453 , n1507 );
or ( n1509 , n1452 , n1508 );
xor ( n1510 , n1449 , n1509 );
and ( n1511 , n1376 , n1377 );
and ( n1512 , n1377 , n1391 );
and ( n1513 , n1376 , n1391 );
or ( n1514 , n1511 , n1512 , n1513 );
and ( n1515 , n1372 , n1392 );
and ( n1516 , n1392 , n1431 );
and ( n1517 , n1372 , n1431 );
or ( n1518 , n1515 , n1516 , n1517 );
xor ( n1519 , n1514 , n1518 );
and ( n1520 , n1397 , n1412 );
and ( n1521 , n1412 , n1430 );
and ( n1522 , n1397 , n1430 );
or ( n1523 , n1520 , n1521 , n1522 );
and ( n1524 , n1417 , n1422 );
and ( n1525 , n1422 , n1429 );
and ( n1526 , n1417 , n1429 );
or ( n1527 , n1524 , n1525 , n1526 );
and ( n1528 , n1407 , n1408 );
and ( n1529 , n1408 , n1410 );
and ( n1530 , n1407 , n1410 );
or ( n1531 , n1528 , n1529 , n1530 );
and ( n1532 , n1418 , n1419 );
and ( n1533 , n1419 , n1421 );
and ( n1534 , n1418 , n1421 );
or ( n1535 , n1532 , n1533 , n1534 );
xor ( n1536 , n1531 , n1535 );
and ( n1537 , n925 , n719 );
buf ( n1538 , n1537 );
xor ( n1539 , n1536 , n1538 );
xor ( n1540 , n1527 , n1539 );
and ( n1541 , n1425 , n1426 );
and ( n1542 , n1426 , n1428 );
and ( n1543 , n1425 , n1428 );
or ( n1544 , n1541 , n1542 , n1543 );
and ( n1545 , n632 , n1134 );
and ( n1546 , n671 , n1034 );
xor ( n1547 , n1545 , n1546 );
and ( n1548 , n715 , n940 );
xor ( n1549 , n1547 , n1548 );
xor ( n1550 , n1544 , n1549 );
buf ( n1551 , n457 );
and ( n1552 , n599 , n1551 );
and ( n1553 , n608 , n1424 );
xor ( n1554 , n1552 , n1553 );
and ( n1555 , n611 , n1254 );
xor ( n1556 , n1554 , n1555 );
xor ( n1557 , n1550 , n1556 );
xor ( n1558 , n1540 , n1557 );
xor ( n1559 , n1523 , n1558 );
and ( n1560 , n1382 , n1384 );
and ( n1561 , n1384 , n1390 );
and ( n1562 , n1382 , n1390 );
or ( n1563 , n1560 , n1561 , n1562 );
and ( n1564 , n1401 , n1405 );
and ( n1565 , n1405 , n1411 );
and ( n1566 , n1401 , n1411 );
or ( n1567 , n1564 , n1565 , n1566 );
xor ( n1568 , n1563 , n1567 );
and ( n1569 , n1386 , n1387 );
and ( n1570 , n1387 , n1389 );
and ( n1571 , n1386 , n1389 );
or ( n1572 , n1569 , n1570 , n1571 );
and ( n1573 , n1047 , n663 );
and ( n1574 , n1164 , n635 );
xor ( n1575 , n1573 , n1574 );
and ( n1576 , n1287 , n606 );
xor ( n1577 , n1575 , n1576 );
xor ( n1578 , n1572 , n1577 );
and ( n1579 , n1383 , n615 );
buf ( n1580 , n457 );
and ( n1581 , n1580 , n612 );
xor ( n1582 , n1579 , n1581 );
xor ( n1583 , n1578 , n1582 );
xor ( n1584 , n1568 , n1583 );
xor ( n1585 , n1559 , n1584 );
xor ( n1586 , n1519 , n1585 );
and ( n1587 , n1363 , n1367 );
and ( n1588 , n1367 , n1432 );
and ( n1589 , n1363 , n1432 );
or ( n1590 , n1587 , n1588 , n1589 );
xor ( n1591 , n1586 , n1590 );
and ( n1592 , n1433 , n1437 );
and ( n1593 , n1438 , n1441 );
or ( n1594 , n1592 , n1593 );
xor ( n1595 , n1591 , n1594 );
buf ( n1596 , n1595 );
buf ( n1597 , n1596 );
not ( n1598 , n1597 );
buf ( n1599 , n511 );
not ( n1600 , n1599 );
nor ( n1601 , n1598 , n1600 );
xor ( n1602 , n1510 , n1601 );
xor ( n1603 , n1453 , n1507 );
nor ( n1604 , n1445 , n1600 );
and ( n1605 , n1603 , n1604 );
xor ( n1606 , n1603 , n1604 );
xor ( n1607 , n1457 , n1505 );
nor ( n1608 , n1303 , n1600 );
and ( n1609 , n1607 , n1608 );
xor ( n1610 , n1607 , n1608 );
xor ( n1611 , n1461 , n1503 );
nor ( n1612 , n1176 , n1600 );
and ( n1613 , n1611 , n1612 );
xor ( n1614 , n1611 , n1612 );
xor ( n1615 , n1465 , n1501 );
nor ( n1616 , n1062 , n1600 );
and ( n1617 , n1615 , n1616 );
xor ( n1618 , n1615 , n1616 );
xor ( n1619 , n1469 , n1499 );
nor ( n1620 , n958 , n1600 );
and ( n1621 , n1619 , n1620 );
xor ( n1622 , n1619 , n1620 );
xor ( n1623 , n1473 , n1497 );
nor ( n1624 , n868 , n1600 );
and ( n1625 , n1623 , n1624 );
xor ( n1626 , n1623 , n1624 );
xor ( n1627 , n1477 , n1495 );
nor ( n1628 , n796 , n1600 );
and ( n1629 , n1627 , n1628 );
xor ( n1630 , n1627 , n1628 );
xor ( n1631 , n1481 , n1493 );
nor ( n1632 , n733 , n1600 );
and ( n1633 , n1631 , n1632 );
xor ( n1634 , n1631 , n1632 );
xor ( n1635 , n1486 , n1491 );
nor ( n1636 , n684 , n1600 );
and ( n1637 , n1635 , n1636 );
xor ( n1638 , n1635 , n1636 );
xor ( n1639 , n1488 , n1489 );
buf ( n1640 , n1639 );
nor ( n1641 , n646 , n1600 );
and ( n1642 , n1640 , n1641 );
xor ( n1643 , n1640 , n1641 );
nor ( n1644 , n601 , n1305 );
buf ( n1645 , n1644 );
nor ( n1646 , n622 , n1600 );
and ( n1647 , n1645 , n1646 );
buf ( n1648 , n1647 );
and ( n1649 , n1643 , n1648 );
or ( n1650 , n1642 , n1649 );
and ( n1651 , n1638 , n1650 );
or ( n1652 , n1637 , n1651 );
and ( n1653 , n1634 , n1652 );
or ( n1654 , n1633 , n1653 );
and ( n1655 , n1630 , n1654 );
or ( n1656 , n1629 , n1655 );
and ( n1657 , n1626 , n1656 );
or ( n1658 , n1625 , n1657 );
and ( n1659 , n1622 , n1658 );
or ( n1660 , n1621 , n1659 );
and ( n1661 , n1618 , n1660 );
or ( n1662 , n1617 , n1661 );
and ( n1663 , n1614 , n1662 );
or ( n1664 , n1613 , n1663 );
and ( n1665 , n1610 , n1664 );
or ( n1666 , n1609 , n1665 );
and ( n1667 , n1606 , n1666 );
or ( n1668 , n1605 , n1667 );
xor ( n1669 , n1602 , n1668 );
and ( n1670 , n1523 , n1558 );
and ( n1671 , n1558 , n1584 );
and ( n1672 , n1523 , n1584 );
or ( n1673 , n1670 , n1671 , n1672 );
and ( n1674 , n1527 , n1539 );
and ( n1675 , n1539 , n1557 );
and ( n1676 , n1527 , n1557 );
or ( n1677 , n1674 , n1675 , n1676 );
and ( n1678 , n1531 , n1535 );
and ( n1679 , n1535 , n1538 );
and ( n1680 , n1531 , n1538 );
or ( n1681 , n1678 , n1679 , n1680 );
and ( n1682 , n1572 , n1577 );
and ( n1683 , n1577 , n1582 );
and ( n1684 , n1572 , n1582 );
or ( n1685 , n1682 , n1683 , n1684 );
xor ( n1686 , n1681 , n1685 );
and ( n1687 , n1573 , n1574 );
and ( n1688 , n1574 , n1576 );
and ( n1689 , n1573 , n1576 );
or ( n1690 , n1687 , n1688 , n1689 );
and ( n1691 , n1383 , n606 );
and ( n1692 , n1580 , n615 );
xor ( n1693 , n1691 , n1692 );
buf ( n1694 , n456 );
and ( n1695 , n1694 , n612 );
xor ( n1696 , n1693 , n1695 );
xor ( n1697 , n1690 , n1696 );
and ( n1698 , n1047 , n719 );
and ( n1699 , n1164 , n663 );
xor ( n1700 , n1698 , n1699 );
and ( n1701 , n1287 , n635 );
xor ( n1702 , n1700 , n1701 );
xor ( n1703 , n1697 , n1702 );
xor ( n1704 , n1686 , n1703 );
xor ( n1705 , n1677 , n1704 );
and ( n1706 , n1544 , n1549 );
and ( n1707 , n1549 , n1556 );
and ( n1708 , n1544 , n1556 );
or ( n1709 , n1706 , n1707 , n1708 );
and ( n1710 , n783 , n840 );
and ( n1711 , n856 , n771 );
and ( n1712 , n1710 , n1711 );
and ( n1713 , n1711 , n1537 );
and ( n1714 , n1710 , n1537 );
or ( n1715 , n1712 , n1713 , n1714 );
and ( n1716 , n1545 , n1546 );
and ( n1717 , n1546 , n1548 );
and ( n1718 , n1545 , n1548 );
or ( n1719 , n1716 , n1717 , n1718 );
xor ( n1720 , n1715 , n1719 );
and ( n1721 , n783 , n940 );
buf ( n1722 , n856 );
xor ( n1723 , n1721 , n1722 );
and ( n1724 , n925 , n771 );
xor ( n1725 , n1723 , n1724 );
xor ( n1726 , n1720 , n1725 );
xor ( n1727 , n1709 , n1726 );
and ( n1728 , n1552 , n1553 );
and ( n1729 , n1553 , n1555 );
and ( n1730 , n1552 , n1555 );
or ( n1731 , n1728 , n1729 , n1730 );
and ( n1732 , n632 , n1254 );
and ( n1733 , n671 , n1134 );
xor ( n1734 , n1732 , n1733 );
and ( n1735 , n715 , n1034 );
xor ( n1736 , n1734 , n1735 );
xor ( n1737 , n1731 , n1736 );
buf ( n1738 , n456 );
and ( n1739 , n599 , n1738 );
and ( n1740 , n608 , n1551 );
xor ( n1741 , n1739 , n1740 );
and ( n1742 , n611 , n1424 );
xor ( n1743 , n1741 , n1742 );
xor ( n1744 , n1737 , n1743 );
xor ( n1745 , n1727 , n1744 );
xor ( n1746 , n1705 , n1745 );
xor ( n1747 , n1673 , n1746 );
and ( n1748 , n1579 , n1581 );
and ( n1749 , n1563 , n1567 );
and ( n1750 , n1567 , n1583 );
and ( n1751 , n1563 , n1583 );
or ( n1752 , n1749 , n1750 , n1751 );
xor ( n1753 , n1748 , n1752 );
xor ( n1754 , n1747 , n1753 );
and ( n1755 , n1514 , n1518 );
and ( n1756 , n1518 , n1585 );
and ( n1757 , n1514 , n1585 );
or ( n1758 , n1755 , n1756 , n1757 );
xor ( n1759 , n1754 , n1758 );
and ( n1760 , n1586 , n1590 );
and ( n1761 , n1591 , n1594 );
or ( n1762 , n1760 , n1761 );
xor ( n1763 , n1759 , n1762 );
buf ( n1764 , n1763 );
buf ( n1765 , n1764 );
not ( n1766 , n1765 );
buf ( n1767 , n512 );
not ( n1768 , n1767 );
nor ( n1769 , n1766 , n1768 );
xor ( n1770 , n1669 , n1769 );
xor ( n1771 , n1606 , n1666 );
nor ( n1772 , n1598 , n1768 );
and ( n1773 , n1771 , n1772 );
xor ( n1774 , n1771 , n1772 );
xor ( n1775 , n1610 , n1664 );
nor ( n1776 , n1445 , n1768 );
and ( n1777 , n1775 , n1776 );
xor ( n1778 , n1775 , n1776 );
xor ( n1779 , n1614 , n1662 );
nor ( n1780 , n1303 , n1768 );
and ( n1781 , n1779 , n1780 );
xor ( n1782 , n1779 , n1780 );
xor ( n1783 , n1618 , n1660 );
nor ( n1784 , n1176 , n1768 );
and ( n1785 , n1783 , n1784 );
xor ( n1786 , n1783 , n1784 );
xor ( n1787 , n1622 , n1658 );
nor ( n1788 , n1062 , n1768 );
and ( n1789 , n1787 , n1788 );
xor ( n1790 , n1787 , n1788 );
xor ( n1791 , n1626 , n1656 );
nor ( n1792 , n958 , n1768 );
and ( n1793 , n1791 , n1792 );
xor ( n1794 , n1791 , n1792 );
xor ( n1795 , n1630 , n1654 );
nor ( n1796 , n868 , n1768 );
and ( n1797 , n1795 , n1796 );
xor ( n1798 , n1795 , n1796 );
xor ( n1799 , n1634 , n1652 );
nor ( n1800 , n796 , n1768 );
and ( n1801 , n1799 , n1800 );
xor ( n1802 , n1799 , n1800 );
xor ( n1803 , n1638 , n1650 );
nor ( n1804 , n733 , n1768 );
and ( n1805 , n1803 , n1804 );
xor ( n1806 , n1803 , n1804 );
xor ( n1807 , n1643 , n1648 );
nor ( n1808 , n684 , n1768 );
and ( n1809 , n1807 , n1808 );
xor ( n1810 , n1807 , n1808 );
xor ( n1811 , n1645 , n1646 );
buf ( n1812 , n1811 );
nor ( n1813 , n646 , n1768 );
and ( n1814 , n1812 , n1813 );
xor ( n1815 , n1812 , n1813 );
nor ( n1816 , n601 , n1447 );
buf ( n1817 , n1816 );
nor ( n1818 , n622 , n1768 );
and ( n1819 , n1817 , n1818 );
buf ( n1820 , n1819 );
and ( n1821 , n1815 , n1820 );
or ( n1822 , n1814 , n1821 );
and ( n1823 , n1810 , n1822 );
or ( n1824 , n1809 , n1823 );
and ( n1825 , n1806 , n1824 );
or ( n1826 , n1805 , n1825 );
and ( n1827 , n1802 , n1826 );
or ( n1828 , n1801 , n1827 );
and ( n1829 , n1798 , n1828 );
or ( n1830 , n1797 , n1829 );
and ( n1831 , n1794 , n1830 );
or ( n1832 , n1793 , n1831 );
and ( n1833 , n1790 , n1832 );
or ( n1834 , n1789 , n1833 );
and ( n1835 , n1786 , n1834 );
or ( n1836 , n1785 , n1835 );
and ( n1837 , n1782 , n1836 );
or ( n1838 , n1781 , n1837 );
and ( n1839 , n1778 , n1838 );
or ( n1840 , n1777 , n1839 );
and ( n1841 , n1774 , n1840 );
or ( n1842 , n1773 , n1841 );
xor ( n1843 , n1770 , n1842 );
and ( n1844 , n1748 , n1752 );
and ( n1845 , n1673 , n1746 );
and ( n1846 , n1746 , n1753 );
and ( n1847 , n1673 , n1753 );
or ( n1848 , n1845 , n1846 , n1847 );
xor ( n1849 , n1844 , n1848 );
and ( n1850 , n1677 , n1704 );
and ( n1851 , n1704 , n1745 );
and ( n1852 , n1677 , n1745 );
or ( n1853 , n1850 , n1851 , n1852 );
and ( n1854 , n1709 , n1726 );
and ( n1855 , n1726 , n1744 );
and ( n1856 , n1709 , n1744 );
or ( n1857 , n1854 , n1855 , n1856 );
and ( n1858 , n1731 , n1736 );
and ( n1859 , n1736 , n1743 );
and ( n1860 , n1731 , n1743 );
or ( n1861 , n1858 , n1859 , n1860 );
and ( n1862 , n1721 , n1722 );
and ( n1863 , n1722 , n1724 );
and ( n1864 , n1721 , n1724 );
or ( n1865 , n1862 , n1863 , n1864 );
and ( n1866 , n1732 , n1733 );
and ( n1867 , n1733 , n1735 );
and ( n1868 , n1732 , n1735 );
or ( n1869 , n1866 , n1867 , n1868 );
xor ( n1870 , n1865 , n1869 );
and ( n1871 , n783 , n1034 );
and ( n1872 , n856 , n940 );
xor ( n1873 , n1871 , n1872 );
and ( n1874 , n925 , n840 );
xor ( n1875 , n1873 , n1874 );
xor ( n1876 , n1870 , n1875 );
xor ( n1877 , n1861 , n1876 );
and ( n1878 , n1739 , n1740 );
and ( n1879 , n1740 , n1742 );
and ( n1880 , n1739 , n1742 );
or ( n1881 , n1878 , n1879 , n1880 );
buf ( n1882 , n455 );
and ( n1883 , n599 , n1882 );
and ( n1884 , n608 , n1738 );
xor ( n1885 , n1883 , n1884 );
and ( n1886 , n611 , n1551 );
xor ( n1887 , n1885 , n1886 );
xor ( n1888 , n1881 , n1887 );
and ( n1889 , n632 , n1424 );
and ( n1890 , n671 , n1254 );
xor ( n1891 , n1889 , n1890 );
and ( n1892 , n715 , n1134 );
xor ( n1893 , n1891 , n1892 );
xor ( n1894 , n1888 , n1893 );
xor ( n1895 , n1877 , n1894 );
xor ( n1896 , n1857 , n1895 );
and ( n1897 , n1690 , n1696 );
and ( n1898 , n1696 , n1702 );
and ( n1899 , n1690 , n1702 );
or ( n1900 , n1897 , n1898 , n1899 );
and ( n1901 , n1715 , n1719 );
and ( n1902 , n1719 , n1725 );
and ( n1903 , n1715 , n1725 );
or ( n1904 , n1901 , n1902 , n1903 );
xor ( n1905 , n1900 , n1904 );
and ( n1906 , n1698 , n1699 );
and ( n1907 , n1699 , n1701 );
and ( n1908 , n1698 , n1701 );
or ( n1909 , n1906 , n1907 , n1908 );
and ( n1910 , n1383 , n635 );
and ( n1911 , n1580 , n606 );
xor ( n1912 , n1910 , n1911 );
and ( n1913 , n1694 , n615 );
xor ( n1914 , n1912 , n1913 );
xor ( n1915 , n1909 , n1914 );
and ( n1916 , n1047 , n771 );
and ( n1917 , n1164 , n719 );
xor ( n1918 , n1916 , n1917 );
and ( n1919 , n1287 , n663 );
xor ( n1920 , n1918 , n1919 );
xor ( n1921 , n1915 , n1920 );
xor ( n1922 , n1905 , n1921 );
xor ( n1923 , n1896 , n1922 );
xor ( n1924 , n1853 , n1923 );
and ( n1925 , n1681 , n1685 );
and ( n1926 , n1685 , n1703 );
and ( n1927 , n1681 , n1703 );
or ( n1928 , n1925 , n1926 , n1927 );
and ( n1929 , n1691 , n1692 );
and ( n1930 , n1692 , n1695 );
and ( n1931 , n1691 , n1695 );
or ( n1932 , n1929 , n1930 , n1931 );
buf ( n1933 , n455 );
and ( n1934 , n1933 , n612 );
xor ( n1935 , n1932 , n1934 );
xor ( n1936 , n1928 , n1935 );
xor ( n1937 , n1924 , n1936 );
xor ( n1938 , n1849 , n1937 );
and ( n1939 , n1754 , n1758 );
and ( n1940 , n1759 , n1762 );
or ( n1941 , n1939 , n1940 );
xor ( n1942 , n1938 , n1941 );
buf ( n1943 , n1942 );
buf ( n1944 , n1943 );
not ( n1945 , n1944 );
buf ( n1946 , n513 );
not ( n1947 , n1946 );
nor ( n1948 , n1945 , n1947 );
xor ( n1949 , n1843 , n1948 );
xor ( n1950 , n1774 , n1840 );
nor ( n1951 , n1766 , n1947 );
and ( n1952 , n1950 , n1951 );
xor ( n1953 , n1950 , n1951 );
xor ( n1954 , n1778 , n1838 );
nor ( n1955 , n1598 , n1947 );
and ( n1956 , n1954 , n1955 );
xor ( n1957 , n1954 , n1955 );
xor ( n1958 , n1782 , n1836 );
nor ( n1959 , n1445 , n1947 );
and ( n1960 , n1958 , n1959 );
xor ( n1961 , n1958 , n1959 );
xor ( n1962 , n1786 , n1834 );
nor ( n1963 , n1303 , n1947 );
and ( n1964 , n1962 , n1963 );
xor ( n1965 , n1962 , n1963 );
xor ( n1966 , n1790 , n1832 );
nor ( n1967 , n1176 , n1947 );
and ( n1968 , n1966 , n1967 );
xor ( n1969 , n1966 , n1967 );
xor ( n1970 , n1794 , n1830 );
nor ( n1971 , n1062 , n1947 );
and ( n1972 , n1970 , n1971 );
xor ( n1973 , n1970 , n1971 );
xor ( n1974 , n1798 , n1828 );
nor ( n1975 , n958 , n1947 );
and ( n1976 , n1974 , n1975 );
xor ( n1977 , n1974 , n1975 );
xor ( n1978 , n1802 , n1826 );
nor ( n1979 , n868 , n1947 );
and ( n1980 , n1978 , n1979 );
xor ( n1981 , n1978 , n1979 );
xor ( n1982 , n1806 , n1824 );
nor ( n1983 , n796 , n1947 );
and ( n1984 , n1982 , n1983 );
xor ( n1985 , n1982 , n1983 );
xor ( n1986 , n1810 , n1822 );
nor ( n1987 , n733 , n1947 );
and ( n1988 , n1986 , n1987 );
xor ( n1989 , n1986 , n1987 );
xor ( n1990 , n1815 , n1820 );
nor ( n1991 , n684 , n1947 );
and ( n1992 , n1990 , n1991 );
xor ( n1993 , n1990 , n1991 );
xor ( n1994 , n1817 , n1818 );
buf ( n1995 , n1994 );
nor ( n1996 , n646 , n1947 );
and ( n1997 , n1995 , n1996 );
xor ( n1998 , n1995 , n1996 );
nor ( n1999 , n601 , n1600 );
buf ( n2000 , n1999 );
nor ( n2001 , n622 , n1947 );
and ( n2002 , n2000 , n2001 );
buf ( n2003 , n2002 );
and ( n2004 , n1998 , n2003 );
or ( n2005 , n1997 , n2004 );
and ( n2006 , n1993 , n2005 );
or ( n2007 , n1992 , n2006 );
and ( n2008 , n1989 , n2007 );
or ( n2009 , n1988 , n2008 );
and ( n2010 , n1985 , n2009 );
or ( n2011 , n1984 , n2010 );
and ( n2012 , n1981 , n2011 );
or ( n2013 , n1980 , n2012 );
and ( n2014 , n1977 , n2013 );
or ( n2015 , n1976 , n2014 );
and ( n2016 , n1973 , n2015 );
or ( n2017 , n1972 , n2016 );
and ( n2018 , n1969 , n2017 );
or ( n2019 , n1968 , n2018 );
and ( n2020 , n1965 , n2019 );
or ( n2021 , n1964 , n2020 );
and ( n2022 , n1961 , n2021 );
or ( n2023 , n1960 , n2022 );
and ( n2024 , n1957 , n2023 );
or ( n2025 , n1956 , n2024 );
and ( n2026 , n1953 , n2025 );
or ( n2027 , n1952 , n2026 );
xor ( n2028 , n1949 , n2027 );
and ( n2029 , n1928 , n1935 );
and ( n2030 , n1853 , n1923 );
and ( n2031 , n1923 , n1936 );
and ( n2032 , n1853 , n1936 );
or ( n2033 , n2030 , n2031 , n2032 );
xor ( n2034 , n2029 , n2033 );
and ( n2035 , n1857 , n1895 );
and ( n2036 , n1895 , n1922 );
and ( n2037 , n1857 , n1922 );
or ( n2038 , n2035 , n2036 , n2037 );
and ( n2039 , n1861 , n1876 );
and ( n2040 , n1876 , n1894 );
and ( n2041 , n1861 , n1894 );
or ( n2042 , n2039 , n2040 , n2041 );
and ( n2043 , n1865 , n1869 );
and ( n2044 , n1869 , n1875 );
and ( n2045 , n1865 , n1875 );
or ( n2046 , n2043 , n2044 , n2045 );
and ( n2047 , n1909 , n1914 );
and ( n2048 , n1914 , n1920 );
and ( n2049 , n1909 , n1920 );
or ( n2050 , n2047 , n2048 , n2049 );
xor ( n2051 , n2046 , n2050 );
and ( n2052 , n1916 , n1917 );
and ( n2053 , n1917 , n1919 );
and ( n2054 , n1916 , n1919 );
or ( n2055 , n2052 , n2053 , n2054 );
and ( n2056 , n1383 , n663 );
and ( n2057 , n1580 , n635 );
xor ( n2058 , n2056 , n2057 );
and ( n2059 , n1694 , n606 );
xor ( n2060 , n2058 , n2059 );
xor ( n2061 , n2055 , n2060 );
and ( n2062 , n1047 , n840 );
and ( n2063 , n1164 , n771 );
xor ( n2064 , n2062 , n2063 );
and ( n2065 , n1287 , n719 );
xor ( n2066 , n2064 , n2065 );
xor ( n2067 , n2061 , n2066 );
xor ( n2068 , n2051 , n2067 );
xor ( n2069 , n2042 , n2068 );
and ( n2070 , n1881 , n1887 );
and ( n2071 , n1887 , n1893 );
and ( n2072 , n1881 , n1893 );
or ( n2073 , n2070 , n2071 , n2072 );
and ( n2074 , n1871 , n1872 );
and ( n2075 , n1872 , n1874 );
and ( n2076 , n1871 , n1874 );
or ( n2077 , n2074 , n2075 , n2076 );
and ( n2078 , n1889 , n1890 );
and ( n2079 , n1890 , n1892 );
and ( n2080 , n1889 , n1892 );
or ( n2081 , n2078 , n2079 , n2080 );
xor ( n2082 , n2077 , n2081 );
and ( n2083 , n783 , n1134 );
and ( n2084 , n856 , n1034 );
xor ( n2085 , n2083 , n2084 );
buf ( n2086 , n925 );
xor ( n2087 , n2085 , n2086 );
xor ( n2088 , n2082 , n2087 );
xor ( n2089 , n2073 , n2088 );
and ( n2090 , n1883 , n1884 );
and ( n2091 , n1884 , n1886 );
and ( n2092 , n1883 , n1886 );
or ( n2093 , n2090 , n2091 , n2092 );
and ( n2094 , n632 , n1551 );
and ( n2095 , n671 , n1424 );
xor ( n2096 , n2094 , n2095 );
and ( n2097 , n715 , n1254 );
xor ( n2098 , n2096 , n2097 );
xor ( n2099 , n2093 , n2098 );
buf ( n2100 , n454 );
and ( n2101 , n599 , n2100 );
and ( n2102 , n608 , n1882 );
xor ( n2103 , n2101 , n2102 );
and ( n2104 , n611 , n1738 );
xor ( n2105 , n2103 , n2104 );
xor ( n2106 , n2099 , n2105 );
xor ( n2107 , n2089 , n2106 );
xor ( n2108 , n2069 , n2107 );
xor ( n2109 , n2038 , n2108 );
and ( n2110 , n1900 , n1904 );
and ( n2111 , n1904 , n1921 );
and ( n2112 , n1900 , n1921 );
or ( n2113 , n2110 , n2111 , n2112 );
and ( n2114 , n1932 , n1934 );
and ( n2115 , n1910 , n1911 );
and ( n2116 , n1911 , n1913 );
and ( n2117 , n1910 , n1913 );
or ( n2118 , n2115 , n2116 , n2117 );
and ( n2119 , n1933 , n615 );
buf ( n2120 , n454 );
and ( n2121 , n2120 , n612 );
xor ( n2122 , n2119 , n2121 );
xor ( n2123 , n2118 , n2122 );
xor ( n2124 , n2114 , n2123 );
xor ( n2125 , n2113 , n2124 );
xor ( n2126 , n2109 , n2125 );
xor ( n2127 , n2034 , n2126 );
and ( n2128 , n1844 , n1848 );
and ( n2129 , n1848 , n1937 );
and ( n2130 , n1844 , n1937 );
or ( n2131 , n2128 , n2129 , n2130 );
xor ( n2132 , n2127 , n2131 );
and ( n2133 , n1938 , n1941 );
xor ( n2134 , n2132 , n2133 );
buf ( n2135 , n2134 );
buf ( n2136 , n2135 );
not ( n2137 , n2136 );
buf ( n2138 , n514 );
not ( n2139 , n2138 );
nor ( n2140 , n2137 , n2139 );
xor ( n2141 , n2028 , n2140 );
xor ( n2142 , n1953 , n2025 );
nor ( n2143 , n1945 , n2139 );
and ( n2144 , n2142 , n2143 );
xor ( n2145 , n2142 , n2143 );
xor ( n2146 , n1957 , n2023 );
nor ( n2147 , n1766 , n2139 );
and ( n2148 , n2146 , n2147 );
xor ( n2149 , n2146 , n2147 );
xor ( n2150 , n1961 , n2021 );
nor ( n2151 , n1598 , n2139 );
and ( n2152 , n2150 , n2151 );
xor ( n2153 , n2150 , n2151 );
xor ( n2154 , n1965 , n2019 );
nor ( n2155 , n1445 , n2139 );
and ( n2156 , n2154 , n2155 );
xor ( n2157 , n2154 , n2155 );
xor ( n2158 , n1969 , n2017 );
nor ( n2159 , n1303 , n2139 );
and ( n2160 , n2158 , n2159 );
xor ( n2161 , n2158 , n2159 );
xor ( n2162 , n1973 , n2015 );
nor ( n2163 , n1176 , n2139 );
and ( n2164 , n2162 , n2163 );
xor ( n2165 , n2162 , n2163 );
xor ( n2166 , n1977 , n2013 );
nor ( n2167 , n1062 , n2139 );
and ( n2168 , n2166 , n2167 );
xor ( n2169 , n2166 , n2167 );
xor ( n2170 , n1981 , n2011 );
nor ( n2171 , n958 , n2139 );
and ( n2172 , n2170 , n2171 );
xor ( n2173 , n2170 , n2171 );
xor ( n2174 , n1985 , n2009 );
nor ( n2175 , n868 , n2139 );
and ( n2176 , n2174 , n2175 );
xor ( n2177 , n2174 , n2175 );
xor ( n2178 , n1989 , n2007 );
nor ( n2179 , n796 , n2139 );
and ( n2180 , n2178 , n2179 );
xor ( n2181 , n2178 , n2179 );
xor ( n2182 , n1993 , n2005 );
nor ( n2183 , n733 , n2139 );
and ( n2184 , n2182 , n2183 );
xor ( n2185 , n2182 , n2183 );
xor ( n2186 , n1998 , n2003 );
nor ( n2187 , n684 , n2139 );
and ( n2188 , n2186 , n2187 );
xor ( n2189 , n2186 , n2187 );
xor ( n2190 , n2000 , n2001 );
buf ( n2191 , n2190 );
nor ( n2192 , n646 , n2139 );
and ( n2193 , n2191 , n2192 );
xor ( n2194 , n2191 , n2192 );
nor ( n2195 , n601 , n1768 );
buf ( n2196 , n2195 );
nor ( n2197 , n622 , n2139 );
and ( n2198 , n2196 , n2197 );
buf ( n2199 , n2198 );
and ( n2200 , n2194 , n2199 );
or ( n2201 , n2193 , n2200 );
and ( n2202 , n2189 , n2201 );
or ( n2203 , n2188 , n2202 );
and ( n2204 , n2185 , n2203 );
or ( n2205 , n2184 , n2204 );
and ( n2206 , n2181 , n2205 );
or ( n2207 , n2180 , n2206 );
and ( n2208 , n2177 , n2207 );
or ( n2209 , n2176 , n2208 );
and ( n2210 , n2173 , n2209 );
or ( n2211 , n2172 , n2210 );
and ( n2212 , n2169 , n2211 );
or ( n2213 , n2168 , n2212 );
and ( n2214 , n2165 , n2213 );
or ( n2215 , n2164 , n2214 );
and ( n2216 , n2161 , n2215 );
or ( n2217 , n2160 , n2216 );
and ( n2218 , n2157 , n2217 );
or ( n2219 , n2156 , n2218 );
and ( n2220 , n2153 , n2219 );
or ( n2221 , n2152 , n2220 );
and ( n2222 , n2149 , n2221 );
or ( n2223 , n2148 , n2222 );
and ( n2224 , n2145 , n2223 );
or ( n2225 , n2144 , n2224 );
xor ( n2226 , n2141 , n2225 );
and ( n2227 , n2113 , n2124 );
and ( n2228 , n2038 , n2108 );
and ( n2229 , n2108 , n2125 );
and ( n2230 , n2038 , n2125 );
or ( n2231 , n2228 , n2229 , n2230 );
xor ( n2232 , n2227 , n2231 );
and ( n2233 , n2042 , n2068 );
and ( n2234 , n2068 , n2107 );
and ( n2235 , n2042 , n2107 );
or ( n2236 , n2233 , n2234 , n2235 );
and ( n2237 , n2073 , n2088 );
and ( n2238 , n2088 , n2106 );
and ( n2239 , n2073 , n2106 );
or ( n2240 , n2237 , n2238 , n2239 );
and ( n2241 , n2055 , n2060 );
and ( n2242 , n2060 , n2066 );
and ( n2243 , n2055 , n2066 );
or ( n2244 , n2241 , n2242 , n2243 );
and ( n2245 , n2077 , n2081 );
and ( n2246 , n2081 , n2087 );
and ( n2247 , n2077 , n2087 );
or ( n2248 , n2245 , n2246 , n2247 );
xor ( n2249 , n2244 , n2248 );
and ( n2250 , n2062 , n2063 );
and ( n2251 , n2063 , n2065 );
and ( n2252 , n2062 , n2065 );
or ( n2253 , n2250 , n2251 , n2252 );
and ( n2254 , n1383 , n719 );
and ( n2255 , n1580 , n663 );
xor ( n2256 , n2254 , n2255 );
and ( n2257 , n1694 , n635 );
xor ( n2258 , n2256 , n2257 );
xor ( n2259 , n2253 , n2258 );
and ( n2260 , n1047 , n940 );
and ( n2261 , n1164 , n840 );
xor ( n2262 , n2260 , n2261 );
and ( n2263 , n1287 , n771 );
xor ( n2264 , n2262 , n2263 );
xor ( n2265 , n2259 , n2264 );
xor ( n2266 , n2249 , n2265 );
xor ( n2267 , n2240 , n2266 );
and ( n2268 , n2093 , n2098 );
and ( n2269 , n2098 , n2105 );
and ( n2270 , n2093 , n2105 );
or ( n2271 , n2268 , n2269 , n2270 );
and ( n2272 , n2094 , n2095 );
and ( n2273 , n2095 , n2097 );
and ( n2274 , n2094 , n2097 );
or ( n2275 , n2272 , n2273 , n2274 );
and ( n2276 , n2083 , n2084 );
and ( n2277 , n2084 , n2086 );
and ( n2278 , n2083 , n2086 );
or ( n2279 , n2276 , n2277 , n2278 );
xor ( n2280 , n2275 , n2279 );
and ( n2281 , n783 , n1254 );
and ( n2282 , n856 , n1134 );
xor ( n2283 , n2281 , n2282 );
and ( n2284 , n925 , n1034 );
xor ( n2285 , n2283 , n2284 );
xor ( n2286 , n2280 , n2285 );
xor ( n2287 , n2271 , n2286 );
and ( n2288 , n2101 , n2102 );
and ( n2289 , n2102 , n2104 );
and ( n2290 , n2101 , n2104 );
or ( n2291 , n2288 , n2289 , n2290 );
and ( n2292 , n632 , n1738 );
and ( n2293 , n671 , n1551 );
xor ( n2294 , n2292 , n2293 );
and ( n2295 , n715 , n1424 );
xor ( n2296 , n2294 , n2295 );
xor ( n2297 , n2291 , n2296 );
buf ( n2298 , n453 );
and ( n2299 , n599 , n2298 );
and ( n2300 , n608 , n2100 );
xor ( n2301 , n2299 , n2300 );
and ( n2302 , n611 , n1882 );
xor ( n2303 , n2301 , n2302 );
xor ( n2304 , n2297 , n2303 );
xor ( n2305 , n2287 , n2304 );
xor ( n2306 , n2267 , n2305 );
xor ( n2307 , n2236 , n2306 );
and ( n2308 , n2046 , n2050 );
and ( n2309 , n2050 , n2067 );
and ( n2310 , n2046 , n2067 );
or ( n2311 , n2308 , n2309 , n2310 );
and ( n2312 , n2114 , n2123 );
xor ( n2313 , n2311 , n2312 );
and ( n2314 , n2118 , n2122 );
and ( n2315 , n2056 , n2057 );
and ( n2316 , n2057 , n2059 );
and ( n2317 , n2056 , n2059 );
or ( n2318 , n2315 , n2316 , n2317 );
and ( n2319 , n2119 , n2121 );
xor ( n2320 , n2318 , n2319 );
and ( n2321 , n1933 , n606 );
and ( n2322 , n2120 , n615 );
xor ( n2323 , n2321 , n2322 );
buf ( n2324 , n453 );
and ( n2325 , n2324 , n612 );
xor ( n2326 , n2323 , n2325 );
xor ( n2327 , n2320 , n2326 );
xor ( n2328 , n2314 , n2327 );
xor ( n2329 , n2313 , n2328 );
xor ( n2330 , n2307 , n2329 );
xor ( n2331 , n2232 , n2330 );
and ( n2332 , n2029 , n2033 );
and ( n2333 , n2033 , n2126 );
and ( n2334 , n2029 , n2126 );
or ( n2335 , n2332 , n2333 , n2334 );
xor ( n2336 , n2331 , n2335 );
and ( n2337 , n2127 , n2131 );
and ( n2338 , n2132 , n2133 );
or ( n2339 , n2337 , n2338 );
xor ( n2340 , n2336 , n2339 );
buf ( n2341 , n2340 );
buf ( n2342 , n2341 );
not ( n2343 , n2342 );
buf ( n2344 , n515 );
not ( n2345 , n2344 );
nor ( n2346 , n2343 , n2345 );
xor ( n2347 , n2226 , n2346 );
xor ( n2348 , n2145 , n2223 );
nor ( n2349 , n2137 , n2345 );
and ( n2350 , n2348 , n2349 );
xor ( n2351 , n2348 , n2349 );
xor ( n2352 , n2149 , n2221 );
nor ( n2353 , n1945 , n2345 );
and ( n2354 , n2352 , n2353 );
xor ( n2355 , n2352 , n2353 );
xor ( n2356 , n2153 , n2219 );
nor ( n2357 , n1766 , n2345 );
and ( n2358 , n2356 , n2357 );
xor ( n2359 , n2356 , n2357 );
xor ( n2360 , n2157 , n2217 );
nor ( n2361 , n1598 , n2345 );
and ( n2362 , n2360 , n2361 );
xor ( n2363 , n2360 , n2361 );
xor ( n2364 , n2161 , n2215 );
nor ( n2365 , n1445 , n2345 );
and ( n2366 , n2364 , n2365 );
xor ( n2367 , n2364 , n2365 );
xor ( n2368 , n2165 , n2213 );
nor ( n2369 , n1303 , n2345 );
and ( n2370 , n2368 , n2369 );
xor ( n2371 , n2368 , n2369 );
xor ( n2372 , n2169 , n2211 );
nor ( n2373 , n1176 , n2345 );
and ( n2374 , n2372 , n2373 );
xor ( n2375 , n2372 , n2373 );
xor ( n2376 , n2173 , n2209 );
nor ( n2377 , n1062 , n2345 );
and ( n2378 , n2376 , n2377 );
xor ( n2379 , n2376 , n2377 );
xor ( n2380 , n2177 , n2207 );
nor ( n2381 , n958 , n2345 );
and ( n2382 , n2380 , n2381 );
xor ( n2383 , n2380 , n2381 );
xor ( n2384 , n2181 , n2205 );
nor ( n2385 , n868 , n2345 );
and ( n2386 , n2384 , n2385 );
xor ( n2387 , n2384 , n2385 );
xor ( n2388 , n2185 , n2203 );
nor ( n2389 , n796 , n2345 );
and ( n2390 , n2388 , n2389 );
xor ( n2391 , n2388 , n2389 );
xor ( n2392 , n2189 , n2201 );
nor ( n2393 , n733 , n2345 );
and ( n2394 , n2392 , n2393 );
xor ( n2395 , n2392 , n2393 );
xor ( n2396 , n2194 , n2199 );
nor ( n2397 , n684 , n2345 );
and ( n2398 , n2396 , n2397 );
xor ( n2399 , n2396 , n2397 );
xor ( n2400 , n2196 , n2197 );
buf ( n2401 , n2400 );
nor ( n2402 , n646 , n2345 );
and ( n2403 , n2401 , n2402 );
xor ( n2404 , n2401 , n2402 );
nor ( n2405 , n601 , n1947 );
buf ( n2406 , n2405 );
nor ( n2407 , n622 , n2345 );
and ( n2408 , n2406 , n2407 );
buf ( n2409 , n2408 );
and ( n2410 , n2404 , n2409 );
or ( n2411 , n2403 , n2410 );
and ( n2412 , n2399 , n2411 );
or ( n2413 , n2398 , n2412 );
and ( n2414 , n2395 , n2413 );
or ( n2415 , n2394 , n2414 );
and ( n2416 , n2391 , n2415 );
or ( n2417 , n2390 , n2416 );
and ( n2418 , n2387 , n2417 );
or ( n2419 , n2386 , n2418 );
and ( n2420 , n2383 , n2419 );
or ( n2421 , n2382 , n2420 );
and ( n2422 , n2379 , n2421 );
or ( n2423 , n2378 , n2422 );
and ( n2424 , n2375 , n2423 );
or ( n2425 , n2374 , n2424 );
and ( n2426 , n2371 , n2425 );
or ( n2427 , n2370 , n2426 );
and ( n2428 , n2367 , n2427 );
or ( n2429 , n2366 , n2428 );
and ( n2430 , n2363 , n2429 );
or ( n2431 , n2362 , n2430 );
and ( n2432 , n2359 , n2431 );
or ( n2433 , n2358 , n2432 );
and ( n2434 , n2355 , n2433 );
or ( n2435 , n2354 , n2434 );
and ( n2436 , n2351 , n2435 );
or ( n2437 , n2350 , n2436 );
xor ( n2438 , n2347 , n2437 );
and ( n2439 , n2311 , n2312 );
and ( n2440 , n2312 , n2328 );
and ( n2441 , n2311 , n2328 );
or ( n2442 , n2439 , n2440 , n2441 );
and ( n2443 , n2236 , n2306 );
and ( n2444 , n2306 , n2329 );
and ( n2445 , n2236 , n2329 );
or ( n2446 , n2443 , n2444 , n2445 );
xor ( n2447 , n2442 , n2446 );
and ( n2448 , n2240 , n2266 );
and ( n2449 , n2266 , n2305 );
and ( n2450 , n2240 , n2305 );
or ( n2451 , n2448 , n2449 , n2450 );
and ( n2452 , n2244 , n2248 );
and ( n2453 , n2248 , n2265 );
and ( n2454 , n2244 , n2265 );
or ( n2455 , n2452 , n2453 , n2454 );
and ( n2456 , n2314 , n2327 );
xor ( n2457 , n2455 , n2456 );
and ( n2458 , n2318 , n2319 );
and ( n2459 , n2319 , n2326 );
and ( n2460 , n2318 , n2326 );
or ( n2461 , n2458 , n2459 , n2460 );
buf ( n2462 , n452 );
and ( n2463 , n2462 , n612 );
xor ( n2464 , n2461 , n2463 );
and ( n2465 , n2321 , n2322 );
and ( n2466 , n2322 , n2325 );
and ( n2467 , n2321 , n2325 );
or ( n2468 , n2465 , n2466 , n2467 );
and ( n2469 , n2254 , n2255 );
and ( n2470 , n2255 , n2257 );
and ( n2471 , n2254 , n2257 );
or ( n2472 , n2469 , n2470 , n2471 );
xor ( n2473 , n2468 , n2472 );
and ( n2474 , n1933 , n635 );
and ( n2475 , n2120 , n606 );
xor ( n2476 , n2474 , n2475 );
and ( n2477 , n2324 , n615 );
xor ( n2478 , n2476 , n2477 );
xor ( n2479 , n2473 , n2478 );
xor ( n2480 , n2464 , n2479 );
xor ( n2481 , n2457 , n2480 );
xor ( n2482 , n2451 , n2481 );
and ( n2483 , n2271 , n2286 );
and ( n2484 , n2286 , n2304 );
and ( n2485 , n2271 , n2304 );
or ( n2486 , n2483 , n2484 , n2485 );
and ( n2487 , n2253 , n2258 );
and ( n2488 , n2258 , n2264 );
and ( n2489 , n2253 , n2264 );
or ( n2490 , n2487 , n2488 , n2489 );
and ( n2491 , n2275 , n2279 );
and ( n2492 , n2279 , n2285 );
and ( n2493 , n2275 , n2285 );
or ( n2494 , n2491 , n2492 , n2493 );
xor ( n2495 , n2490 , n2494 );
and ( n2496 , n2260 , n2261 );
and ( n2497 , n2261 , n2263 );
and ( n2498 , n2260 , n2263 );
or ( n2499 , n2496 , n2497 , n2498 );
and ( n2500 , n1383 , n771 );
and ( n2501 , n1580 , n719 );
xor ( n2502 , n2500 , n2501 );
and ( n2503 , n1694 , n663 );
xor ( n2504 , n2502 , n2503 );
xor ( n2505 , n2499 , n2504 );
buf ( n2506 , n1047 );
and ( n2507 , n1164 , n940 );
xor ( n2508 , n2506 , n2507 );
and ( n2509 , n1287 , n840 );
xor ( n2510 , n2508 , n2509 );
xor ( n2511 , n2505 , n2510 );
xor ( n2512 , n2495 , n2511 );
xor ( n2513 , n2486 , n2512 );
and ( n2514 , n2291 , n2296 );
and ( n2515 , n2296 , n2303 );
and ( n2516 , n2291 , n2303 );
or ( n2517 , n2514 , n2515 , n2516 );
and ( n2518 , n2281 , n2282 );
and ( n2519 , n2282 , n2284 );
and ( n2520 , n2281 , n2284 );
or ( n2521 , n2518 , n2519 , n2520 );
and ( n2522 , n2292 , n2293 );
and ( n2523 , n2293 , n2295 );
and ( n2524 , n2292 , n2295 );
or ( n2525 , n2522 , n2523 , n2524 );
xor ( n2526 , n2521 , n2525 );
and ( n2527 , n783 , n1424 );
and ( n2528 , n856 , n1254 );
xor ( n2529 , n2527 , n2528 );
and ( n2530 , n925 , n1134 );
xor ( n2531 , n2529 , n2530 );
xor ( n2532 , n2526 , n2531 );
xor ( n2533 , n2517 , n2532 );
and ( n2534 , n2299 , n2300 );
and ( n2535 , n2300 , n2302 );
and ( n2536 , n2299 , n2302 );
or ( n2537 , n2534 , n2535 , n2536 );
and ( n2538 , n632 , n1882 );
and ( n2539 , n671 , n1738 );
xor ( n2540 , n2538 , n2539 );
and ( n2541 , n715 , n1551 );
xor ( n2542 , n2540 , n2541 );
xor ( n2543 , n2537 , n2542 );
buf ( n2544 , n452 );
and ( n2545 , n599 , n2544 );
and ( n2546 , n608 , n2298 );
xor ( n2547 , n2545 , n2546 );
and ( n2548 , n611 , n2100 );
xor ( n2549 , n2547 , n2548 );
xor ( n2550 , n2543 , n2549 );
xor ( n2551 , n2533 , n2550 );
xor ( n2552 , n2513 , n2551 );
xor ( n2553 , n2482 , n2552 );
xor ( n2554 , n2447 , n2553 );
and ( n2555 , n2227 , n2231 );
and ( n2556 , n2231 , n2330 );
and ( n2557 , n2227 , n2330 );
or ( n2558 , n2555 , n2556 , n2557 );
xor ( n2559 , n2554 , n2558 );
and ( n2560 , n2331 , n2335 );
and ( n2561 , n2336 , n2339 );
or ( n2562 , n2560 , n2561 );
xor ( n2563 , n2559 , n2562 );
buf ( n2564 , n2563 );
buf ( n2565 , n2564 );
not ( n2566 , n2565 );
buf ( n2567 , n516 );
not ( n2568 , n2567 );
nor ( n2569 , n2566 , n2568 );
xor ( n2570 , n2438 , n2569 );
xor ( n2571 , n2351 , n2435 );
nor ( n2572 , n2343 , n2568 );
and ( n2573 , n2571 , n2572 );
xor ( n2574 , n2571 , n2572 );
xor ( n2575 , n2355 , n2433 );
nor ( n2576 , n2137 , n2568 );
and ( n2577 , n2575 , n2576 );
xor ( n2578 , n2575 , n2576 );
xor ( n2579 , n2359 , n2431 );
nor ( n2580 , n1945 , n2568 );
and ( n2581 , n2579 , n2580 );
xor ( n2582 , n2579 , n2580 );
xor ( n2583 , n2363 , n2429 );
nor ( n2584 , n1766 , n2568 );
and ( n2585 , n2583 , n2584 );
xor ( n2586 , n2583 , n2584 );
xor ( n2587 , n2367 , n2427 );
nor ( n2588 , n1598 , n2568 );
and ( n2589 , n2587 , n2588 );
xor ( n2590 , n2587 , n2588 );
xor ( n2591 , n2371 , n2425 );
nor ( n2592 , n1445 , n2568 );
and ( n2593 , n2591 , n2592 );
xor ( n2594 , n2591 , n2592 );
xor ( n2595 , n2375 , n2423 );
nor ( n2596 , n1303 , n2568 );
and ( n2597 , n2595 , n2596 );
xor ( n2598 , n2595 , n2596 );
xor ( n2599 , n2379 , n2421 );
nor ( n2600 , n1176 , n2568 );
and ( n2601 , n2599 , n2600 );
xor ( n2602 , n2599 , n2600 );
xor ( n2603 , n2383 , n2419 );
nor ( n2604 , n1062 , n2568 );
and ( n2605 , n2603 , n2604 );
xor ( n2606 , n2603 , n2604 );
xor ( n2607 , n2387 , n2417 );
nor ( n2608 , n958 , n2568 );
and ( n2609 , n2607 , n2608 );
xor ( n2610 , n2607 , n2608 );
xor ( n2611 , n2391 , n2415 );
nor ( n2612 , n868 , n2568 );
and ( n2613 , n2611 , n2612 );
xor ( n2614 , n2611 , n2612 );
xor ( n2615 , n2395 , n2413 );
nor ( n2616 , n796 , n2568 );
and ( n2617 , n2615 , n2616 );
xor ( n2618 , n2615 , n2616 );
xor ( n2619 , n2399 , n2411 );
nor ( n2620 , n733 , n2568 );
and ( n2621 , n2619 , n2620 );
xor ( n2622 , n2619 , n2620 );
xor ( n2623 , n2404 , n2409 );
nor ( n2624 , n684 , n2568 );
and ( n2625 , n2623 , n2624 );
xor ( n2626 , n2623 , n2624 );
xor ( n2627 , n2406 , n2407 );
buf ( n2628 , n2627 );
nor ( n2629 , n646 , n2568 );
and ( n2630 , n2628 , n2629 );
xor ( n2631 , n2628 , n2629 );
nor ( n2632 , n601 , n2139 );
buf ( n2633 , n2632 );
nor ( n2634 , n622 , n2568 );
and ( n2635 , n2633 , n2634 );
buf ( n2636 , n2635 );
and ( n2637 , n2631 , n2636 );
or ( n2638 , n2630 , n2637 );
and ( n2639 , n2626 , n2638 );
or ( n2640 , n2625 , n2639 );
and ( n2641 , n2622 , n2640 );
or ( n2642 , n2621 , n2641 );
and ( n2643 , n2618 , n2642 );
or ( n2644 , n2617 , n2643 );
and ( n2645 , n2614 , n2644 );
or ( n2646 , n2613 , n2645 );
and ( n2647 , n2610 , n2646 );
or ( n2648 , n2609 , n2647 );
and ( n2649 , n2606 , n2648 );
or ( n2650 , n2605 , n2649 );
and ( n2651 , n2602 , n2650 );
or ( n2652 , n2601 , n2651 );
and ( n2653 , n2598 , n2652 );
or ( n2654 , n2597 , n2653 );
and ( n2655 , n2594 , n2654 );
or ( n2656 , n2593 , n2655 );
and ( n2657 , n2590 , n2656 );
or ( n2658 , n2589 , n2657 );
and ( n2659 , n2586 , n2658 );
or ( n2660 , n2585 , n2659 );
and ( n2661 , n2582 , n2660 );
or ( n2662 , n2581 , n2661 );
and ( n2663 , n2578 , n2662 );
or ( n2664 , n2577 , n2663 );
and ( n2665 , n2574 , n2664 );
or ( n2666 , n2573 , n2665 );
xor ( n2667 , n2570 , n2666 );
and ( n2668 , n2455 , n2456 );
and ( n2669 , n2456 , n2480 );
and ( n2670 , n2455 , n2480 );
or ( n2671 , n2668 , n2669 , n2670 );
and ( n2672 , n2451 , n2481 );
and ( n2673 , n2481 , n2552 );
and ( n2674 , n2451 , n2552 );
or ( n2675 , n2672 , n2673 , n2674 );
xor ( n2676 , n2671 , n2675 );
and ( n2677 , n2486 , n2512 );
and ( n2678 , n2512 , n2551 );
and ( n2679 , n2486 , n2551 );
or ( n2680 , n2677 , n2678 , n2679 );
and ( n2681 , n2517 , n2532 );
and ( n2682 , n2532 , n2550 );
and ( n2683 , n2517 , n2550 );
or ( n2684 , n2681 , n2682 , n2683 );
and ( n2685 , n2499 , n2504 );
and ( n2686 , n2504 , n2510 );
and ( n2687 , n2499 , n2510 );
or ( n2688 , n2685 , n2686 , n2687 );
and ( n2689 , n2521 , n2525 );
and ( n2690 , n2525 , n2531 );
and ( n2691 , n2521 , n2531 );
or ( n2692 , n2689 , n2690 , n2691 );
xor ( n2693 , n2688 , n2692 );
and ( n2694 , n2506 , n2507 );
and ( n2695 , n2507 , n2509 );
and ( n2696 , n2506 , n2509 );
or ( n2697 , n2694 , n2695 , n2696 );
and ( n2698 , n1383 , n840 );
and ( n2699 , n1580 , n771 );
xor ( n2700 , n2698 , n2699 );
and ( n2701 , n1694 , n719 );
xor ( n2702 , n2700 , n2701 );
xor ( n2703 , n2697 , n2702 );
and ( n2704 , n1287 , n940 );
buf ( n2705 , n2704 );
xor ( n2706 , n2703 , n2705 );
xor ( n2707 , n2693 , n2706 );
xor ( n2708 , n2684 , n2707 );
and ( n2709 , n2537 , n2542 );
and ( n2710 , n2542 , n2549 );
and ( n2711 , n2537 , n2549 );
or ( n2712 , n2709 , n2710 , n2711 );
and ( n2713 , n2527 , n2528 );
and ( n2714 , n2528 , n2530 );
and ( n2715 , n2527 , n2530 );
or ( n2716 , n2713 , n2714 , n2715 );
and ( n2717 , n2538 , n2539 );
and ( n2718 , n2539 , n2541 );
and ( n2719 , n2538 , n2541 );
or ( n2720 , n2717 , n2718 , n2719 );
xor ( n2721 , n2716 , n2720 );
and ( n2722 , n783 , n1551 );
and ( n2723 , n856 , n1424 );
xor ( n2724 , n2722 , n2723 );
and ( n2725 , n925 , n1254 );
xor ( n2726 , n2724 , n2725 );
xor ( n2727 , n2721 , n2726 );
xor ( n2728 , n2712 , n2727 );
and ( n2729 , n2545 , n2546 );
and ( n2730 , n2546 , n2548 );
and ( n2731 , n2545 , n2548 );
or ( n2732 , n2729 , n2730 , n2731 );
and ( n2733 , n632 , n2100 );
and ( n2734 , n671 , n1882 );
xor ( n2735 , n2733 , n2734 );
and ( n2736 , n715 , n1738 );
xor ( n2737 , n2735 , n2736 );
xor ( n2738 , n2732 , n2737 );
buf ( n2739 , n451 );
and ( n2740 , n599 , n2739 );
and ( n2741 , n608 , n2544 );
xor ( n2742 , n2740 , n2741 );
and ( n2743 , n611 , n2298 );
xor ( n2744 , n2742 , n2743 );
xor ( n2745 , n2738 , n2744 );
xor ( n2746 , n2728 , n2745 );
xor ( n2747 , n2708 , n2746 );
xor ( n2748 , n2680 , n2747 );
and ( n2749 , n2461 , n2463 );
and ( n2750 , n2463 , n2479 );
and ( n2751 , n2461 , n2479 );
or ( n2752 , n2749 , n2750 , n2751 );
and ( n2753 , n2490 , n2494 );
and ( n2754 , n2494 , n2511 );
and ( n2755 , n2490 , n2511 );
or ( n2756 , n2753 , n2754 , n2755 );
xor ( n2757 , n2752 , n2756 );
and ( n2758 , n2468 , n2472 );
and ( n2759 , n2472 , n2478 );
and ( n2760 , n2468 , n2478 );
or ( n2761 , n2758 , n2759 , n2760 );
and ( n2762 , n2474 , n2475 );
and ( n2763 , n2475 , n2477 );
and ( n2764 , n2474 , n2477 );
or ( n2765 , n2762 , n2763 , n2764 );
and ( n2766 , n2500 , n2501 );
and ( n2767 , n2501 , n2503 );
and ( n2768 , n2500 , n2503 );
or ( n2769 , n2766 , n2767 , n2768 );
xor ( n2770 , n2765 , n2769 );
and ( n2771 , n1933 , n663 );
and ( n2772 , n2120 , n635 );
xor ( n2773 , n2771 , n2772 );
and ( n2774 , n2324 , n606 );
xor ( n2775 , n2773 , n2774 );
xor ( n2776 , n2770 , n2775 );
xor ( n2777 , n2761 , n2776 );
and ( n2778 , n2462 , n615 );
buf ( n2779 , n451 );
and ( n2780 , n2779 , n612 );
xor ( n2781 , n2778 , n2780 );
xor ( n2782 , n2777 , n2781 );
xor ( n2783 , n2757 , n2782 );
xor ( n2784 , n2748 , n2783 );
xor ( n2785 , n2676 , n2784 );
and ( n2786 , n2442 , n2446 );
and ( n2787 , n2446 , n2553 );
and ( n2788 , n2442 , n2553 );
or ( n2789 , n2786 , n2787 , n2788 );
xor ( n2790 , n2785 , n2789 );
and ( n2791 , n2554 , n2558 );
and ( n2792 , n2559 , n2562 );
or ( n2793 , n2791 , n2792 );
xor ( n2794 , n2790 , n2793 );
buf ( n2795 , n2794 );
buf ( n2796 , n2795 );
not ( n2797 , n2796 );
buf ( n2798 , n517 );
not ( n2799 , n2798 );
nor ( n2800 , n2797 , n2799 );
xor ( n2801 , n2667 , n2800 );
xor ( n2802 , n2574 , n2664 );
nor ( n2803 , n2566 , n2799 );
and ( n2804 , n2802 , n2803 );
xor ( n2805 , n2802 , n2803 );
xor ( n2806 , n2578 , n2662 );
nor ( n2807 , n2343 , n2799 );
and ( n2808 , n2806 , n2807 );
xor ( n2809 , n2806 , n2807 );
xor ( n2810 , n2582 , n2660 );
nor ( n2811 , n2137 , n2799 );
and ( n2812 , n2810 , n2811 );
xor ( n2813 , n2810 , n2811 );
xor ( n2814 , n2586 , n2658 );
nor ( n2815 , n1945 , n2799 );
and ( n2816 , n2814 , n2815 );
xor ( n2817 , n2814 , n2815 );
xor ( n2818 , n2590 , n2656 );
nor ( n2819 , n1766 , n2799 );
and ( n2820 , n2818 , n2819 );
xor ( n2821 , n2818 , n2819 );
xor ( n2822 , n2594 , n2654 );
nor ( n2823 , n1598 , n2799 );
and ( n2824 , n2822 , n2823 );
xor ( n2825 , n2822 , n2823 );
xor ( n2826 , n2598 , n2652 );
nor ( n2827 , n1445 , n2799 );
and ( n2828 , n2826 , n2827 );
xor ( n2829 , n2826 , n2827 );
xor ( n2830 , n2602 , n2650 );
nor ( n2831 , n1303 , n2799 );
and ( n2832 , n2830 , n2831 );
xor ( n2833 , n2830 , n2831 );
xor ( n2834 , n2606 , n2648 );
nor ( n2835 , n1176 , n2799 );
and ( n2836 , n2834 , n2835 );
xor ( n2837 , n2834 , n2835 );
xor ( n2838 , n2610 , n2646 );
nor ( n2839 , n1062 , n2799 );
and ( n2840 , n2838 , n2839 );
xor ( n2841 , n2838 , n2839 );
xor ( n2842 , n2614 , n2644 );
nor ( n2843 , n958 , n2799 );
and ( n2844 , n2842 , n2843 );
xor ( n2845 , n2842 , n2843 );
xor ( n2846 , n2618 , n2642 );
nor ( n2847 , n868 , n2799 );
and ( n2848 , n2846 , n2847 );
xor ( n2849 , n2846 , n2847 );
xor ( n2850 , n2622 , n2640 );
nor ( n2851 , n796 , n2799 );
and ( n2852 , n2850 , n2851 );
xor ( n2853 , n2850 , n2851 );
xor ( n2854 , n2626 , n2638 );
nor ( n2855 , n733 , n2799 );
and ( n2856 , n2854 , n2855 );
xor ( n2857 , n2854 , n2855 );
xor ( n2858 , n2631 , n2636 );
nor ( n2859 , n684 , n2799 );
and ( n2860 , n2858 , n2859 );
xor ( n2861 , n2858 , n2859 );
xor ( n2862 , n2633 , n2634 );
buf ( n2863 , n2862 );
nor ( n2864 , n646 , n2799 );
and ( n2865 , n2863 , n2864 );
xor ( n2866 , n2863 , n2864 );
nor ( n2867 , n601 , n2345 );
buf ( n2868 , n2867 );
nor ( n2869 , n622 , n2799 );
and ( n2870 , n2868 , n2869 );
buf ( n2871 , n2870 );
and ( n2872 , n2866 , n2871 );
or ( n2873 , n2865 , n2872 );
and ( n2874 , n2861 , n2873 );
or ( n2875 , n2860 , n2874 );
and ( n2876 , n2857 , n2875 );
or ( n2877 , n2856 , n2876 );
and ( n2878 , n2853 , n2877 );
or ( n2879 , n2852 , n2878 );
and ( n2880 , n2849 , n2879 );
or ( n2881 , n2848 , n2880 );
and ( n2882 , n2845 , n2881 );
or ( n2883 , n2844 , n2882 );
and ( n2884 , n2841 , n2883 );
or ( n2885 , n2840 , n2884 );
and ( n2886 , n2837 , n2885 );
or ( n2887 , n2836 , n2886 );
and ( n2888 , n2833 , n2887 );
or ( n2889 , n2832 , n2888 );
and ( n2890 , n2829 , n2889 );
or ( n2891 , n2828 , n2890 );
and ( n2892 , n2825 , n2891 );
or ( n2893 , n2824 , n2892 );
and ( n2894 , n2821 , n2893 );
or ( n2895 , n2820 , n2894 );
and ( n2896 , n2817 , n2895 );
or ( n2897 , n2816 , n2896 );
and ( n2898 , n2813 , n2897 );
or ( n2899 , n2812 , n2898 );
and ( n2900 , n2809 , n2899 );
or ( n2901 , n2808 , n2900 );
and ( n2902 , n2805 , n2901 );
or ( n2903 , n2804 , n2902 );
xor ( n2904 , n2801 , n2903 );
and ( n2905 , n2752 , n2756 );
and ( n2906 , n2756 , n2782 );
and ( n2907 , n2752 , n2782 );
or ( n2908 , n2905 , n2906 , n2907 );
and ( n2909 , n2680 , n2747 );
and ( n2910 , n2747 , n2783 );
and ( n2911 , n2680 , n2783 );
or ( n2912 , n2909 , n2910 , n2911 );
xor ( n2913 , n2908 , n2912 );
and ( n2914 , n2684 , n2707 );
and ( n2915 , n2707 , n2746 );
and ( n2916 , n2684 , n2746 );
or ( n2917 , n2914 , n2915 , n2916 );
and ( n2918 , n2712 , n2727 );
and ( n2919 , n2727 , n2745 );
and ( n2920 , n2712 , n2745 );
or ( n2921 , n2918 , n2919 , n2920 );
and ( n2922 , n2697 , n2702 );
and ( n2923 , n2702 , n2705 );
and ( n2924 , n2697 , n2705 );
or ( n2925 , n2922 , n2923 , n2924 );
and ( n2926 , n2716 , n2720 );
and ( n2927 , n2720 , n2726 );
and ( n2928 , n2716 , n2726 );
or ( n2929 , n2926 , n2927 , n2928 );
xor ( n2930 , n2925 , n2929 );
and ( n2931 , n1047 , n1134 );
and ( n2932 , n1164 , n1034 );
and ( n2933 , n2931 , n2932 );
and ( n2934 , n2932 , n2704 );
and ( n2935 , n2931 , n2704 );
or ( n2936 , n2933 , n2934 , n2935 );
and ( n2937 , n1383 , n940 );
and ( n2938 , n1580 , n840 );
xor ( n2939 , n2937 , n2938 );
and ( n2940 , n1694 , n771 );
xor ( n2941 , n2939 , n2940 );
xor ( n2942 , n2936 , n2941 );
and ( n2943 , n1047 , n1254 );
buf ( n2944 , n1164 );
xor ( n2945 , n2943 , n2944 );
and ( n2946 , n1287 , n1034 );
xor ( n2947 , n2945 , n2946 );
xor ( n2948 , n2942 , n2947 );
xor ( n2949 , n2930 , n2948 );
xor ( n2950 , n2921 , n2949 );
and ( n2951 , n2732 , n2737 );
and ( n2952 , n2737 , n2744 );
and ( n2953 , n2732 , n2744 );
or ( n2954 , n2951 , n2952 , n2953 );
and ( n2955 , n2722 , n2723 );
and ( n2956 , n2723 , n2725 );
and ( n2957 , n2722 , n2725 );
or ( n2958 , n2955 , n2956 , n2957 );
and ( n2959 , n2733 , n2734 );
and ( n2960 , n2734 , n2736 );
and ( n2961 , n2733 , n2736 );
or ( n2962 , n2959 , n2960 , n2961 );
xor ( n2963 , n2958 , n2962 );
and ( n2964 , n783 , n1738 );
and ( n2965 , n856 , n1551 );
xor ( n2966 , n2964 , n2965 );
and ( n2967 , n925 , n1424 );
xor ( n2968 , n2966 , n2967 );
xor ( n2969 , n2963 , n2968 );
xor ( n2970 , n2954 , n2969 );
and ( n2971 , n2740 , n2741 );
and ( n2972 , n2741 , n2743 );
and ( n2973 , n2740 , n2743 );
or ( n2974 , n2971 , n2972 , n2973 );
and ( n2975 , n632 , n2298 );
and ( n2976 , n671 , n2100 );
xor ( n2977 , n2975 , n2976 );
and ( n2978 , n715 , n1882 );
xor ( n2979 , n2977 , n2978 );
xor ( n2980 , n2974 , n2979 );
buf ( n2981 , n450 );
and ( n2982 , n599 , n2981 );
and ( n2983 , n608 , n2739 );
xor ( n2984 , n2982 , n2983 );
and ( n2985 , n611 , n2544 );
xor ( n2986 , n2984 , n2985 );
xor ( n2987 , n2980 , n2986 );
xor ( n2988 , n2970 , n2987 );
xor ( n2989 , n2950 , n2988 );
xor ( n2990 , n2917 , n2989 );
and ( n2991 , n2688 , n2692 );
and ( n2992 , n2692 , n2706 );
and ( n2993 , n2688 , n2706 );
or ( n2994 , n2991 , n2992 , n2993 );
and ( n2995 , n2761 , n2776 );
and ( n2996 , n2776 , n2781 );
and ( n2997 , n2761 , n2781 );
or ( n2998 , n2995 , n2996 , n2997 );
xor ( n2999 , n2994 , n2998 );
and ( n3000 , n2765 , n2769 );
and ( n3001 , n2769 , n2775 );
and ( n3002 , n2765 , n2775 );
or ( n3003 , n3000 , n3001 , n3002 );
and ( n3004 , n2771 , n2772 );
and ( n3005 , n2772 , n2774 );
and ( n3006 , n2771 , n2774 );
or ( n3007 , n3004 , n3005 , n3006 );
and ( n3008 , n2698 , n2699 );
and ( n3009 , n2699 , n2701 );
and ( n3010 , n2698 , n2701 );
or ( n3011 , n3008 , n3009 , n3010 );
xor ( n3012 , n3007 , n3011 );
and ( n3013 , n1933 , n719 );
and ( n3014 , n2120 , n663 );
xor ( n3015 , n3013 , n3014 );
and ( n3016 , n2324 , n635 );
xor ( n3017 , n3015 , n3016 );
xor ( n3018 , n3012 , n3017 );
xor ( n3019 , n3003 , n3018 );
and ( n3020 , n2778 , n2780 );
and ( n3021 , n2462 , n606 );
and ( n3022 , n2779 , n615 );
xor ( n3023 , n3021 , n3022 );
buf ( n3024 , n450 );
and ( n3025 , n3024 , n612 );
xor ( n3026 , n3023 , n3025 );
xor ( n3027 , n3020 , n3026 );
xor ( n3028 , n3019 , n3027 );
xor ( n3029 , n2999 , n3028 );
xor ( n3030 , n2990 , n3029 );
xor ( n3031 , n2913 , n3030 );
and ( n3032 , n2671 , n2675 );
and ( n3033 , n2675 , n2784 );
and ( n3034 , n2671 , n2784 );
or ( n3035 , n3032 , n3033 , n3034 );
xor ( n3036 , n3031 , n3035 );
and ( n3037 , n2785 , n2789 );
and ( n3038 , n2790 , n2793 );
or ( n3039 , n3037 , n3038 );
xor ( n3040 , n3036 , n3039 );
buf ( n3041 , n3040 );
buf ( n3042 , n3041 );
not ( n3043 , n3042 );
buf ( n3044 , n518 );
not ( n3045 , n3044 );
nor ( n3046 , n3043 , n3045 );
xor ( n3047 , n2904 , n3046 );
xor ( n3048 , n2805 , n2901 );
nor ( n3049 , n2797 , n3045 );
and ( n3050 , n3048 , n3049 );
xor ( n3051 , n3048 , n3049 );
xor ( n3052 , n2809 , n2899 );
nor ( n3053 , n2566 , n3045 );
and ( n3054 , n3052 , n3053 );
xor ( n3055 , n3052 , n3053 );
xor ( n3056 , n2813 , n2897 );
nor ( n3057 , n2343 , n3045 );
and ( n3058 , n3056 , n3057 );
xor ( n3059 , n3056 , n3057 );
xor ( n3060 , n2817 , n2895 );
nor ( n3061 , n2137 , n3045 );
and ( n3062 , n3060 , n3061 );
xor ( n3063 , n3060 , n3061 );
xor ( n3064 , n2821 , n2893 );
nor ( n3065 , n1945 , n3045 );
and ( n3066 , n3064 , n3065 );
xor ( n3067 , n3064 , n3065 );
xor ( n3068 , n2825 , n2891 );
nor ( n3069 , n1766 , n3045 );
and ( n3070 , n3068 , n3069 );
xor ( n3071 , n3068 , n3069 );
xor ( n3072 , n2829 , n2889 );
nor ( n3073 , n1598 , n3045 );
and ( n3074 , n3072 , n3073 );
xor ( n3075 , n3072 , n3073 );
xor ( n3076 , n2833 , n2887 );
nor ( n3077 , n1445 , n3045 );
and ( n3078 , n3076 , n3077 );
xor ( n3079 , n3076 , n3077 );
xor ( n3080 , n2837 , n2885 );
nor ( n3081 , n1303 , n3045 );
and ( n3082 , n3080 , n3081 );
xor ( n3083 , n3080 , n3081 );
xor ( n3084 , n2841 , n2883 );
nor ( n3085 , n1176 , n3045 );
and ( n3086 , n3084 , n3085 );
xor ( n3087 , n3084 , n3085 );
xor ( n3088 , n2845 , n2881 );
nor ( n3089 , n1062 , n3045 );
and ( n3090 , n3088 , n3089 );
xor ( n3091 , n3088 , n3089 );
xor ( n3092 , n2849 , n2879 );
nor ( n3093 , n958 , n3045 );
and ( n3094 , n3092 , n3093 );
xor ( n3095 , n3092 , n3093 );
xor ( n3096 , n2853 , n2877 );
nor ( n3097 , n868 , n3045 );
and ( n3098 , n3096 , n3097 );
xor ( n3099 , n3096 , n3097 );
xor ( n3100 , n2857 , n2875 );
nor ( n3101 , n796 , n3045 );
and ( n3102 , n3100 , n3101 );
xor ( n3103 , n3100 , n3101 );
xor ( n3104 , n2861 , n2873 );
nor ( n3105 , n733 , n3045 );
and ( n3106 , n3104 , n3105 );
xor ( n3107 , n3104 , n3105 );
xor ( n3108 , n2866 , n2871 );
nor ( n3109 , n684 , n3045 );
and ( n3110 , n3108 , n3109 );
xor ( n3111 , n3108 , n3109 );
xor ( n3112 , n2868 , n2869 );
buf ( n3113 , n3112 );
nor ( n3114 , n646 , n3045 );
and ( n3115 , n3113 , n3114 );
xor ( n3116 , n3113 , n3114 );
nor ( n3117 , n601 , n2568 );
buf ( n3118 , n3117 );
nor ( n3119 , n622 , n3045 );
and ( n3120 , n3118 , n3119 );
buf ( n3121 , n3120 );
and ( n3122 , n3116 , n3121 );
or ( n3123 , n3115 , n3122 );
and ( n3124 , n3111 , n3123 );
or ( n3125 , n3110 , n3124 );
and ( n3126 , n3107 , n3125 );
or ( n3127 , n3106 , n3126 );
and ( n3128 , n3103 , n3127 );
or ( n3129 , n3102 , n3128 );
and ( n3130 , n3099 , n3129 );
or ( n3131 , n3098 , n3130 );
and ( n3132 , n3095 , n3131 );
or ( n3133 , n3094 , n3132 );
and ( n3134 , n3091 , n3133 );
or ( n3135 , n3090 , n3134 );
and ( n3136 , n3087 , n3135 );
or ( n3137 , n3086 , n3136 );
and ( n3138 , n3083 , n3137 );
or ( n3139 , n3082 , n3138 );
and ( n3140 , n3079 , n3139 );
or ( n3141 , n3078 , n3140 );
and ( n3142 , n3075 , n3141 );
or ( n3143 , n3074 , n3142 );
and ( n3144 , n3071 , n3143 );
or ( n3145 , n3070 , n3144 );
and ( n3146 , n3067 , n3145 );
or ( n3147 , n3066 , n3146 );
and ( n3148 , n3063 , n3147 );
or ( n3149 , n3062 , n3148 );
and ( n3150 , n3059 , n3149 );
or ( n3151 , n3058 , n3150 );
and ( n3152 , n3055 , n3151 );
or ( n3153 , n3054 , n3152 );
and ( n3154 , n3051 , n3153 );
or ( n3155 , n3050 , n3154 );
xor ( n3156 , n3047 , n3155 );
and ( n3157 , n2917 , n2989 );
and ( n3158 , n2989 , n3029 );
and ( n3159 , n2917 , n3029 );
or ( n3160 , n3157 , n3158 , n3159 );
and ( n3161 , n2921 , n2949 );
and ( n3162 , n2949 , n2988 );
and ( n3163 , n2921 , n2988 );
or ( n3164 , n3161 , n3162 , n3163 );
and ( n3165 , n2925 , n2929 );
and ( n3166 , n2929 , n2948 );
and ( n3167 , n2925 , n2948 );
or ( n3168 , n3165 , n3166 , n3167 );
and ( n3169 , n3003 , n3018 );
and ( n3170 , n3018 , n3027 );
and ( n3171 , n3003 , n3027 );
or ( n3172 , n3169 , n3170 , n3171 );
xor ( n3173 , n3168 , n3172 );
and ( n3174 , n3007 , n3011 );
and ( n3175 , n3011 , n3017 );
and ( n3176 , n3007 , n3017 );
or ( n3177 , n3174 , n3175 , n3176 );
and ( n3178 , n3021 , n3022 );
and ( n3179 , n3022 , n3025 );
and ( n3180 , n3021 , n3025 );
or ( n3181 , n3178 , n3179 , n3180 );
buf ( n3182 , n449 );
and ( n3183 , n3182 , n612 );
xor ( n3184 , n3181 , n3183 );
and ( n3185 , n2462 , n635 );
and ( n3186 , n2779 , n606 );
xor ( n3187 , n3185 , n3186 );
and ( n3188 , n3024 , n615 );
xor ( n3189 , n3187 , n3188 );
xor ( n3190 , n3184 , n3189 );
xor ( n3191 , n3177 , n3190 );
and ( n3192 , n3013 , n3014 );
and ( n3193 , n3014 , n3016 );
and ( n3194 , n3013 , n3016 );
or ( n3195 , n3192 , n3193 , n3194 );
and ( n3196 , n2937 , n2938 );
and ( n3197 , n2938 , n2940 );
and ( n3198 , n2937 , n2940 );
or ( n3199 , n3196 , n3197 , n3198 );
xor ( n3200 , n3195 , n3199 );
and ( n3201 , n1933 , n771 );
and ( n3202 , n2120 , n719 );
xor ( n3203 , n3201 , n3202 );
and ( n3204 , n2324 , n663 );
xor ( n3205 , n3203 , n3204 );
xor ( n3206 , n3200 , n3205 );
xor ( n3207 , n3191 , n3206 );
xor ( n3208 , n3173 , n3207 );
xor ( n3209 , n3164 , n3208 );
and ( n3210 , n2954 , n2969 );
and ( n3211 , n2969 , n2987 );
and ( n3212 , n2954 , n2987 );
or ( n3213 , n3210 , n3211 , n3212 );
and ( n3214 , n2936 , n2941 );
and ( n3215 , n2941 , n2947 );
and ( n3216 , n2936 , n2947 );
or ( n3217 , n3214 , n3215 , n3216 );
and ( n3218 , n2958 , n2962 );
and ( n3219 , n2962 , n2968 );
and ( n3220 , n2958 , n2968 );
or ( n3221 , n3218 , n3219 , n3220 );
xor ( n3222 , n3217 , n3221 );
and ( n3223 , n2943 , n2944 );
and ( n3224 , n2944 , n2946 );
and ( n3225 , n2943 , n2946 );
or ( n3226 , n3223 , n3224 , n3225 );
and ( n3227 , n1383 , n1034 );
and ( n3228 , n1580 , n940 );
xor ( n3229 , n3227 , n3228 );
and ( n3230 , n1694 , n840 );
xor ( n3231 , n3229 , n3230 );
xor ( n3232 , n3226 , n3231 );
and ( n3233 , n1047 , n1424 );
and ( n3234 , n1164 , n1254 );
xor ( n3235 , n3233 , n3234 );
and ( n3236 , n1287 , n1134 );
xor ( n3237 , n3235 , n3236 );
xor ( n3238 , n3232 , n3237 );
xor ( n3239 , n3222 , n3238 );
xor ( n3240 , n3213 , n3239 );
and ( n3241 , n2974 , n2979 );
and ( n3242 , n2979 , n2986 );
and ( n3243 , n2974 , n2986 );
or ( n3244 , n3241 , n3242 , n3243 );
and ( n3245 , n2964 , n2965 );
and ( n3246 , n2965 , n2967 );
and ( n3247 , n2964 , n2967 );
or ( n3248 , n3245 , n3246 , n3247 );
and ( n3249 , n2975 , n2976 );
and ( n3250 , n2976 , n2978 );
and ( n3251 , n2975 , n2978 );
or ( n3252 , n3249 , n3250 , n3251 );
xor ( n3253 , n3248 , n3252 );
and ( n3254 , n783 , n1882 );
and ( n3255 , n856 , n1738 );
xor ( n3256 , n3254 , n3255 );
and ( n3257 , n925 , n1551 );
xor ( n3258 , n3256 , n3257 );
xor ( n3259 , n3253 , n3258 );
xor ( n3260 , n3244 , n3259 );
and ( n3261 , n2982 , n2983 );
and ( n3262 , n2983 , n2985 );
and ( n3263 , n2982 , n2985 );
or ( n3264 , n3261 , n3262 , n3263 );
and ( n3265 , n632 , n2544 );
and ( n3266 , n671 , n2298 );
xor ( n3267 , n3265 , n3266 );
and ( n3268 , n715 , n2100 );
xor ( n3269 , n3267 , n3268 );
xor ( n3270 , n3264 , n3269 );
buf ( n3271 , n449 );
and ( n3272 , n599 , n3271 );
and ( n3273 , n608 , n2981 );
xor ( n3274 , n3272 , n3273 );
and ( n3275 , n611 , n2739 );
xor ( n3276 , n3274 , n3275 );
xor ( n3277 , n3270 , n3276 );
xor ( n3278 , n3260 , n3277 );
xor ( n3279 , n3240 , n3278 );
xor ( n3280 , n3209 , n3279 );
xor ( n3281 , n3160 , n3280 );
and ( n3282 , n3020 , n3026 );
and ( n3283 , n2994 , n2998 );
and ( n3284 , n2998 , n3028 );
and ( n3285 , n2994 , n3028 );
or ( n3286 , n3283 , n3284 , n3285 );
xor ( n3287 , n3282 , n3286 );
xor ( n3288 , n3281 , n3287 );
and ( n3289 , n2908 , n2912 );
and ( n3290 , n2912 , n3030 );
and ( n3291 , n2908 , n3030 );
or ( n3292 , n3289 , n3290 , n3291 );
xor ( n3293 , n3288 , n3292 );
and ( n3294 , n3031 , n3035 );
and ( n3295 , n3036 , n3039 );
or ( n3296 , n3294 , n3295 );
xor ( n3297 , n3293 , n3296 );
buf ( n3298 , n3297 );
buf ( n3299 , n3298 );
not ( n3300 , n3299 );
buf ( n3301 , n519 );
not ( n3302 , n3301 );
nor ( n3303 , n3300 , n3302 );
xor ( n3304 , n3156 , n3303 );
xor ( n3305 , n3051 , n3153 );
nor ( n3306 , n3043 , n3302 );
and ( n3307 , n3305 , n3306 );
xor ( n3308 , n3305 , n3306 );
xor ( n3309 , n3055 , n3151 );
nor ( n3310 , n2797 , n3302 );
and ( n3311 , n3309 , n3310 );
xor ( n3312 , n3309 , n3310 );
xor ( n3313 , n3059 , n3149 );
nor ( n3314 , n2566 , n3302 );
and ( n3315 , n3313 , n3314 );
xor ( n3316 , n3313 , n3314 );
xor ( n3317 , n3063 , n3147 );
nor ( n3318 , n2343 , n3302 );
and ( n3319 , n3317 , n3318 );
xor ( n3320 , n3317 , n3318 );
xor ( n3321 , n3067 , n3145 );
nor ( n3322 , n2137 , n3302 );
and ( n3323 , n3321 , n3322 );
xor ( n3324 , n3321 , n3322 );
xor ( n3325 , n3071 , n3143 );
nor ( n3326 , n1945 , n3302 );
and ( n3327 , n3325 , n3326 );
xor ( n3328 , n3325 , n3326 );
xor ( n3329 , n3075 , n3141 );
nor ( n3330 , n1766 , n3302 );
and ( n3331 , n3329 , n3330 );
xor ( n3332 , n3329 , n3330 );
xor ( n3333 , n3079 , n3139 );
nor ( n3334 , n1598 , n3302 );
and ( n3335 , n3333 , n3334 );
xor ( n3336 , n3333 , n3334 );
xor ( n3337 , n3083 , n3137 );
nor ( n3338 , n1445 , n3302 );
and ( n3339 , n3337 , n3338 );
xor ( n3340 , n3337 , n3338 );
xor ( n3341 , n3087 , n3135 );
nor ( n3342 , n1303 , n3302 );
and ( n3343 , n3341 , n3342 );
xor ( n3344 , n3341 , n3342 );
xor ( n3345 , n3091 , n3133 );
nor ( n3346 , n1176 , n3302 );
and ( n3347 , n3345 , n3346 );
xor ( n3348 , n3345 , n3346 );
xor ( n3349 , n3095 , n3131 );
nor ( n3350 , n1062 , n3302 );
and ( n3351 , n3349 , n3350 );
xor ( n3352 , n3349 , n3350 );
xor ( n3353 , n3099 , n3129 );
nor ( n3354 , n958 , n3302 );
and ( n3355 , n3353 , n3354 );
xor ( n3356 , n3353 , n3354 );
xor ( n3357 , n3103 , n3127 );
nor ( n3358 , n868 , n3302 );
and ( n3359 , n3357 , n3358 );
xor ( n3360 , n3357 , n3358 );
xor ( n3361 , n3107 , n3125 );
nor ( n3362 , n796 , n3302 );
and ( n3363 , n3361 , n3362 );
xor ( n3364 , n3361 , n3362 );
xor ( n3365 , n3111 , n3123 );
nor ( n3366 , n733 , n3302 );
and ( n3367 , n3365 , n3366 );
xor ( n3368 , n3365 , n3366 );
xor ( n3369 , n3116 , n3121 );
nor ( n3370 , n684 , n3302 );
and ( n3371 , n3369 , n3370 );
xor ( n3372 , n3369 , n3370 );
xor ( n3373 , n3118 , n3119 );
buf ( n3374 , n3373 );
nor ( n3375 , n646 , n3302 );
and ( n3376 , n3374 , n3375 );
xor ( n3377 , n3374 , n3375 );
nor ( n3378 , n601 , n2799 );
buf ( n3379 , n3378 );
nor ( n3380 , n622 , n3302 );
and ( n3381 , n3379 , n3380 );
buf ( n3382 , n3381 );
and ( n3383 , n3377 , n3382 );
or ( n3384 , n3376 , n3383 );
and ( n3385 , n3372 , n3384 );
or ( n3386 , n3371 , n3385 );
and ( n3387 , n3368 , n3386 );
or ( n3388 , n3367 , n3387 );
and ( n3389 , n3364 , n3388 );
or ( n3390 , n3363 , n3389 );
and ( n3391 , n3360 , n3390 );
or ( n3392 , n3359 , n3391 );
and ( n3393 , n3356 , n3392 );
or ( n3394 , n3355 , n3393 );
and ( n3395 , n3352 , n3394 );
or ( n3396 , n3351 , n3395 );
and ( n3397 , n3348 , n3396 );
or ( n3398 , n3347 , n3397 );
and ( n3399 , n3344 , n3398 );
or ( n3400 , n3343 , n3399 );
and ( n3401 , n3340 , n3400 );
or ( n3402 , n3339 , n3401 );
and ( n3403 , n3336 , n3402 );
or ( n3404 , n3335 , n3403 );
and ( n3405 , n3332 , n3404 );
or ( n3406 , n3331 , n3405 );
and ( n3407 , n3328 , n3406 );
or ( n3408 , n3327 , n3407 );
and ( n3409 , n3324 , n3408 );
or ( n3410 , n3323 , n3409 );
and ( n3411 , n3320 , n3410 );
or ( n3412 , n3319 , n3411 );
and ( n3413 , n3316 , n3412 );
or ( n3414 , n3315 , n3413 );
and ( n3415 , n3312 , n3414 );
or ( n3416 , n3311 , n3415 );
and ( n3417 , n3308 , n3416 );
or ( n3418 , n3307 , n3417 );
xor ( n3419 , n3304 , n3418 );
and ( n3420 , n3282 , n3286 );
and ( n3421 , n3160 , n3280 );
and ( n3422 , n3280 , n3287 );
and ( n3423 , n3160 , n3287 );
or ( n3424 , n3421 , n3422 , n3423 );
xor ( n3425 , n3420 , n3424 );
and ( n3426 , n3164 , n3208 );
and ( n3427 , n3208 , n3279 );
and ( n3428 , n3164 , n3279 );
or ( n3429 , n3426 , n3427 , n3428 );
and ( n3430 , n3213 , n3239 );
and ( n3431 , n3239 , n3278 );
and ( n3432 , n3213 , n3278 );
or ( n3433 , n3430 , n3431 , n3432 );
and ( n3434 , n3244 , n3259 );
and ( n3435 , n3259 , n3277 );
and ( n3436 , n3244 , n3277 );
or ( n3437 , n3434 , n3435 , n3436 );
and ( n3438 , n3226 , n3231 );
and ( n3439 , n3231 , n3237 );
and ( n3440 , n3226 , n3237 );
or ( n3441 , n3438 , n3439 , n3440 );
and ( n3442 , n3248 , n3252 );
and ( n3443 , n3252 , n3258 );
and ( n3444 , n3248 , n3258 );
or ( n3445 , n3442 , n3443 , n3444 );
xor ( n3446 , n3441 , n3445 );
and ( n3447 , n3233 , n3234 );
and ( n3448 , n3234 , n3236 );
and ( n3449 , n3233 , n3236 );
or ( n3450 , n3447 , n3448 , n3449 );
and ( n3451 , n1383 , n1134 );
and ( n3452 , n1580 , n1034 );
xor ( n3453 , n3451 , n3452 );
and ( n3454 , n1694 , n940 );
xor ( n3455 , n3453 , n3454 );
xor ( n3456 , n3450 , n3455 );
and ( n3457 , n1047 , n1551 );
and ( n3458 , n1164 , n1424 );
xor ( n3459 , n3457 , n3458 );
buf ( n3460 , n1287 );
xor ( n3461 , n3459 , n3460 );
xor ( n3462 , n3456 , n3461 );
xor ( n3463 , n3446 , n3462 );
xor ( n3464 , n3437 , n3463 );
and ( n3465 , n3264 , n3269 );
and ( n3466 , n3269 , n3276 );
and ( n3467 , n3264 , n3276 );
or ( n3468 , n3465 , n3466 , n3467 );
and ( n3469 , n3254 , n3255 );
and ( n3470 , n3255 , n3257 );
and ( n3471 , n3254 , n3257 );
or ( n3472 , n3469 , n3470 , n3471 );
and ( n3473 , n3265 , n3266 );
and ( n3474 , n3266 , n3268 );
and ( n3475 , n3265 , n3268 );
or ( n3476 , n3473 , n3474 , n3475 );
xor ( n3477 , n3472 , n3476 );
and ( n3478 , n783 , n2100 );
and ( n3479 , n856 , n1882 );
xor ( n3480 , n3478 , n3479 );
and ( n3481 , n925 , n1738 );
xor ( n3482 , n3480 , n3481 );
xor ( n3483 , n3477 , n3482 );
xor ( n3484 , n3468 , n3483 );
and ( n3485 , n3272 , n3273 );
and ( n3486 , n3273 , n3275 );
and ( n3487 , n3272 , n3275 );
or ( n3488 , n3485 , n3486 , n3487 );
and ( n3489 , n632 , n2739 );
and ( n3490 , n671 , n2544 );
xor ( n3491 , n3489 , n3490 );
and ( n3492 , n715 , n2298 );
xor ( n3493 , n3491 , n3492 );
xor ( n3494 , n3488 , n3493 );
buf ( n3495 , n448 );
and ( n3496 , n599 , n3495 );
and ( n3497 , n608 , n3271 );
xor ( n3498 , n3496 , n3497 );
and ( n3499 , n611 , n2981 );
xor ( n3500 , n3498 , n3499 );
xor ( n3501 , n3494 , n3500 );
xor ( n3502 , n3484 , n3501 );
xor ( n3503 , n3464 , n3502 );
xor ( n3504 , n3433 , n3503 );
and ( n3505 , n3177 , n3190 );
and ( n3506 , n3190 , n3206 );
and ( n3507 , n3177 , n3206 );
or ( n3508 , n3505 , n3506 , n3507 );
and ( n3509 , n3217 , n3221 );
and ( n3510 , n3221 , n3238 );
and ( n3511 , n3217 , n3238 );
or ( n3512 , n3509 , n3510 , n3511 );
xor ( n3513 , n3508 , n3512 );
and ( n3514 , n3195 , n3199 );
and ( n3515 , n3199 , n3205 );
and ( n3516 , n3195 , n3205 );
or ( n3517 , n3514 , n3515 , n3516 );
and ( n3518 , n3201 , n3202 );
and ( n3519 , n3202 , n3204 );
and ( n3520 , n3201 , n3204 );
or ( n3521 , n3518 , n3519 , n3520 );
and ( n3522 , n3227 , n3228 );
and ( n3523 , n3228 , n3230 );
and ( n3524 , n3227 , n3230 );
or ( n3525 , n3522 , n3523 , n3524 );
xor ( n3526 , n3521 , n3525 );
and ( n3527 , n1933 , n840 );
and ( n3528 , n2120 , n771 );
xor ( n3529 , n3527 , n3528 );
and ( n3530 , n2324 , n719 );
xor ( n3531 , n3529 , n3530 );
xor ( n3532 , n3526 , n3531 );
xor ( n3533 , n3517 , n3532 );
and ( n3534 , n3185 , n3186 );
and ( n3535 , n3186 , n3188 );
and ( n3536 , n3185 , n3188 );
or ( n3537 , n3534 , n3535 , n3536 );
and ( n3538 , n2462 , n663 );
and ( n3539 , n2779 , n635 );
xor ( n3540 , n3538 , n3539 );
and ( n3541 , n3024 , n606 );
xor ( n3542 , n3540 , n3541 );
xor ( n3543 , n3537 , n3542 );
and ( n3544 , n3182 , n615 );
buf ( n3545 , n448 );
and ( n3546 , n3545 , n612 );
xor ( n3547 , n3544 , n3546 );
xor ( n3548 , n3543 , n3547 );
xor ( n3549 , n3533 , n3548 );
xor ( n3550 , n3513 , n3549 );
xor ( n3551 , n3504 , n3550 );
xor ( n3552 , n3429 , n3551 );
and ( n3553 , n3181 , n3183 );
and ( n3554 , n3183 , n3189 );
and ( n3555 , n3181 , n3189 );
or ( n3556 , n3553 , n3554 , n3555 );
and ( n3557 , n3168 , n3172 );
and ( n3558 , n3172 , n3207 );
and ( n3559 , n3168 , n3207 );
or ( n3560 , n3557 , n3558 , n3559 );
xor ( n3561 , n3556 , n3560 );
xor ( n3562 , n3552 , n3561 );
xor ( n3563 , n3425 , n3562 );
and ( n3564 , n3288 , n3292 );
and ( n3565 , n3293 , n3296 );
or ( n3566 , n3564 , n3565 );
xor ( n3567 , n3563 , n3566 );
buf ( n3568 , n3567 );
buf ( n3569 , n3568 );
not ( n3570 , n3569 );
buf ( n3571 , n520 );
not ( n3572 , n3571 );
nor ( n3573 , n3570 , n3572 );
xor ( n3574 , n3419 , n3573 );
xor ( n3575 , n3308 , n3416 );
nor ( n3576 , n3300 , n3572 );
and ( n3577 , n3575 , n3576 );
xor ( n3578 , n3575 , n3576 );
xor ( n3579 , n3312 , n3414 );
nor ( n3580 , n3043 , n3572 );
and ( n3581 , n3579 , n3580 );
xor ( n3582 , n3579 , n3580 );
xor ( n3583 , n3316 , n3412 );
nor ( n3584 , n2797 , n3572 );
and ( n3585 , n3583 , n3584 );
xor ( n3586 , n3583 , n3584 );
xor ( n3587 , n3320 , n3410 );
nor ( n3588 , n2566 , n3572 );
and ( n3589 , n3587 , n3588 );
xor ( n3590 , n3587 , n3588 );
xor ( n3591 , n3324 , n3408 );
nor ( n3592 , n2343 , n3572 );
and ( n3593 , n3591 , n3592 );
xor ( n3594 , n3591 , n3592 );
xor ( n3595 , n3328 , n3406 );
nor ( n3596 , n2137 , n3572 );
and ( n3597 , n3595 , n3596 );
xor ( n3598 , n3595 , n3596 );
xor ( n3599 , n3332 , n3404 );
nor ( n3600 , n1945 , n3572 );
and ( n3601 , n3599 , n3600 );
xor ( n3602 , n3599 , n3600 );
xor ( n3603 , n3336 , n3402 );
nor ( n3604 , n1766 , n3572 );
and ( n3605 , n3603 , n3604 );
xor ( n3606 , n3603 , n3604 );
xor ( n3607 , n3340 , n3400 );
nor ( n3608 , n1598 , n3572 );
and ( n3609 , n3607 , n3608 );
xor ( n3610 , n3607 , n3608 );
xor ( n3611 , n3344 , n3398 );
nor ( n3612 , n1445 , n3572 );
and ( n3613 , n3611 , n3612 );
xor ( n3614 , n3611 , n3612 );
xor ( n3615 , n3348 , n3396 );
nor ( n3616 , n1303 , n3572 );
and ( n3617 , n3615 , n3616 );
xor ( n3618 , n3615 , n3616 );
xor ( n3619 , n3352 , n3394 );
nor ( n3620 , n1176 , n3572 );
and ( n3621 , n3619 , n3620 );
xor ( n3622 , n3619 , n3620 );
xor ( n3623 , n3356 , n3392 );
nor ( n3624 , n1062 , n3572 );
and ( n3625 , n3623 , n3624 );
xor ( n3626 , n3623 , n3624 );
xor ( n3627 , n3360 , n3390 );
nor ( n3628 , n958 , n3572 );
and ( n3629 , n3627 , n3628 );
xor ( n3630 , n3627 , n3628 );
xor ( n3631 , n3364 , n3388 );
nor ( n3632 , n868 , n3572 );
and ( n3633 , n3631 , n3632 );
xor ( n3634 , n3631 , n3632 );
xor ( n3635 , n3368 , n3386 );
nor ( n3636 , n796 , n3572 );
and ( n3637 , n3635 , n3636 );
xor ( n3638 , n3635 , n3636 );
xor ( n3639 , n3372 , n3384 );
nor ( n3640 , n733 , n3572 );
and ( n3641 , n3639 , n3640 );
xor ( n3642 , n3639 , n3640 );
xor ( n3643 , n3377 , n3382 );
nor ( n3644 , n684 , n3572 );
and ( n3645 , n3643 , n3644 );
xor ( n3646 , n3643 , n3644 );
xor ( n3647 , n3379 , n3380 );
buf ( n3648 , n3647 );
nor ( n3649 , n646 , n3572 );
and ( n3650 , n3648 , n3649 );
xor ( n3651 , n3648 , n3649 );
nor ( n3652 , n601 , n3045 );
buf ( n3653 , n3652 );
nor ( n3654 , n622 , n3572 );
and ( n3655 , n3653 , n3654 );
buf ( n3656 , n3655 );
and ( n3657 , n3651 , n3656 );
or ( n3658 , n3650 , n3657 );
and ( n3659 , n3646 , n3658 );
or ( n3660 , n3645 , n3659 );
and ( n3661 , n3642 , n3660 );
or ( n3662 , n3641 , n3661 );
and ( n3663 , n3638 , n3662 );
or ( n3664 , n3637 , n3663 );
and ( n3665 , n3634 , n3664 );
or ( n3666 , n3633 , n3665 );
and ( n3667 , n3630 , n3666 );
or ( n3668 , n3629 , n3667 );
and ( n3669 , n3626 , n3668 );
or ( n3670 , n3625 , n3669 );
and ( n3671 , n3622 , n3670 );
or ( n3672 , n3621 , n3671 );
and ( n3673 , n3618 , n3672 );
or ( n3674 , n3617 , n3673 );
and ( n3675 , n3614 , n3674 );
or ( n3676 , n3613 , n3675 );
and ( n3677 , n3610 , n3676 );
or ( n3678 , n3609 , n3677 );
and ( n3679 , n3606 , n3678 );
or ( n3680 , n3605 , n3679 );
and ( n3681 , n3602 , n3680 );
or ( n3682 , n3601 , n3681 );
and ( n3683 , n3598 , n3682 );
or ( n3684 , n3597 , n3683 );
and ( n3685 , n3594 , n3684 );
or ( n3686 , n3593 , n3685 );
and ( n3687 , n3590 , n3686 );
or ( n3688 , n3589 , n3687 );
and ( n3689 , n3586 , n3688 );
or ( n3690 , n3585 , n3689 );
and ( n3691 , n3582 , n3690 );
or ( n3692 , n3581 , n3691 );
and ( n3693 , n3578 , n3692 );
or ( n3694 , n3577 , n3693 );
xor ( n3695 , n3574 , n3694 );
and ( n3696 , n3556 , n3560 );
and ( n3697 , n3429 , n3551 );
and ( n3698 , n3551 , n3561 );
and ( n3699 , n3429 , n3561 );
or ( n3700 , n3697 , n3698 , n3699 );
xor ( n3701 , n3696 , n3700 );
and ( n3702 , n3433 , n3503 );
and ( n3703 , n3503 , n3550 );
and ( n3704 , n3433 , n3550 );
or ( n3705 , n3702 , n3703 , n3704 );
and ( n3706 , n3437 , n3463 );
and ( n3707 , n3463 , n3502 );
and ( n3708 , n3437 , n3502 );
or ( n3709 , n3706 , n3707 , n3708 );
and ( n3710 , n3468 , n3483 );
and ( n3711 , n3483 , n3501 );
and ( n3712 , n3468 , n3501 );
or ( n3713 , n3710 , n3711 , n3712 );
and ( n3714 , n3450 , n3455 );
and ( n3715 , n3455 , n3461 );
and ( n3716 , n3450 , n3461 );
or ( n3717 , n3714 , n3715 , n3716 );
and ( n3718 , n3472 , n3476 );
and ( n3719 , n3476 , n3482 );
and ( n3720 , n3472 , n3482 );
or ( n3721 , n3718 , n3719 , n3720 );
xor ( n3722 , n3717 , n3721 );
and ( n3723 , n3457 , n3458 );
and ( n3724 , n3458 , n3460 );
and ( n3725 , n3457 , n3460 );
or ( n3726 , n3723 , n3724 , n3725 );
and ( n3727 , n1047 , n1738 );
and ( n3728 , n1164 , n1551 );
xor ( n3729 , n3727 , n3728 );
and ( n3730 , n1287 , n1424 );
xor ( n3731 , n3729 , n3730 );
xor ( n3732 , n3726 , n3731 );
and ( n3733 , n1383 , n1254 );
and ( n3734 , n1580 , n1134 );
xor ( n3735 , n3733 , n3734 );
and ( n3736 , n1694 , n1034 );
xor ( n3737 , n3735 , n3736 );
xor ( n3738 , n3732 , n3737 );
xor ( n3739 , n3722 , n3738 );
xor ( n3740 , n3713 , n3739 );
and ( n3741 , n3488 , n3493 );
and ( n3742 , n3493 , n3500 );
and ( n3743 , n3488 , n3500 );
or ( n3744 , n3741 , n3742 , n3743 );
and ( n3745 , n3496 , n3497 );
and ( n3746 , n3497 , n3499 );
and ( n3747 , n3496 , n3499 );
or ( n3748 , n3745 , n3746 , n3747 );
buf ( n3749 , n447 );
and ( n3750 , n599 , n3749 );
and ( n3751 , n608 , n3495 );
xor ( n3752 , n3750 , n3751 );
and ( n3753 , n611 , n3271 );
xor ( n3754 , n3752 , n3753 );
xor ( n3755 , n3748 , n3754 );
and ( n3756 , n632 , n2981 );
and ( n3757 , n671 , n2739 );
xor ( n3758 , n3756 , n3757 );
and ( n3759 , n715 , n2544 );
xor ( n3760 , n3758 , n3759 );
xor ( n3761 , n3755 , n3760 );
xor ( n3762 , n3744 , n3761 );
and ( n3763 , n3478 , n3479 );
and ( n3764 , n3479 , n3481 );
and ( n3765 , n3478 , n3481 );
or ( n3766 , n3763 , n3764 , n3765 );
and ( n3767 , n3489 , n3490 );
and ( n3768 , n3490 , n3492 );
and ( n3769 , n3489 , n3492 );
or ( n3770 , n3767 , n3768 , n3769 );
xor ( n3771 , n3766 , n3770 );
and ( n3772 , n783 , n2298 );
and ( n3773 , n856 , n2100 );
xor ( n3774 , n3772 , n3773 );
and ( n3775 , n925 , n1882 );
xor ( n3776 , n3774 , n3775 );
xor ( n3777 , n3771 , n3776 );
xor ( n3778 , n3762 , n3777 );
xor ( n3779 , n3740 , n3778 );
xor ( n3780 , n3709 , n3779 );
and ( n3781 , n3441 , n3445 );
and ( n3782 , n3445 , n3462 );
and ( n3783 , n3441 , n3462 );
or ( n3784 , n3781 , n3782 , n3783 );
and ( n3785 , n3517 , n3532 );
and ( n3786 , n3532 , n3548 );
and ( n3787 , n3517 , n3548 );
or ( n3788 , n3785 , n3786 , n3787 );
xor ( n3789 , n3784 , n3788 );
and ( n3790 , n3521 , n3525 );
and ( n3791 , n3525 , n3531 );
and ( n3792 , n3521 , n3531 );
or ( n3793 , n3790 , n3791 , n3792 );
and ( n3794 , n3538 , n3539 );
and ( n3795 , n3539 , n3541 );
and ( n3796 , n3538 , n3541 );
or ( n3797 , n3794 , n3795 , n3796 );
and ( n3798 , n3182 , n606 );
and ( n3799 , n3545 , n615 );
xor ( n3800 , n3798 , n3799 );
buf ( n3801 , n447 );
and ( n3802 , n3801 , n612 );
xor ( n3803 , n3800 , n3802 );
xor ( n3804 , n3797 , n3803 );
and ( n3805 , n2462 , n719 );
and ( n3806 , n2779 , n663 );
xor ( n3807 , n3805 , n3806 );
and ( n3808 , n3024 , n635 );
xor ( n3809 , n3807 , n3808 );
xor ( n3810 , n3804 , n3809 );
xor ( n3811 , n3793 , n3810 );
and ( n3812 , n3527 , n3528 );
and ( n3813 , n3528 , n3530 );
and ( n3814 , n3527 , n3530 );
or ( n3815 , n3812 , n3813 , n3814 );
and ( n3816 , n3451 , n3452 );
and ( n3817 , n3452 , n3454 );
and ( n3818 , n3451 , n3454 );
or ( n3819 , n3816 , n3817 , n3818 );
xor ( n3820 , n3815 , n3819 );
and ( n3821 , n1933 , n940 );
and ( n3822 , n2120 , n840 );
xor ( n3823 , n3821 , n3822 );
and ( n3824 , n2324 , n771 );
xor ( n3825 , n3823 , n3824 );
xor ( n3826 , n3820 , n3825 );
xor ( n3827 , n3811 , n3826 );
xor ( n3828 , n3789 , n3827 );
xor ( n3829 , n3780 , n3828 );
xor ( n3830 , n3705 , n3829 );
and ( n3831 , n3508 , n3512 );
and ( n3832 , n3512 , n3549 );
and ( n3833 , n3508 , n3549 );
or ( n3834 , n3831 , n3832 , n3833 );
and ( n3835 , n3544 , n3546 );
and ( n3836 , n3537 , n3542 );
and ( n3837 , n3542 , n3547 );
and ( n3838 , n3537 , n3547 );
or ( n3839 , n3836 , n3837 , n3838 );
xor ( n3840 , n3835 , n3839 );
xor ( n3841 , n3834 , n3840 );
xor ( n3842 , n3830 , n3841 );
xor ( n3843 , n3701 , n3842 );
and ( n3844 , n3420 , n3424 );
and ( n3845 , n3424 , n3562 );
and ( n3846 , n3420 , n3562 );
or ( n3847 , n3844 , n3845 , n3846 );
xor ( n3848 , n3843 , n3847 );
and ( n3849 , n3563 , n3566 );
xor ( n3850 , n3848 , n3849 );
buf ( n3851 , n3850 );
buf ( n3852 , n3851 );
not ( n3853 , n3852 );
buf ( n3854 , n521 );
not ( n3855 , n3854 );
nor ( n3856 , n3853 , n3855 );
xor ( n3857 , n3695 , n3856 );
xor ( n3858 , n3578 , n3692 );
nor ( n3859 , n3570 , n3855 );
and ( n3860 , n3858 , n3859 );
xor ( n3861 , n3858 , n3859 );
xor ( n3862 , n3582 , n3690 );
nor ( n3863 , n3300 , n3855 );
and ( n3864 , n3862 , n3863 );
xor ( n3865 , n3862 , n3863 );
xor ( n3866 , n3586 , n3688 );
nor ( n3867 , n3043 , n3855 );
and ( n3868 , n3866 , n3867 );
xor ( n3869 , n3866 , n3867 );
xor ( n3870 , n3590 , n3686 );
nor ( n3871 , n2797 , n3855 );
and ( n3872 , n3870 , n3871 );
xor ( n3873 , n3870 , n3871 );
xor ( n3874 , n3594 , n3684 );
nor ( n3875 , n2566 , n3855 );
and ( n3876 , n3874 , n3875 );
xor ( n3877 , n3874 , n3875 );
xor ( n3878 , n3598 , n3682 );
nor ( n3879 , n2343 , n3855 );
and ( n3880 , n3878 , n3879 );
xor ( n3881 , n3878 , n3879 );
xor ( n3882 , n3602 , n3680 );
nor ( n3883 , n2137 , n3855 );
and ( n3884 , n3882 , n3883 );
xor ( n3885 , n3882 , n3883 );
xor ( n3886 , n3606 , n3678 );
nor ( n3887 , n1945 , n3855 );
and ( n3888 , n3886 , n3887 );
xor ( n3889 , n3886 , n3887 );
xor ( n3890 , n3610 , n3676 );
nor ( n3891 , n1766 , n3855 );
and ( n3892 , n3890 , n3891 );
xor ( n3893 , n3890 , n3891 );
xor ( n3894 , n3614 , n3674 );
nor ( n3895 , n1598 , n3855 );
and ( n3896 , n3894 , n3895 );
xor ( n3897 , n3894 , n3895 );
xor ( n3898 , n3618 , n3672 );
nor ( n3899 , n1445 , n3855 );
and ( n3900 , n3898 , n3899 );
xor ( n3901 , n3898 , n3899 );
xor ( n3902 , n3622 , n3670 );
nor ( n3903 , n1303 , n3855 );
and ( n3904 , n3902 , n3903 );
xor ( n3905 , n3902 , n3903 );
xor ( n3906 , n3626 , n3668 );
nor ( n3907 , n1176 , n3855 );
and ( n3908 , n3906 , n3907 );
xor ( n3909 , n3906 , n3907 );
xor ( n3910 , n3630 , n3666 );
nor ( n3911 , n1062 , n3855 );
and ( n3912 , n3910 , n3911 );
xor ( n3913 , n3910 , n3911 );
xor ( n3914 , n3634 , n3664 );
nor ( n3915 , n958 , n3855 );
and ( n3916 , n3914 , n3915 );
xor ( n3917 , n3914 , n3915 );
xor ( n3918 , n3638 , n3662 );
nor ( n3919 , n868 , n3855 );
and ( n3920 , n3918 , n3919 );
xor ( n3921 , n3918 , n3919 );
xor ( n3922 , n3642 , n3660 );
nor ( n3923 , n796 , n3855 );
and ( n3924 , n3922 , n3923 );
xor ( n3925 , n3922 , n3923 );
xor ( n3926 , n3646 , n3658 );
nor ( n3927 , n733 , n3855 );
and ( n3928 , n3926 , n3927 );
xor ( n3929 , n3926 , n3927 );
xor ( n3930 , n3651 , n3656 );
nor ( n3931 , n684 , n3855 );
and ( n3932 , n3930 , n3931 );
xor ( n3933 , n3930 , n3931 );
xor ( n3934 , n3653 , n3654 );
buf ( n3935 , n3934 );
nor ( n3936 , n646 , n3855 );
and ( n3937 , n3935 , n3936 );
xor ( n3938 , n3935 , n3936 );
nor ( n3939 , n601 , n3302 );
buf ( n3940 , n3939 );
nor ( n3941 , n622 , n3855 );
and ( n3942 , n3940 , n3941 );
buf ( n3943 , n3942 );
and ( n3944 , n3938 , n3943 );
or ( n3945 , n3937 , n3944 );
and ( n3946 , n3933 , n3945 );
or ( n3947 , n3932 , n3946 );
and ( n3948 , n3929 , n3947 );
or ( n3949 , n3928 , n3948 );
and ( n3950 , n3925 , n3949 );
or ( n3951 , n3924 , n3950 );
and ( n3952 , n3921 , n3951 );
or ( n3953 , n3920 , n3952 );
and ( n3954 , n3917 , n3953 );
or ( n3955 , n3916 , n3954 );
and ( n3956 , n3913 , n3955 );
or ( n3957 , n3912 , n3956 );
and ( n3958 , n3909 , n3957 );
or ( n3959 , n3908 , n3958 );
and ( n3960 , n3905 , n3959 );
or ( n3961 , n3904 , n3960 );
and ( n3962 , n3901 , n3961 );
or ( n3963 , n3900 , n3962 );
and ( n3964 , n3897 , n3963 );
or ( n3965 , n3896 , n3964 );
and ( n3966 , n3893 , n3965 );
or ( n3967 , n3892 , n3966 );
and ( n3968 , n3889 , n3967 );
or ( n3969 , n3888 , n3968 );
and ( n3970 , n3885 , n3969 );
or ( n3971 , n3884 , n3970 );
and ( n3972 , n3881 , n3971 );
or ( n3973 , n3880 , n3972 );
and ( n3974 , n3877 , n3973 );
or ( n3975 , n3876 , n3974 );
and ( n3976 , n3873 , n3975 );
or ( n3977 , n3872 , n3976 );
and ( n3978 , n3869 , n3977 );
or ( n3979 , n3868 , n3978 );
and ( n3980 , n3865 , n3979 );
or ( n3981 , n3864 , n3980 );
and ( n3982 , n3861 , n3981 );
or ( n3983 , n3860 , n3982 );
xor ( n3984 , n3857 , n3983 );
and ( n3985 , n3834 , n3840 );
and ( n3986 , n3705 , n3829 );
and ( n3987 , n3829 , n3841 );
and ( n3988 , n3705 , n3841 );
or ( n3989 , n3986 , n3987 , n3988 );
xor ( n3990 , n3985 , n3989 );
and ( n3991 , n3709 , n3779 );
and ( n3992 , n3779 , n3828 );
and ( n3993 , n3709 , n3828 );
or ( n3994 , n3991 , n3992 , n3993 );
and ( n3995 , n3713 , n3739 );
and ( n3996 , n3739 , n3778 );
and ( n3997 , n3713 , n3778 );
or ( n3998 , n3995 , n3996 , n3997 );
and ( n3999 , n3717 , n3721 );
and ( n4000 , n3721 , n3738 );
and ( n4001 , n3717 , n3738 );
or ( n4002 , n3999 , n4000 , n4001 );
and ( n4003 , n3793 , n3810 );
and ( n4004 , n3810 , n3826 );
and ( n4005 , n3793 , n3826 );
or ( n4006 , n4003 , n4004 , n4005 );
xor ( n4007 , n4002 , n4006 );
and ( n4008 , n3815 , n3819 );
and ( n4009 , n3819 , n3825 );
and ( n4010 , n3815 , n3825 );
or ( n4011 , n4008 , n4009 , n4010 );
and ( n4012 , n3805 , n3806 );
and ( n4013 , n3806 , n3808 );
and ( n4014 , n3805 , n3808 );
or ( n4015 , n4012 , n4013 , n4014 );
and ( n4016 , n3182 , n635 );
and ( n4017 , n3545 , n606 );
xor ( n4018 , n4016 , n4017 );
and ( n4019 , n3801 , n615 );
xor ( n4020 , n4018 , n4019 );
xor ( n4021 , n4015 , n4020 );
and ( n4022 , n2462 , n771 );
and ( n4023 , n2779 , n719 );
xor ( n4024 , n4022 , n4023 );
and ( n4025 , n3024 , n663 );
xor ( n4026 , n4024 , n4025 );
xor ( n4027 , n4021 , n4026 );
xor ( n4028 , n4011 , n4027 );
and ( n4029 , n3821 , n3822 );
and ( n4030 , n3822 , n3824 );
and ( n4031 , n3821 , n3824 );
or ( n4032 , n4029 , n4030 , n4031 );
and ( n4033 , n3733 , n3734 );
and ( n4034 , n3734 , n3736 );
and ( n4035 , n3733 , n3736 );
or ( n4036 , n4033 , n4034 , n4035 );
xor ( n4037 , n4032 , n4036 );
and ( n4038 , n1933 , n1034 );
and ( n4039 , n2120 , n940 );
xor ( n4040 , n4038 , n4039 );
and ( n4041 , n2324 , n840 );
xor ( n4042 , n4040 , n4041 );
xor ( n4043 , n4037 , n4042 );
xor ( n4044 , n4028 , n4043 );
xor ( n4045 , n4007 , n4044 );
xor ( n4046 , n3998 , n4045 );
and ( n4047 , n3744 , n3761 );
and ( n4048 , n3761 , n3777 );
and ( n4049 , n3744 , n3777 );
or ( n4050 , n4047 , n4048 , n4049 );
and ( n4051 , n3726 , n3731 );
and ( n4052 , n3731 , n3737 );
and ( n4053 , n3726 , n3737 );
or ( n4054 , n4051 , n4052 , n4053 );
and ( n4055 , n3766 , n3770 );
and ( n4056 , n3770 , n3776 );
and ( n4057 , n3766 , n3776 );
or ( n4058 , n4055 , n4056 , n4057 );
xor ( n4059 , n4054 , n4058 );
and ( n4060 , n3727 , n3728 );
and ( n4061 , n3728 , n3730 );
and ( n4062 , n3727 , n3730 );
or ( n4063 , n4060 , n4061 , n4062 );
and ( n4064 , n1047 , n1882 );
and ( n4065 , n1164 , n1738 );
xor ( n4066 , n4064 , n4065 );
and ( n4067 , n1287 , n1551 );
xor ( n4068 , n4066 , n4067 );
xor ( n4069 , n4063 , n4068 );
buf ( n4070 , n1383 );
and ( n4071 , n1580 , n1254 );
xor ( n4072 , n4070 , n4071 );
and ( n4073 , n1694 , n1134 );
xor ( n4074 , n4072 , n4073 );
xor ( n4075 , n4069 , n4074 );
xor ( n4076 , n4059 , n4075 );
xor ( n4077 , n4050 , n4076 );
and ( n4078 , n3748 , n3754 );
and ( n4079 , n3754 , n3760 );
and ( n4080 , n3748 , n3760 );
or ( n4081 , n4078 , n4079 , n4080 );
and ( n4082 , n3756 , n3757 );
and ( n4083 , n3757 , n3759 );
and ( n4084 , n3756 , n3759 );
or ( n4085 , n4082 , n4083 , n4084 );
and ( n4086 , n3772 , n3773 );
and ( n4087 , n3773 , n3775 );
and ( n4088 , n3772 , n3775 );
or ( n4089 , n4086 , n4087 , n4088 );
xor ( n4090 , n4085 , n4089 );
and ( n4091 , n783 , n2544 );
and ( n4092 , n856 , n2298 );
xor ( n4093 , n4091 , n4092 );
and ( n4094 , n925 , n2100 );
xor ( n4095 , n4093 , n4094 );
xor ( n4096 , n4090 , n4095 );
xor ( n4097 , n4081 , n4096 );
and ( n4098 , n3750 , n3751 );
and ( n4099 , n3751 , n3753 );
and ( n4100 , n3750 , n3753 );
or ( n4101 , n4098 , n4099 , n4100 );
buf ( n4102 , n446 );
and ( n4103 , n599 , n4102 );
and ( n4104 , n608 , n3749 );
xor ( n4105 , n4103 , n4104 );
and ( n4106 , n611 , n3495 );
xor ( n4107 , n4105 , n4106 );
xor ( n4108 , n4101 , n4107 );
and ( n4109 , n632 , n3271 );
and ( n4110 , n671 , n2981 );
xor ( n4111 , n4109 , n4110 );
and ( n4112 , n715 , n2739 );
xor ( n4113 , n4111 , n4112 );
xor ( n4114 , n4108 , n4113 );
xor ( n4115 , n4097 , n4114 );
xor ( n4116 , n4077 , n4115 );
xor ( n4117 , n4046 , n4116 );
xor ( n4118 , n3994 , n4117 );
and ( n4119 , n3784 , n3788 );
and ( n4120 , n3788 , n3827 );
and ( n4121 , n3784 , n3827 );
or ( n4122 , n4119 , n4120 , n4121 );
and ( n4123 , n3835 , n3839 );
and ( n4124 , n3797 , n3803 );
and ( n4125 , n3803 , n3809 );
and ( n4126 , n3797 , n3809 );
or ( n4127 , n4124 , n4125 , n4126 );
and ( n4128 , n3798 , n3799 );
and ( n4129 , n3799 , n3802 );
and ( n4130 , n3798 , n3802 );
or ( n4131 , n4128 , n4129 , n4130 );
buf ( n4132 , n446 );
and ( n4133 , n4132 , n612 );
xor ( n4134 , n4131 , n4133 );
xor ( n4135 , n4127 , n4134 );
xor ( n4136 , n4123 , n4135 );
xor ( n4137 , n4122 , n4136 );
xor ( n4138 , n4118 , n4137 );
xor ( n4139 , n3990 , n4138 );
and ( n4140 , n3696 , n3700 );
and ( n4141 , n3700 , n3842 );
and ( n4142 , n3696 , n3842 );
or ( n4143 , n4140 , n4141 , n4142 );
xor ( n4144 , n4139 , n4143 );
and ( n4145 , n3843 , n3847 );
and ( n4146 , n3848 , n3849 );
or ( n4147 , n4145 , n4146 );
xor ( n4148 , n4144 , n4147 );
buf ( n4149 , n4148 );
buf ( n4150 , n4149 );
not ( n4151 , n4150 );
buf ( n4152 , n522 );
not ( n4153 , n4152 );
nor ( n4154 , n4151 , n4153 );
xor ( n4155 , n3984 , n4154 );
xor ( n4156 , n3861 , n3981 );
nor ( n4157 , n3853 , n4153 );
and ( n4158 , n4156 , n4157 );
xor ( n4159 , n4156 , n4157 );
xor ( n4160 , n3865 , n3979 );
nor ( n4161 , n3570 , n4153 );
and ( n4162 , n4160 , n4161 );
xor ( n4163 , n4160 , n4161 );
xor ( n4164 , n3869 , n3977 );
nor ( n4165 , n3300 , n4153 );
and ( n4166 , n4164 , n4165 );
xor ( n4167 , n4164 , n4165 );
xor ( n4168 , n3873 , n3975 );
nor ( n4169 , n3043 , n4153 );
and ( n4170 , n4168 , n4169 );
xor ( n4171 , n4168 , n4169 );
xor ( n4172 , n3877 , n3973 );
nor ( n4173 , n2797 , n4153 );
and ( n4174 , n4172 , n4173 );
xor ( n4175 , n4172 , n4173 );
xor ( n4176 , n3881 , n3971 );
nor ( n4177 , n2566 , n4153 );
and ( n4178 , n4176 , n4177 );
xor ( n4179 , n4176 , n4177 );
xor ( n4180 , n3885 , n3969 );
nor ( n4181 , n2343 , n4153 );
and ( n4182 , n4180 , n4181 );
xor ( n4183 , n4180 , n4181 );
xor ( n4184 , n3889 , n3967 );
nor ( n4185 , n2137 , n4153 );
and ( n4186 , n4184 , n4185 );
xor ( n4187 , n4184 , n4185 );
xor ( n4188 , n3893 , n3965 );
nor ( n4189 , n1945 , n4153 );
and ( n4190 , n4188 , n4189 );
xor ( n4191 , n4188 , n4189 );
xor ( n4192 , n3897 , n3963 );
nor ( n4193 , n1766 , n4153 );
and ( n4194 , n4192 , n4193 );
xor ( n4195 , n4192 , n4193 );
xor ( n4196 , n3901 , n3961 );
nor ( n4197 , n1598 , n4153 );
and ( n4198 , n4196 , n4197 );
xor ( n4199 , n4196 , n4197 );
xor ( n4200 , n3905 , n3959 );
nor ( n4201 , n1445 , n4153 );
and ( n4202 , n4200 , n4201 );
xor ( n4203 , n4200 , n4201 );
xor ( n4204 , n3909 , n3957 );
nor ( n4205 , n1303 , n4153 );
and ( n4206 , n4204 , n4205 );
xor ( n4207 , n4204 , n4205 );
xor ( n4208 , n3913 , n3955 );
nor ( n4209 , n1176 , n4153 );
and ( n4210 , n4208 , n4209 );
xor ( n4211 , n4208 , n4209 );
xor ( n4212 , n3917 , n3953 );
nor ( n4213 , n1062 , n4153 );
and ( n4214 , n4212 , n4213 );
xor ( n4215 , n4212 , n4213 );
xor ( n4216 , n3921 , n3951 );
nor ( n4217 , n958 , n4153 );
and ( n4218 , n4216 , n4217 );
xor ( n4219 , n4216 , n4217 );
xor ( n4220 , n3925 , n3949 );
nor ( n4221 , n868 , n4153 );
and ( n4222 , n4220 , n4221 );
xor ( n4223 , n4220 , n4221 );
xor ( n4224 , n3929 , n3947 );
nor ( n4225 , n796 , n4153 );
and ( n4226 , n4224 , n4225 );
xor ( n4227 , n4224 , n4225 );
xor ( n4228 , n3933 , n3945 );
nor ( n4229 , n733 , n4153 );
and ( n4230 , n4228 , n4229 );
xor ( n4231 , n4228 , n4229 );
xor ( n4232 , n3938 , n3943 );
nor ( n4233 , n684 , n4153 );
and ( n4234 , n4232 , n4233 );
xor ( n4235 , n4232 , n4233 );
xor ( n4236 , n3940 , n3941 );
buf ( n4237 , n4236 );
nor ( n4238 , n646 , n4153 );
and ( n4239 , n4237 , n4238 );
xor ( n4240 , n4237 , n4238 );
nor ( n4241 , n601 , n3572 );
buf ( n4242 , n4241 );
nor ( n4243 , n622 , n4153 );
and ( n4244 , n4242 , n4243 );
buf ( n4245 , n4244 );
and ( n4246 , n4240 , n4245 );
or ( n4247 , n4239 , n4246 );
and ( n4248 , n4235 , n4247 );
or ( n4249 , n4234 , n4248 );
and ( n4250 , n4231 , n4249 );
or ( n4251 , n4230 , n4250 );
and ( n4252 , n4227 , n4251 );
or ( n4253 , n4226 , n4252 );
and ( n4254 , n4223 , n4253 );
or ( n4255 , n4222 , n4254 );
and ( n4256 , n4219 , n4255 );
or ( n4257 , n4218 , n4256 );
and ( n4258 , n4215 , n4257 );
or ( n4259 , n4214 , n4258 );
and ( n4260 , n4211 , n4259 );
or ( n4261 , n4210 , n4260 );
and ( n4262 , n4207 , n4261 );
or ( n4263 , n4206 , n4262 );
and ( n4264 , n4203 , n4263 );
or ( n4265 , n4202 , n4264 );
and ( n4266 , n4199 , n4265 );
or ( n4267 , n4198 , n4266 );
and ( n4268 , n4195 , n4267 );
or ( n4269 , n4194 , n4268 );
and ( n4270 , n4191 , n4269 );
or ( n4271 , n4190 , n4270 );
and ( n4272 , n4187 , n4271 );
or ( n4273 , n4186 , n4272 );
and ( n4274 , n4183 , n4273 );
or ( n4275 , n4182 , n4274 );
and ( n4276 , n4179 , n4275 );
or ( n4277 , n4178 , n4276 );
and ( n4278 , n4175 , n4277 );
or ( n4279 , n4174 , n4278 );
and ( n4280 , n4171 , n4279 );
or ( n4281 , n4170 , n4280 );
and ( n4282 , n4167 , n4281 );
or ( n4283 , n4166 , n4282 );
and ( n4284 , n4163 , n4283 );
or ( n4285 , n4162 , n4284 );
and ( n4286 , n4159 , n4285 );
or ( n4287 , n4158 , n4286 );
xor ( n4288 , n4155 , n4287 );
and ( n4289 , n4122 , n4136 );
and ( n4290 , n3994 , n4117 );
and ( n4291 , n4117 , n4137 );
and ( n4292 , n3994 , n4137 );
or ( n4293 , n4290 , n4291 , n4292 );
xor ( n4294 , n4289 , n4293 );
and ( n4295 , n3998 , n4045 );
and ( n4296 , n4045 , n4116 );
and ( n4297 , n3998 , n4116 );
or ( n4298 , n4295 , n4296 , n4297 );
and ( n4299 , n4050 , n4076 );
and ( n4300 , n4076 , n4115 );
and ( n4301 , n4050 , n4115 );
or ( n4302 , n4299 , n4300 , n4301 );
and ( n4303 , n4011 , n4027 );
and ( n4304 , n4027 , n4043 );
and ( n4305 , n4011 , n4043 );
or ( n4306 , n4303 , n4304 , n4305 );
and ( n4307 , n4054 , n4058 );
and ( n4308 , n4058 , n4075 );
and ( n4309 , n4054 , n4075 );
or ( n4310 , n4307 , n4308 , n4309 );
xor ( n4311 , n4306 , n4310 );
and ( n4312 , n4032 , n4036 );
and ( n4313 , n4036 , n4042 );
and ( n4314 , n4032 , n4042 );
or ( n4315 , n4312 , n4313 , n4314 );
and ( n4316 , n4022 , n4023 );
and ( n4317 , n4023 , n4025 );
and ( n4318 , n4022 , n4025 );
or ( n4319 , n4316 , n4317 , n4318 );
and ( n4320 , n3182 , n663 );
and ( n4321 , n3545 , n635 );
xor ( n4322 , n4320 , n4321 );
and ( n4323 , n3801 , n606 );
xor ( n4324 , n4322 , n4323 );
xor ( n4325 , n4319 , n4324 );
and ( n4326 , n2462 , n840 );
and ( n4327 , n2779 , n771 );
xor ( n4328 , n4326 , n4327 );
and ( n4329 , n3024 , n719 );
xor ( n4330 , n4328 , n4329 );
xor ( n4331 , n4325 , n4330 );
xor ( n4332 , n4315 , n4331 );
and ( n4333 , n4038 , n4039 );
and ( n4334 , n4039 , n4041 );
and ( n4335 , n4038 , n4041 );
or ( n4336 , n4333 , n4334 , n4335 );
and ( n4337 , n4070 , n4071 );
and ( n4338 , n4071 , n4073 );
and ( n4339 , n4070 , n4073 );
or ( n4340 , n4337 , n4338 , n4339 );
xor ( n4341 , n4336 , n4340 );
and ( n4342 , n1933 , n1134 );
and ( n4343 , n2120 , n1034 );
xor ( n4344 , n4342 , n4343 );
and ( n4345 , n2324 , n940 );
xor ( n4346 , n4344 , n4345 );
xor ( n4347 , n4341 , n4346 );
xor ( n4348 , n4332 , n4347 );
xor ( n4349 , n4311 , n4348 );
xor ( n4350 , n4302 , n4349 );
and ( n4351 , n4081 , n4096 );
and ( n4352 , n4096 , n4114 );
and ( n4353 , n4081 , n4114 );
or ( n4354 , n4351 , n4352 , n4353 );
and ( n4355 , n4063 , n4068 );
and ( n4356 , n4068 , n4074 );
and ( n4357 , n4063 , n4074 );
or ( n4358 , n4355 , n4356 , n4357 );
and ( n4359 , n4085 , n4089 );
and ( n4360 , n4089 , n4095 );
and ( n4361 , n4085 , n4095 );
or ( n4362 , n4359 , n4360 , n4361 );
xor ( n4363 , n4358 , n4362 );
and ( n4364 , n4064 , n4065 );
and ( n4365 , n4065 , n4067 );
and ( n4366 , n4064 , n4067 );
or ( n4367 , n4364 , n4365 , n4366 );
and ( n4368 , n1047 , n2100 );
and ( n4369 , n1164 , n1882 );
xor ( n4370 , n4368 , n4369 );
and ( n4371 , n1287 , n1738 );
xor ( n4372 , n4370 , n4371 );
xor ( n4373 , n4367 , n4372 );
and ( n4374 , n1694 , n1254 );
buf ( n4375 , n4374 );
xor ( n4376 , n4373 , n4375 );
xor ( n4377 , n4363 , n4376 );
xor ( n4378 , n4354 , n4377 );
and ( n4379 , n4101 , n4107 );
and ( n4380 , n4107 , n4113 );
and ( n4381 , n4101 , n4113 );
or ( n4382 , n4379 , n4380 , n4381 );
and ( n4383 , n4091 , n4092 );
and ( n4384 , n4092 , n4094 );
and ( n4385 , n4091 , n4094 );
or ( n4386 , n4383 , n4384 , n4385 );
and ( n4387 , n4109 , n4110 );
and ( n4388 , n4110 , n4112 );
and ( n4389 , n4109 , n4112 );
or ( n4390 , n4387 , n4388 , n4389 );
xor ( n4391 , n4386 , n4390 );
and ( n4392 , n783 , n2739 );
and ( n4393 , n856 , n2544 );
xor ( n4394 , n4392 , n4393 );
and ( n4395 , n925 , n2298 );
xor ( n4396 , n4394 , n4395 );
xor ( n4397 , n4391 , n4396 );
xor ( n4398 , n4382 , n4397 );
and ( n4399 , n4103 , n4104 );
and ( n4400 , n4104 , n4106 );
and ( n4401 , n4103 , n4106 );
or ( n4402 , n4399 , n4400 , n4401 );
buf ( n4403 , n445 );
and ( n4404 , n599 , n4403 );
and ( n4405 , n608 , n4102 );
xor ( n4406 , n4404 , n4405 );
and ( n4407 , n611 , n3749 );
xor ( n4408 , n4406 , n4407 );
xor ( n4409 , n4402 , n4408 );
and ( n4410 , n632 , n3495 );
and ( n4411 , n671 , n3271 );
xor ( n4412 , n4410 , n4411 );
and ( n4413 , n715 , n2981 );
xor ( n4414 , n4412 , n4413 );
xor ( n4415 , n4409 , n4414 );
xor ( n4416 , n4398 , n4415 );
xor ( n4417 , n4378 , n4416 );
xor ( n4418 , n4350 , n4417 );
xor ( n4419 , n4298 , n4418 );
and ( n4420 , n4002 , n4006 );
and ( n4421 , n4006 , n4044 );
and ( n4422 , n4002 , n4044 );
or ( n4423 , n4420 , n4421 , n4422 );
and ( n4424 , n4123 , n4135 );
xor ( n4425 , n4423 , n4424 );
and ( n4426 , n4127 , n4134 );
and ( n4427 , n4015 , n4020 );
and ( n4428 , n4020 , n4026 );
and ( n4429 , n4015 , n4026 );
or ( n4430 , n4427 , n4428 , n4429 );
and ( n4431 , n4131 , n4133 );
xor ( n4432 , n4430 , n4431 );
and ( n4433 , n4016 , n4017 );
and ( n4434 , n4017 , n4019 );
and ( n4435 , n4016 , n4019 );
or ( n4436 , n4433 , n4434 , n4435 );
and ( n4437 , n4132 , n615 );
buf ( n4438 , n445 );
and ( n4439 , n4438 , n612 );
xor ( n4440 , n4437 , n4439 );
xor ( n4441 , n4436 , n4440 );
xor ( n4442 , n4432 , n4441 );
xor ( n4443 , n4426 , n4442 );
xor ( n4444 , n4425 , n4443 );
xor ( n4445 , n4419 , n4444 );
xor ( n4446 , n4294 , n4445 );
and ( n4447 , n3985 , n3989 );
and ( n4448 , n3989 , n4138 );
and ( n4449 , n3985 , n4138 );
or ( n4450 , n4447 , n4448 , n4449 );
xor ( n4451 , n4446 , n4450 );
and ( n4452 , n4139 , n4143 );
and ( n4453 , n4144 , n4147 );
or ( n4454 , n4452 , n4453 );
xor ( n4455 , n4451 , n4454 );
buf ( n4456 , n4455 );
buf ( n4457 , n4456 );
not ( n4458 , n4457 );
buf ( n4459 , n523 );
not ( n4460 , n4459 );
nor ( n4461 , n4458 , n4460 );
xor ( n4462 , n4288 , n4461 );
xor ( n4463 , n4159 , n4285 );
nor ( n4464 , n4151 , n4460 );
and ( n4465 , n4463 , n4464 );
xor ( n4466 , n4463 , n4464 );
xor ( n4467 , n4163 , n4283 );
nor ( n4468 , n3853 , n4460 );
and ( n4469 , n4467 , n4468 );
xor ( n4470 , n4467 , n4468 );
xor ( n4471 , n4167 , n4281 );
nor ( n4472 , n3570 , n4460 );
and ( n4473 , n4471 , n4472 );
xor ( n4474 , n4471 , n4472 );
xor ( n4475 , n4171 , n4279 );
nor ( n4476 , n3300 , n4460 );
and ( n4477 , n4475 , n4476 );
xor ( n4478 , n4475 , n4476 );
xor ( n4479 , n4175 , n4277 );
nor ( n4480 , n3043 , n4460 );
and ( n4481 , n4479 , n4480 );
xor ( n4482 , n4479 , n4480 );
xor ( n4483 , n4179 , n4275 );
nor ( n4484 , n2797 , n4460 );
and ( n4485 , n4483 , n4484 );
xor ( n4486 , n4483 , n4484 );
xor ( n4487 , n4183 , n4273 );
nor ( n4488 , n2566 , n4460 );
and ( n4489 , n4487 , n4488 );
xor ( n4490 , n4487 , n4488 );
xor ( n4491 , n4187 , n4271 );
nor ( n4492 , n2343 , n4460 );
and ( n4493 , n4491 , n4492 );
xor ( n4494 , n4491 , n4492 );
xor ( n4495 , n4191 , n4269 );
nor ( n4496 , n2137 , n4460 );
and ( n4497 , n4495 , n4496 );
xor ( n4498 , n4495 , n4496 );
xor ( n4499 , n4195 , n4267 );
nor ( n4500 , n1945 , n4460 );
and ( n4501 , n4499 , n4500 );
xor ( n4502 , n4499 , n4500 );
xor ( n4503 , n4199 , n4265 );
nor ( n4504 , n1766 , n4460 );
and ( n4505 , n4503 , n4504 );
xor ( n4506 , n4503 , n4504 );
xor ( n4507 , n4203 , n4263 );
nor ( n4508 , n1598 , n4460 );
and ( n4509 , n4507 , n4508 );
xor ( n4510 , n4507 , n4508 );
xor ( n4511 , n4207 , n4261 );
nor ( n4512 , n1445 , n4460 );
and ( n4513 , n4511 , n4512 );
xor ( n4514 , n4511 , n4512 );
xor ( n4515 , n4211 , n4259 );
nor ( n4516 , n1303 , n4460 );
and ( n4517 , n4515 , n4516 );
xor ( n4518 , n4515 , n4516 );
xor ( n4519 , n4215 , n4257 );
nor ( n4520 , n1176 , n4460 );
and ( n4521 , n4519 , n4520 );
xor ( n4522 , n4519 , n4520 );
xor ( n4523 , n4219 , n4255 );
nor ( n4524 , n1062 , n4460 );
and ( n4525 , n4523 , n4524 );
xor ( n4526 , n4523 , n4524 );
xor ( n4527 , n4223 , n4253 );
nor ( n4528 , n958 , n4460 );
and ( n4529 , n4527 , n4528 );
xor ( n4530 , n4527 , n4528 );
xor ( n4531 , n4227 , n4251 );
nor ( n4532 , n868 , n4460 );
and ( n4533 , n4531 , n4532 );
xor ( n4534 , n4531 , n4532 );
xor ( n4535 , n4231 , n4249 );
nor ( n4536 , n796 , n4460 );
and ( n4537 , n4535 , n4536 );
xor ( n4538 , n4535 , n4536 );
xor ( n4539 , n4235 , n4247 );
nor ( n4540 , n733 , n4460 );
and ( n4541 , n4539 , n4540 );
xor ( n4542 , n4539 , n4540 );
xor ( n4543 , n4240 , n4245 );
nor ( n4544 , n684 , n4460 );
and ( n4545 , n4543 , n4544 );
xor ( n4546 , n4543 , n4544 );
xor ( n4547 , n4242 , n4243 );
buf ( n4548 , n4547 );
nor ( n4549 , n646 , n4460 );
and ( n4550 , n4548 , n4549 );
xor ( n4551 , n4548 , n4549 );
nor ( n4552 , n601 , n3855 );
buf ( n4553 , n4552 );
nor ( n4554 , n622 , n4460 );
and ( n4555 , n4553 , n4554 );
buf ( n4556 , n4555 );
and ( n4557 , n4551 , n4556 );
or ( n4558 , n4550 , n4557 );
and ( n4559 , n4546 , n4558 );
or ( n4560 , n4545 , n4559 );
and ( n4561 , n4542 , n4560 );
or ( n4562 , n4541 , n4561 );
and ( n4563 , n4538 , n4562 );
or ( n4564 , n4537 , n4563 );
and ( n4565 , n4534 , n4564 );
or ( n4566 , n4533 , n4565 );
and ( n4567 , n4530 , n4566 );
or ( n4568 , n4529 , n4567 );
and ( n4569 , n4526 , n4568 );
or ( n4570 , n4525 , n4569 );
and ( n4571 , n4522 , n4570 );
or ( n4572 , n4521 , n4571 );
and ( n4573 , n4518 , n4572 );
or ( n4574 , n4517 , n4573 );
and ( n4575 , n4514 , n4574 );
or ( n4576 , n4513 , n4575 );
and ( n4577 , n4510 , n4576 );
or ( n4578 , n4509 , n4577 );
and ( n4579 , n4506 , n4578 );
or ( n4580 , n4505 , n4579 );
and ( n4581 , n4502 , n4580 );
or ( n4582 , n4501 , n4581 );
and ( n4583 , n4498 , n4582 );
or ( n4584 , n4497 , n4583 );
and ( n4585 , n4494 , n4584 );
or ( n4586 , n4493 , n4585 );
and ( n4587 , n4490 , n4586 );
or ( n4588 , n4489 , n4587 );
and ( n4589 , n4486 , n4588 );
or ( n4590 , n4485 , n4589 );
and ( n4591 , n4482 , n4590 );
or ( n4592 , n4481 , n4591 );
and ( n4593 , n4478 , n4592 );
or ( n4594 , n4477 , n4593 );
and ( n4595 , n4474 , n4594 );
or ( n4596 , n4473 , n4595 );
and ( n4597 , n4470 , n4596 );
or ( n4598 , n4469 , n4597 );
and ( n4599 , n4466 , n4598 );
or ( n4600 , n4465 , n4599 );
xor ( n4601 , n4462 , n4600 );
and ( n4602 , n4423 , n4424 );
and ( n4603 , n4424 , n4443 );
and ( n4604 , n4423 , n4443 );
or ( n4605 , n4602 , n4603 , n4604 );
and ( n4606 , n4298 , n4418 );
and ( n4607 , n4418 , n4444 );
and ( n4608 , n4298 , n4444 );
or ( n4609 , n4606 , n4607 , n4608 );
xor ( n4610 , n4605 , n4609 );
and ( n4611 , n4302 , n4349 );
and ( n4612 , n4349 , n4417 );
and ( n4613 , n4302 , n4417 );
or ( n4614 , n4611 , n4612 , n4613 );
and ( n4615 , n4354 , n4377 );
and ( n4616 , n4377 , n4416 );
and ( n4617 , n4354 , n4416 );
or ( n4618 , n4615 , n4616 , n4617 );
and ( n4619 , n4315 , n4331 );
and ( n4620 , n4331 , n4347 );
and ( n4621 , n4315 , n4347 );
or ( n4622 , n4619 , n4620 , n4621 );
and ( n4623 , n4358 , n4362 );
and ( n4624 , n4362 , n4376 );
and ( n4625 , n4358 , n4376 );
or ( n4626 , n4623 , n4624 , n4625 );
xor ( n4627 , n4622 , n4626 );
and ( n4628 , n4336 , n4340 );
and ( n4629 , n4340 , n4346 );
and ( n4630 , n4336 , n4346 );
or ( n4631 , n4628 , n4629 , n4630 );
and ( n4632 , n4326 , n4327 );
and ( n4633 , n4327 , n4329 );
and ( n4634 , n4326 , n4329 );
or ( n4635 , n4632 , n4633 , n4634 );
and ( n4636 , n3182 , n719 );
and ( n4637 , n3545 , n663 );
xor ( n4638 , n4636 , n4637 );
and ( n4639 , n3801 , n635 );
xor ( n4640 , n4638 , n4639 );
xor ( n4641 , n4635 , n4640 );
and ( n4642 , n2462 , n940 );
and ( n4643 , n2779 , n840 );
xor ( n4644 , n4642 , n4643 );
and ( n4645 , n3024 , n771 );
xor ( n4646 , n4644 , n4645 );
xor ( n4647 , n4641 , n4646 );
xor ( n4648 , n4631 , n4647 );
and ( n4649 , n4342 , n4343 );
and ( n4650 , n4343 , n4345 );
and ( n4651 , n4342 , n4345 );
or ( n4652 , n4649 , n4650 , n4651 );
and ( n4653 , n1383 , n1551 );
and ( n4654 , n1580 , n1424 );
and ( n4655 , n4653 , n4654 );
and ( n4656 , n4654 , n4374 );
and ( n4657 , n4653 , n4374 );
or ( n4658 , n4655 , n4656 , n4657 );
xor ( n4659 , n4652 , n4658 );
and ( n4660 , n1933 , n1254 );
and ( n4661 , n2120 , n1134 );
xor ( n4662 , n4660 , n4661 );
and ( n4663 , n2324 , n1034 );
xor ( n4664 , n4662 , n4663 );
xor ( n4665 , n4659 , n4664 );
xor ( n4666 , n4648 , n4665 );
xor ( n4667 , n4627 , n4666 );
xor ( n4668 , n4618 , n4667 );
and ( n4669 , n4382 , n4397 );
and ( n4670 , n4397 , n4415 );
and ( n4671 , n4382 , n4415 );
or ( n4672 , n4669 , n4670 , n4671 );
and ( n4673 , n4367 , n4372 );
and ( n4674 , n4372 , n4375 );
and ( n4675 , n4367 , n4375 );
or ( n4676 , n4673 , n4674 , n4675 );
and ( n4677 , n4386 , n4390 );
and ( n4678 , n4390 , n4396 );
and ( n4679 , n4386 , n4396 );
or ( n4680 , n4677 , n4678 , n4679 );
xor ( n4681 , n4676 , n4680 );
and ( n4682 , n4368 , n4369 );
and ( n4683 , n4369 , n4371 );
and ( n4684 , n4368 , n4371 );
or ( n4685 , n4682 , n4683 , n4684 );
and ( n4686 , n1383 , n1738 );
buf ( n4687 , n1580 );
xor ( n4688 , n4686 , n4687 );
and ( n4689 , n1694 , n1424 );
xor ( n4690 , n4688 , n4689 );
xor ( n4691 , n4685 , n4690 );
and ( n4692 , n1047 , n2298 );
and ( n4693 , n1164 , n2100 );
xor ( n4694 , n4692 , n4693 );
and ( n4695 , n1287 , n1882 );
xor ( n4696 , n4694 , n4695 );
xor ( n4697 , n4691 , n4696 );
xor ( n4698 , n4681 , n4697 );
xor ( n4699 , n4672 , n4698 );
and ( n4700 , n4402 , n4408 );
and ( n4701 , n4408 , n4414 );
and ( n4702 , n4402 , n4414 );
or ( n4703 , n4700 , n4701 , n4702 );
and ( n4704 , n4410 , n4411 );
and ( n4705 , n4411 , n4413 );
and ( n4706 , n4410 , n4413 );
or ( n4707 , n4704 , n4705 , n4706 );
and ( n4708 , n4392 , n4393 );
and ( n4709 , n4393 , n4395 );
and ( n4710 , n4392 , n4395 );
or ( n4711 , n4708 , n4709 , n4710 );
xor ( n4712 , n4707 , n4711 );
and ( n4713 , n783 , n2981 );
and ( n4714 , n856 , n2739 );
xor ( n4715 , n4713 , n4714 );
and ( n4716 , n925 , n2544 );
xor ( n4717 , n4715 , n4716 );
xor ( n4718 , n4712 , n4717 );
xor ( n4719 , n4703 , n4718 );
and ( n4720 , n4404 , n4405 );
and ( n4721 , n4405 , n4407 );
and ( n4722 , n4404 , n4407 );
or ( n4723 , n4720 , n4721 , n4722 );
and ( n4724 , n632 , n3749 );
and ( n4725 , n671 , n3495 );
xor ( n4726 , n4724 , n4725 );
and ( n4727 , n715 , n3271 );
xor ( n4728 , n4726 , n4727 );
xor ( n4729 , n4723 , n4728 );
buf ( n4730 , n444 );
and ( n4731 , n599 , n4730 );
and ( n4732 , n608 , n4403 );
xor ( n4733 , n4731 , n4732 );
and ( n4734 , n611 , n4102 );
xor ( n4735 , n4733 , n4734 );
xor ( n4736 , n4729 , n4735 );
xor ( n4737 , n4719 , n4736 );
xor ( n4738 , n4699 , n4737 );
xor ( n4739 , n4668 , n4738 );
xor ( n4740 , n4614 , n4739 );
and ( n4741 , n4306 , n4310 );
and ( n4742 , n4310 , n4348 );
and ( n4743 , n4306 , n4348 );
or ( n4744 , n4741 , n4742 , n4743 );
and ( n4745 , n4426 , n4442 );
xor ( n4746 , n4744 , n4745 );
and ( n4747 , n4430 , n4431 );
and ( n4748 , n4431 , n4441 );
and ( n4749 , n4430 , n4441 );
or ( n4750 , n4747 , n4748 , n4749 );
and ( n4751 , n4319 , n4324 );
and ( n4752 , n4324 , n4330 );
and ( n4753 , n4319 , n4330 );
or ( n4754 , n4751 , n4752 , n4753 );
and ( n4755 , n4436 , n4440 );
xor ( n4756 , n4754 , n4755 );
and ( n4757 , n4320 , n4321 );
and ( n4758 , n4321 , n4323 );
and ( n4759 , n4320 , n4323 );
or ( n4760 , n4757 , n4758 , n4759 );
and ( n4761 , n4437 , n4439 );
xor ( n4762 , n4760 , n4761 );
and ( n4763 , n4132 , n606 );
and ( n4764 , n4438 , n615 );
xor ( n4765 , n4763 , n4764 );
buf ( n4766 , n444 );
and ( n4767 , n4766 , n612 );
xor ( n4768 , n4765 , n4767 );
xor ( n4769 , n4762 , n4768 );
xor ( n4770 , n4756 , n4769 );
xor ( n4771 , n4750 , n4770 );
xor ( n4772 , n4746 , n4771 );
xor ( n4773 , n4740 , n4772 );
xor ( n4774 , n4610 , n4773 );
and ( n4775 , n4289 , n4293 );
and ( n4776 , n4293 , n4445 );
and ( n4777 , n4289 , n4445 );
or ( n4778 , n4775 , n4776 , n4777 );
xor ( n4779 , n4774 , n4778 );
and ( n4780 , n4446 , n4450 );
and ( n4781 , n4451 , n4454 );
or ( n4782 , n4780 , n4781 );
xor ( n4783 , n4779 , n4782 );
buf ( n4784 , n4783 );
buf ( n4785 , n4784 );
not ( n4786 , n4785 );
buf ( n4787 , n524 );
not ( n4788 , n4787 );
nor ( n4789 , n4786 , n4788 );
xor ( n4790 , n4601 , n4789 );
xor ( n4791 , n4466 , n4598 );
nor ( n4792 , n4458 , n4788 );
and ( n4793 , n4791 , n4792 );
xor ( n4794 , n4791 , n4792 );
xor ( n4795 , n4470 , n4596 );
nor ( n4796 , n4151 , n4788 );
and ( n4797 , n4795 , n4796 );
xor ( n4798 , n4795 , n4796 );
xor ( n4799 , n4474 , n4594 );
nor ( n4800 , n3853 , n4788 );
and ( n4801 , n4799 , n4800 );
xor ( n4802 , n4799 , n4800 );
xor ( n4803 , n4478 , n4592 );
nor ( n4804 , n3570 , n4788 );
and ( n4805 , n4803 , n4804 );
xor ( n4806 , n4803 , n4804 );
xor ( n4807 , n4482 , n4590 );
nor ( n4808 , n3300 , n4788 );
and ( n4809 , n4807 , n4808 );
xor ( n4810 , n4807 , n4808 );
xor ( n4811 , n4486 , n4588 );
nor ( n4812 , n3043 , n4788 );
and ( n4813 , n4811 , n4812 );
xor ( n4814 , n4811 , n4812 );
xor ( n4815 , n4490 , n4586 );
nor ( n4816 , n2797 , n4788 );
and ( n4817 , n4815 , n4816 );
xor ( n4818 , n4815 , n4816 );
xor ( n4819 , n4494 , n4584 );
nor ( n4820 , n2566 , n4788 );
and ( n4821 , n4819 , n4820 );
xor ( n4822 , n4819 , n4820 );
xor ( n4823 , n4498 , n4582 );
nor ( n4824 , n2343 , n4788 );
and ( n4825 , n4823 , n4824 );
xor ( n4826 , n4823 , n4824 );
xor ( n4827 , n4502 , n4580 );
nor ( n4828 , n2137 , n4788 );
and ( n4829 , n4827 , n4828 );
xor ( n4830 , n4827 , n4828 );
xor ( n4831 , n4506 , n4578 );
nor ( n4832 , n1945 , n4788 );
and ( n4833 , n4831 , n4832 );
xor ( n4834 , n4831 , n4832 );
xor ( n4835 , n4510 , n4576 );
nor ( n4836 , n1766 , n4788 );
and ( n4837 , n4835 , n4836 );
xor ( n4838 , n4835 , n4836 );
xor ( n4839 , n4514 , n4574 );
nor ( n4840 , n1598 , n4788 );
and ( n4841 , n4839 , n4840 );
xor ( n4842 , n4839 , n4840 );
xor ( n4843 , n4518 , n4572 );
nor ( n4844 , n1445 , n4788 );
and ( n4845 , n4843 , n4844 );
xor ( n4846 , n4843 , n4844 );
xor ( n4847 , n4522 , n4570 );
nor ( n4848 , n1303 , n4788 );
and ( n4849 , n4847 , n4848 );
xor ( n4850 , n4847 , n4848 );
xor ( n4851 , n4526 , n4568 );
nor ( n4852 , n1176 , n4788 );
and ( n4853 , n4851 , n4852 );
xor ( n4854 , n4851 , n4852 );
xor ( n4855 , n4530 , n4566 );
nor ( n4856 , n1062 , n4788 );
and ( n4857 , n4855 , n4856 );
xor ( n4858 , n4855 , n4856 );
xor ( n4859 , n4534 , n4564 );
nor ( n4860 , n958 , n4788 );
and ( n4861 , n4859 , n4860 );
xor ( n4862 , n4859 , n4860 );
xor ( n4863 , n4538 , n4562 );
nor ( n4864 , n868 , n4788 );
and ( n4865 , n4863 , n4864 );
xor ( n4866 , n4863 , n4864 );
xor ( n4867 , n4542 , n4560 );
nor ( n4868 , n796 , n4788 );
and ( n4869 , n4867 , n4868 );
xor ( n4870 , n4867 , n4868 );
xor ( n4871 , n4546 , n4558 );
nor ( n4872 , n733 , n4788 );
and ( n4873 , n4871 , n4872 );
xor ( n4874 , n4871 , n4872 );
xor ( n4875 , n4551 , n4556 );
nor ( n4876 , n684 , n4788 );
and ( n4877 , n4875 , n4876 );
xor ( n4878 , n4875 , n4876 );
xor ( n4879 , n4553 , n4554 );
buf ( n4880 , n4879 );
nor ( n4881 , n646 , n4788 );
and ( n4882 , n4880 , n4881 );
xor ( n4883 , n4880 , n4881 );
nor ( n4884 , n601 , n4153 );
buf ( n4885 , n4884 );
nor ( n4886 , n622 , n4788 );
and ( n4887 , n4885 , n4886 );
buf ( n4888 , n4887 );
and ( n4889 , n4883 , n4888 );
or ( n4890 , n4882 , n4889 );
and ( n4891 , n4878 , n4890 );
or ( n4892 , n4877 , n4891 );
and ( n4893 , n4874 , n4892 );
or ( n4894 , n4873 , n4893 );
and ( n4895 , n4870 , n4894 );
or ( n4896 , n4869 , n4895 );
and ( n4897 , n4866 , n4896 );
or ( n4898 , n4865 , n4897 );
and ( n4899 , n4862 , n4898 );
or ( n4900 , n4861 , n4899 );
and ( n4901 , n4858 , n4900 );
or ( n4902 , n4857 , n4901 );
and ( n4903 , n4854 , n4902 );
or ( n4904 , n4853 , n4903 );
and ( n4905 , n4850 , n4904 );
or ( n4906 , n4849 , n4905 );
and ( n4907 , n4846 , n4906 );
or ( n4908 , n4845 , n4907 );
and ( n4909 , n4842 , n4908 );
or ( n4910 , n4841 , n4909 );
and ( n4911 , n4838 , n4910 );
or ( n4912 , n4837 , n4911 );
and ( n4913 , n4834 , n4912 );
or ( n4914 , n4833 , n4913 );
and ( n4915 , n4830 , n4914 );
or ( n4916 , n4829 , n4915 );
and ( n4917 , n4826 , n4916 );
or ( n4918 , n4825 , n4917 );
and ( n4919 , n4822 , n4918 );
or ( n4920 , n4821 , n4919 );
and ( n4921 , n4818 , n4920 );
or ( n4922 , n4817 , n4921 );
and ( n4923 , n4814 , n4922 );
or ( n4924 , n4813 , n4923 );
and ( n4925 , n4810 , n4924 );
or ( n4926 , n4809 , n4925 );
and ( n4927 , n4806 , n4926 );
or ( n4928 , n4805 , n4927 );
and ( n4929 , n4802 , n4928 );
or ( n4930 , n4801 , n4929 );
and ( n4931 , n4798 , n4930 );
or ( n4932 , n4797 , n4931 );
and ( n4933 , n4794 , n4932 );
or ( n4934 , n4793 , n4933 );
xor ( n4935 , n4790 , n4934 );
and ( n4936 , n4744 , n4745 );
and ( n4937 , n4745 , n4771 );
and ( n4938 , n4744 , n4771 );
or ( n4939 , n4936 , n4937 , n4938 );
and ( n4940 , n4614 , n4739 );
and ( n4941 , n4739 , n4772 );
and ( n4942 , n4614 , n4772 );
or ( n4943 , n4940 , n4941 , n4942 );
xor ( n4944 , n4939 , n4943 );
and ( n4945 , n4618 , n4667 );
and ( n4946 , n4667 , n4738 );
and ( n4947 , n4618 , n4738 );
or ( n4948 , n4945 , n4946 , n4947 );
and ( n4949 , n4622 , n4626 );
and ( n4950 , n4626 , n4666 );
and ( n4951 , n4622 , n4666 );
or ( n4952 , n4949 , n4950 , n4951 );
and ( n4953 , n4750 , n4770 );
xor ( n4954 , n4952 , n4953 );
and ( n4955 , n4754 , n4755 );
and ( n4956 , n4755 , n4769 );
and ( n4957 , n4754 , n4769 );
or ( n4958 , n4955 , n4956 , n4957 );
buf ( n4959 , n443 );
and ( n4960 , n4959 , n612 );
xor ( n4961 , n4958 , n4960 );
and ( n4962 , n4760 , n4761 );
and ( n4963 , n4761 , n4768 );
and ( n4964 , n4760 , n4768 );
or ( n4965 , n4962 , n4963 , n4964 );
and ( n4966 , n4635 , n4640 );
and ( n4967 , n4640 , n4646 );
and ( n4968 , n4635 , n4646 );
or ( n4969 , n4966 , n4967 , n4968 );
xor ( n4970 , n4965 , n4969 );
and ( n4971 , n4763 , n4764 );
and ( n4972 , n4764 , n4767 );
and ( n4973 , n4763 , n4767 );
or ( n4974 , n4971 , n4972 , n4973 );
and ( n4975 , n4636 , n4637 );
and ( n4976 , n4637 , n4639 );
and ( n4977 , n4636 , n4639 );
or ( n4978 , n4975 , n4976 , n4977 );
xor ( n4979 , n4974 , n4978 );
and ( n4980 , n4132 , n635 );
and ( n4981 , n4438 , n606 );
xor ( n4982 , n4980 , n4981 );
and ( n4983 , n4766 , n615 );
xor ( n4984 , n4982 , n4983 );
xor ( n4985 , n4979 , n4984 );
xor ( n4986 , n4970 , n4985 );
xor ( n4987 , n4961 , n4986 );
xor ( n4988 , n4954 , n4987 );
xor ( n4989 , n4948 , n4988 );
and ( n4990 , n4672 , n4698 );
and ( n4991 , n4698 , n4737 );
and ( n4992 , n4672 , n4737 );
or ( n4993 , n4990 , n4991 , n4992 );
and ( n4994 , n4631 , n4647 );
and ( n4995 , n4647 , n4665 );
and ( n4996 , n4631 , n4665 );
or ( n4997 , n4994 , n4995 , n4996 );
and ( n4998 , n4676 , n4680 );
and ( n4999 , n4680 , n4697 );
and ( n5000 , n4676 , n4697 );
or ( n5001 , n4998 , n4999 , n5000 );
xor ( n5002 , n4997 , n5001 );
and ( n5003 , n4652 , n4658 );
and ( n5004 , n4658 , n4664 );
and ( n5005 , n4652 , n4664 );
or ( n5006 , n5003 , n5004 , n5005 );
and ( n5007 , n4642 , n4643 );
and ( n5008 , n4643 , n4645 );
and ( n5009 , n4642 , n4645 );
or ( n5010 , n5007 , n5008 , n5009 );
and ( n5011 , n3182 , n771 );
and ( n5012 , n3545 , n719 );
xor ( n5013 , n5011 , n5012 );
and ( n5014 , n3801 , n663 );
xor ( n5015 , n5013 , n5014 );
xor ( n5016 , n5010 , n5015 );
and ( n5017 , n2462 , n1034 );
and ( n5018 , n2779 , n940 );
xor ( n5019 , n5017 , n5018 );
and ( n5020 , n3024 , n840 );
xor ( n5021 , n5019 , n5020 );
xor ( n5022 , n5016 , n5021 );
xor ( n5023 , n5006 , n5022 );
and ( n5024 , n4660 , n4661 );
and ( n5025 , n4661 , n4663 );
and ( n5026 , n4660 , n4663 );
or ( n5027 , n5024 , n5025 , n5026 );
and ( n5028 , n4686 , n4687 );
and ( n5029 , n4687 , n4689 );
and ( n5030 , n4686 , n4689 );
or ( n5031 , n5028 , n5029 , n5030 );
xor ( n5032 , n5027 , n5031 );
and ( n5033 , n1933 , n1424 );
and ( n5034 , n2120 , n1254 );
xor ( n5035 , n5033 , n5034 );
and ( n5036 , n2324 , n1134 );
xor ( n5037 , n5035 , n5036 );
xor ( n5038 , n5032 , n5037 );
xor ( n5039 , n5023 , n5038 );
xor ( n5040 , n5002 , n5039 );
xor ( n5041 , n4993 , n5040 );
and ( n5042 , n4703 , n4718 );
and ( n5043 , n4718 , n4736 );
and ( n5044 , n4703 , n4736 );
or ( n5045 , n5042 , n5043 , n5044 );
and ( n5046 , n4685 , n4690 );
and ( n5047 , n4690 , n4696 );
and ( n5048 , n4685 , n4696 );
or ( n5049 , n5046 , n5047 , n5048 );
and ( n5050 , n4707 , n4711 );
and ( n5051 , n4711 , n4717 );
and ( n5052 , n4707 , n4717 );
or ( n5053 , n5050 , n5051 , n5052 );
xor ( n5054 , n5049 , n5053 );
and ( n5055 , n4692 , n4693 );
and ( n5056 , n4693 , n4695 );
and ( n5057 , n4692 , n4695 );
or ( n5058 , n5055 , n5056 , n5057 );
and ( n5059 , n1383 , n1882 );
and ( n5060 , n1580 , n1738 );
xor ( n5061 , n5059 , n5060 );
and ( n5062 , n1694 , n1551 );
xor ( n5063 , n5061 , n5062 );
xor ( n5064 , n5058 , n5063 );
and ( n5065 , n1047 , n2544 );
and ( n5066 , n1164 , n2298 );
xor ( n5067 , n5065 , n5066 );
and ( n5068 , n1287 , n2100 );
xor ( n5069 , n5067 , n5068 );
xor ( n5070 , n5064 , n5069 );
xor ( n5071 , n5054 , n5070 );
xor ( n5072 , n5045 , n5071 );
and ( n5073 , n4723 , n4728 );
and ( n5074 , n4728 , n4735 );
and ( n5075 , n4723 , n4735 );
or ( n5076 , n5073 , n5074 , n5075 );
and ( n5077 , n4713 , n4714 );
and ( n5078 , n4714 , n4716 );
and ( n5079 , n4713 , n4716 );
or ( n5080 , n5077 , n5078 , n5079 );
and ( n5081 , n4724 , n4725 );
and ( n5082 , n4725 , n4727 );
and ( n5083 , n4724 , n4727 );
or ( n5084 , n5081 , n5082 , n5083 );
xor ( n5085 , n5080 , n5084 );
and ( n5086 , n783 , n3271 );
and ( n5087 , n856 , n2981 );
xor ( n5088 , n5086 , n5087 );
and ( n5089 , n925 , n2739 );
xor ( n5090 , n5088 , n5089 );
xor ( n5091 , n5085 , n5090 );
xor ( n5092 , n5076 , n5091 );
and ( n5093 , n4731 , n4732 );
and ( n5094 , n4732 , n4734 );
and ( n5095 , n4731 , n4734 );
or ( n5096 , n5093 , n5094 , n5095 );
and ( n5097 , n632 , n4102 );
and ( n5098 , n671 , n3749 );
xor ( n5099 , n5097 , n5098 );
and ( n5100 , n715 , n3495 );
xor ( n5101 , n5099 , n5100 );
xor ( n5102 , n5096 , n5101 );
buf ( n5103 , n443 );
and ( n5104 , n599 , n5103 );
and ( n5105 , n608 , n4730 );
xor ( n5106 , n5104 , n5105 );
and ( n5107 , n611 , n4403 );
xor ( n5108 , n5106 , n5107 );
xor ( n5109 , n5102 , n5108 );
xor ( n5110 , n5092 , n5109 );
xor ( n5111 , n5072 , n5110 );
xor ( n5112 , n5041 , n5111 );
xor ( n5113 , n4989 , n5112 );
xor ( n5114 , n4944 , n5113 );
and ( n5115 , n4605 , n4609 );
and ( n5116 , n4609 , n4773 );
and ( n5117 , n4605 , n4773 );
or ( n5118 , n5115 , n5116 , n5117 );
xor ( n5119 , n5114 , n5118 );
and ( n5120 , n4774 , n4778 );
and ( n5121 , n4779 , n4782 );
or ( n5122 , n5120 , n5121 );
xor ( n5123 , n5119 , n5122 );
buf ( n5124 , n5123 );
buf ( n5125 , n5124 );
not ( n5126 , n5125 );
buf ( n5127 , n525 );
not ( n5128 , n5127 );
nor ( n5129 , n5126 , n5128 );
xor ( n5130 , n4935 , n5129 );
xor ( n5131 , n4794 , n4932 );
nor ( n5132 , n4786 , n5128 );
and ( n5133 , n5131 , n5132 );
xor ( n5134 , n5131 , n5132 );
xor ( n5135 , n4798 , n4930 );
nor ( n5136 , n4458 , n5128 );
and ( n5137 , n5135 , n5136 );
xor ( n5138 , n5135 , n5136 );
xor ( n5139 , n4802 , n4928 );
nor ( n5140 , n4151 , n5128 );
and ( n5141 , n5139 , n5140 );
xor ( n5142 , n5139 , n5140 );
xor ( n5143 , n4806 , n4926 );
nor ( n5144 , n3853 , n5128 );
and ( n5145 , n5143 , n5144 );
xor ( n5146 , n5143 , n5144 );
xor ( n5147 , n4810 , n4924 );
nor ( n5148 , n3570 , n5128 );
and ( n5149 , n5147 , n5148 );
xor ( n5150 , n5147 , n5148 );
xor ( n5151 , n4814 , n4922 );
nor ( n5152 , n3300 , n5128 );
and ( n5153 , n5151 , n5152 );
xor ( n5154 , n5151 , n5152 );
xor ( n5155 , n4818 , n4920 );
nor ( n5156 , n3043 , n5128 );
and ( n5157 , n5155 , n5156 );
xor ( n5158 , n5155 , n5156 );
xor ( n5159 , n4822 , n4918 );
nor ( n5160 , n2797 , n5128 );
and ( n5161 , n5159 , n5160 );
xor ( n5162 , n5159 , n5160 );
xor ( n5163 , n4826 , n4916 );
nor ( n5164 , n2566 , n5128 );
and ( n5165 , n5163 , n5164 );
xor ( n5166 , n5163 , n5164 );
xor ( n5167 , n4830 , n4914 );
nor ( n5168 , n2343 , n5128 );
and ( n5169 , n5167 , n5168 );
xor ( n5170 , n5167 , n5168 );
xor ( n5171 , n4834 , n4912 );
nor ( n5172 , n2137 , n5128 );
and ( n5173 , n5171 , n5172 );
xor ( n5174 , n5171 , n5172 );
xor ( n5175 , n4838 , n4910 );
nor ( n5176 , n1945 , n5128 );
and ( n5177 , n5175 , n5176 );
xor ( n5178 , n5175 , n5176 );
xor ( n5179 , n4842 , n4908 );
nor ( n5180 , n1766 , n5128 );
and ( n5181 , n5179 , n5180 );
xor ( n5182 , n5179 , n5180 );
xor ( n5183 , n4846 , n4906 );
nor ( n5184 , n1598 , n5128 );
and ( n5185 , n5183 , n5184 );
xor ( n5186 , n5183 , n5184 );
xor ( n5187 , n4850 , n4904 );
nor ( n5188 , n1445 , n5128 );
and ( n5189 , n5187 , n5188 );
xor ( n5190 , n5187 , n5188 );
xor ( n5191 , n4854 , n4902 );
nor ( n5192 , n1303 , n5128 );
and ( n5193 , n5191 , n5192 );
xor ( n5194 , n5191 , n5192 );
xor ( n5195 , n4858 , n4900 );
nor ( n5196 , n1176 , n5128 );
and ( n5197 , n5195 , n5196 );
xor ( n5198 , n5195 , n5196 );
xor ( n5199 , n4862 , n4898 );
nor ( n5200 , n1062 , n5128 );
and ( n5201 , n5199 , n5200 );
xor ( n5202 , n5199 , n5200 );
xor ( n5203 , n4866 , n4896 );
nor ( n5204 , n958 , n5128 );
and ( n5205 , n5203 , n5204 );
xor ( n5206 , n5203 , n5204 );
xor ( n5207 , n4870 , n4894 );
nor ( n5208 , n868 , n5128 );
and ( n5209 , n5207 , n5208 );
xor ( n5210 , n5207 , n5208 );
xor ( n5211 , n4874 , n4892 );
nor ( n5212 , n796 , n5128 );
and ( n5213 , n5211 , n5212 );
xor ( n5214 , n5211 , n5212 );
xor ( n5215 , n4878 , n4890 );
nor ( n5216 , n733 , n5128 );
and ( n5217 , n5215 , n5216 );
xor ( n5218 , n5215 , n5216 );
xor ( n5219 , n4883 , n4888 );
nor ( n5220 , n684 , n5128 );
and ( n5221 , n5219 , n5220 );
xor ( n5222 , n5219 , n5220 );
xor ( n5223 , n4885 , n4886 );
buf ( n5224 , n5223 );
nor ( n5225 , n646 , n5128 );
and ( n5226 , n5224 , n5225 );
xor ( n5227 , n5224 , n5225 );
nor ( n5228 , n601 , n4460 );
buf ( n5229 , n5228 );
nor ( n5230 , n622 , n5128 );
and ( n5231 , n5229 , n5230 );
buf ( n5232 , n5231 );
and ( n5233 , n5227 , n5232 );
or ( n5234 , n5226 , n5233 );
and ( n5235 , n5222 , n5234 );
or ( n5236 , n5221 , n5235 );
and ( n5237 , n5218 , n5236 );
or ( n5238 , n5217 , n5237 );
and ( n5239 , n5214 , n5238 );
or ( n5240 , n5213 , n5239 );
and ( n5241 , n5210 , n5240 );
or ( n5242 , n5209 , n5241 );
and ( n5243 , n5206 , n5242 );
or ( n5244 , n5205 , n5243 );
and ( n5245 , n5202 , n5244 );
or ( n5246 , n5201 , n5245 );
and ( n5247 , n5198 , n5246 );
or ( n5248 , n5197 , n5247 );
and ( n5249 , n5194 , n5248 );
or ( n5250 , n5193 , n5249 );
and ( n5251 , n5190 , n5250 );
or ( n5252 , n5189 , n5251 );
and ( n5253 , n5186 , n5252 );
or ( n5254 , n5185 , n5253 );
and ( n5255 , n5182 , n5254 );
or ( n5256 , n5181 , n5255 );
and ( n5257 , n5178 , n5256 );
or ( n5258 , n5177 , n5257 );
and ( n5259 , n5174 , n5258 );
or ( n5260 , n5173 , n5259 );
and ( n5261 , n5170 , n5260 );
or ( n5262 , n5169 , n5261 );
and ( n5263 , n5166 , n5262 );
or ( n5264 , n5165 , n5263 );
and ( n5265 , n5162 , n5264 );
or ( n5266 , n5161 , n5265 );
and ( n5267 , n5158 , n5266 );
or ( n5268 , n5157 , n5267 );
and ( n5269 , n5154 , n5268 );
or ( n5270 , n5153 , n5269 );
and ( n5271 , n5150 , n5270 );
or ( n5272 , n5149 , n5271 );
and ( n5273 , n5146 , n5272 );
or ( n5274 , n5145 , n5273 );
and ( n5275 , n5142 , n5274 );
or ( n5276 , n5141 , n5275 );
and ( n5277 , n5138 , n5276 );
or ( n5278 , n5137 , n5277 );
and ( n5279 , n5134 , n5278 );
or ( n5280 , n5133 , n5279 );
xor ( n5281 , n5130 , n5280 );
and ( n5282 , n4952 , n4953 );
and ( n5283 , n4953 , n4987 );
and ( n5284 , n4952 , n4987 );
or ( n5285 , n5282 , n5283 , n5284 );
and ( n5286 , n4948 , n4988 );
and ( n5287 , n4988 , n5112 );
and ( n5288 , n4948 , n5112 );
or ( n5289 , n5286 , n5287 , n5288 );
xor ( n5290 , n5285 , n5289 );
and ( n5291 , n4993 , n5040 );
and ( n5292 , n5040 , n5111 );
and ( n5293 , n4993 , n5111 );
or ( n5294 , n5291 , n5292 , n5293 );
and ( n5295 , n5045 , n5071 );
and ( n5296 , n5071 , n5110 );
and ( n5297 , n5045 , n5110 );
or ( n5298 , n5295 , n5296 , n5297 );
and ( n5299 , n5006 , n5022 );
and ( n5300 , n5022 , n5038 );
and ( n5301 , n5006 , n5038 );
or ( n5302 , n5299 , n5300 , n5301 );
and ( n5303 , n5049 , n5053 );
and ( n5304 , n5053 , n5070 );
and ( n5305 , n5049 , n5070 );
or ( n5306 , n5303 , n5304 , n5305 );
xor ( n5307 , n5302 , n5306 );
and ( n5308 , n5027 , n5031 );
and ( n5309 , n5031 , n5037 );
and ( n5310 , n5027 , n5037 );
or ( n5311 , n5308 , n5309 , n5310 );
and ( n5312 , n5017 , n5018 );
and ( n5313 , n5018 , n5020 );
and ( n5314 , n5017 , n5020 );
or ( n5315 , n5312 , n5313 , n5314 );
and ( n5316 , n3182 , n840 );
and ( n5317 , n3545 , n771 );
xor ( n5318 , n5316 , n5317 );
and ( n5319 , n3801 , n719 );
xor ( n5320 , n5318 , n5319 );
xor ( n5321 , n5315 , n5320 );
and ( n5322 , n2462 , n1134 );
and ( n5323 , n2779 , n1034 );
xor ( n5324 , n5322 , n5323 );
and ( n5325 , n3024 , n940 );
xor ( n5326 , n5324 , n5325 );
xor ( n5327 , n5321 , n5326 );
xor ( n5328 , n5311 , n5327 );
and ( n5329 , n5033 , n5034 );
and ( n5330 , n5034 , n5036 );
and ( n5331 , n5033 , n5036 );
or ( n5332 , n5329 , n5330 , n5331 );
and ( n5333 , n5059 , n5060 );
and ( n5334 , n5060 , n5062 );
and ( n5335 , n5059 , n5062 );
or ( n5336 , n5333 , n5334 , n5335 );
xor ( n5337 , n5332 , n5336 );
and ( n5338 , n1933 , n1551 );
and ( n5339 , n2120 , n1424 );
xor ( n5340 , n5338 , n5339 );
and ( n5341 , n2324 , n1254 );
xor ( n5342 , n5340 , n5341 );
xor ( n5343 , n5337 , n5342 );
xor ( n5344 , n5328 , n5343 );
xor ( n5345 , n5307 , n5344 );
xor ( n5346 , n5298 , n5345 );
and ( n5347 , n5076 , n5091 );
and ( n5348 , n5091 , n5109 );
and ( n5349 , n5076 , n5109 );
or ( n5350 , n5347 , n5348 , n5349 );
and ( n5351 , n5058 , n5063 );
and ( n5352 , n5063 , n5069 );
and ( n5353 , n5058 , n5069 );
or ( n5354 , n5351 , n5352 , n5353 );
and ( n5355 , n5080 , n5084 );
and ( n5356 , n5084 , n5090 );
and ( n5357 , n5080 , n5090 );
or ( n5358 , n5355 , n5356 , n5357 );
xor ( n5359 , n5354 , n5358 );
and ( n5360 , n5065 , n5066 );
and ( n5361 , n5066 , n5068 );
and ( n5362 , n5065 , n5068 );
or ( n5363 , n5360 , n5361 , n5362 );
and ( n5364 , n1383 , n2100 );
and ( n5365 , n1580 , n1882 );
xor ( n5366 , n5364 , n5365 );
buf ( n5367 , n1694 );
xor ( n5368 , n5366 , n5367 );
xor ( n5369 , n5363 , n5368 );
and ( n5370 , n1047 , n2739 );
and ( n5371 , n1164 , n2544 );
xor ( n5372 , n5370 , n5371 );
and ( n5373 , n1287 , n2298 );
xor ( n5374 , n5372 , n5373 );
xor ( n5375 , n5369 , n5374 );
xor ( n5376 , n5359 , n5375 );
xor ( n5377 , n5350 , n5376 );
and ( n5378 , n5096 , n5101 );
and ( n5379 , n5101 , n5108 );
and ( n5380 , n5096 , n5108 );
or ( n5381 , n5378 , n5379 , n5380 );
and ( n5382 , n5086 , n5087 );
and ( n5383 , n5087 , n5089 );
and ( n5384 , n5086 , n5089 );
or ( n5385 , n5382 , n5383 , n5384 );
and ( n5386 , n5097 , n5098 );
and ( n5387 , n5098 , n5100 );
and ( n5388 , n5097 , n5100 );
or ( n5389 , n5386 , n5387 , n5388 );
xor ( n5390 , n5385 , n5389 );
and ( n5391 , n783 , n3495 );
and ( n5392 , n856 , n3271 );
xor ( n5393 , n5391 , n5392 );
and ( n5394 , n925 , n2981 );
xor ( n5395 , n5393 , n5394 );
xor ( n5396 , n5390 , n5395 );
xor ( n5397 , n5381 , n5396 );
and ( n5398 , n5104 , n5105 );
and ( n5399 , n5105 , n5107 );
and ( n5400 , n5104 , n5107 );
or ( n5401 , n5398 , n5399 , n5400 );
and ( n5402 , n632 , n4403 );
and ( n5403 , n671 , n4102 );
xor ( n5404 , n5402 , n5403 );
and ( n5405 , n715 , n3749 );
xor ( n5406 , n5404 , n5405 );
xor ( n5407 , n5401 , n5406 );
buf ( n5408 , n442 );
and ( n5409 , n599 , n5408 );
and ( n5410 , n608 , n5103 );
xor ( n5411 , n5409 , n5410 );
and ( n5412 , n611 , n4730 );
xor ( n5413 , n5411 , n5412 );
xor ( n5414 , n5407 , n5413 );
xor ( n5415 , n5397 , n5414 );
xor ( n5416 , n5377 , n5415 );
xor ( n5417 , n5346 , n5416 );
xor ( n5418 , n5294 , n5417 );
and ( n5419 , n4958 , n4960 );
and ( n5420 , n4960 , n4986 );
and ( n5421 , n4958 , n4986 );
or ( n5422 , n5419 , n5420 , n5421 );
and ( n5423 , n4997 , n5001 );
and ( n5424 , n5001 , n5039 );
and ( n5425 , n4997 , n5039 );
or ( n5426 , n5423 , n5424 , n5425 );
xor ( n5427 , n5422 , n5426 );
and ( n5428 , n4965 , n4969 );
and ( n5429 , n4969 , n4985 );
and ( n5430 , n4965 , n4985 );
or ( n5431 , n5428 , n5429 , n5430 );
and ( n5432 , n4974 , n4978 );
and ( n5433 , n4978 , n4984 );
and ( n5434 , n4974 , n4984 );
or ( n5435 , n5432 , n5433 , n5434 );
and ( n5436 , n5010 , n5015 );
and ( n5437 , n5015 , n5021 );
and ( n5438 , n5010 , n5021 );
or ( n5439 , n5436 , n5437 , n5438 );
xor ( n5440 , n5435 , n5439 );
and ( n5441 , n4980 , n4981 );
and ( n5442 , n4981 , n4983 );
and ( n5443 , n4980 , n4983 );
or ( n5444 , n5441 , n5442 , n5443 );
and ( n5445 , n5011 , n5012 );
and ( n5446 , n5012 , n5014 );
and ( n5447 , n5011 , n5014 );
or ( n5448 , n5445 , n5446 , n5447 );
xor ( n5449 , n5444 , n5448 );
and ( n5450 , n4132 , n663 );
and ( n5451 , n4438 , n635 );
xor ( n5452 , n5450 , n5451 );
and ( n5453 , n4766 , n606 );
xor ( n5454 , n5452 , n5453 );
xor ( n5455 , n5449 , n5454 );
xor ( n5456 , n5440 , n5455 );
xor ( n5457 , n5431 , n5456 );
and ( n5458 , n4959 , n615 );
buf ( n5459 , n442 );
and ( n5460 , n5459 , n612 );
xor ( n5461 , n5458 , n5460 );
xor ( n5462 , n5457 , n5461 );
xor ( n5463 , n5427 , n5462 );
xor ( n5464 , n5418 , n5463 );
xor ( n5465 , n5290 , n5464 );
and ( n5466 , n4939 , n4943 );
and ( n5467 , n4943 , n5113 );
and ( n5468 , n4939 , n5113 );
or ( n5469 , n5466 , n5467 , n5468 );
xor ( n5470 , n5465 , n5469 );
and ( n5471 , n5114 , n5118 );
and ( n5472 , n5119 , n5122 );
or ( n5473 , n5471 , n5472 );
xor ( n5474 , n5470 , n5473 );
buf ( n5475 , n5474 );
buf ( n5476 , n5475 );
not ( n5477 , n5476 );
buf ( n5478 , n526 );
not ( n5479 , n5478 );
nor ( n5480 , n5477 , n5479 );
xor ( n5481 , n5281 , n5480 );
xor ( n5482 , n5134 , n5278 );
nor ( n5483 , n5126 , n5479 );
and ( n5484 , n5482 , n5483 );
xor ( n5485 , n5482 , n5483 );
xor ( n5486 , n5138 , n5276 );
nor ( n5487 , n4786 , n5479 );
and ( n5488 , n5486 , n5487 );
xor ( n5489 , n5486 , n5487 );
xor ( n5490 , n5142 , n5274 );
nor ( n5491 , n4458 , n5479 );
and ( n5492 , n5490 , n5491 );
xor ( n5493 , n5490 , n5491 );
xor ( n5494 , n5146 , n5272 );
nor ( n5495 , n4151 , n5479 );
and ( n5496 , n5494 , n5495 );
xor ( n5497 , n5494 , n5495 );
xor ( n5498 , n5150 , n5270 );
nor ( n5499 , n3853 , n5479 );
and ( n5500 , n5498 , n5499 );
xor ( n5501 , n5498 , n5499 );
xor ( n5502 , n5154 , n5268 );
nor ( n5503 , n3570 , n5479 );
and ( n5504 , n5502 , n5503 );
xor ( n5505 , n5502 , n5503 );
xor ( n5506 , n5158 , n5266 );
nor ( n5507 , n3300 , n5479 );
and ( n5508 , n5506 , n5507 );
xor ( n5509 , n5506 , n5507 );
xor ( n5510 , n5162 , n5264 );
nor ( n5511 , n3043 , n5479 );
and ( n5512 , n5510 , n5511 );
xor ( n5513 , n5510 , n5511 );
xor ( n5514 , n5166 , n5262 );
nor ( n5515 , n2797 , n5479 );
and ( n5516 , n5514 , n5515 );
xor ( n5517 , n5514 , n5515 );
xor ( n5518 , n5170 , n5260 );
nor ( n5519 , n2566 , n5479 );
and ( n5520 , n5518 , n5519 );
xor ( n5521 , n5518 , n5519 );
xor ( n5522 , n5174 , n5258 );
nor ( n5523 , n2343 , n5479 );
and ( n5524 , n5522 , n5523 );
xor ( n5525 , n5522 , n5523 );
xor ( n5526 , n5178 , n5256 );
nor ( n5527 , n2137 , n5479 );
and ( n5528 , n5526 , n5527 );
xor ( n5529 , n5526 , n5527 );
xor ( n5530 , n5182 , n5254 );
nor ( n5531 , n1945 , n5479 );
and ( n5532 , n5530 , n5531 );
xor ( n5533 , n5530 , n5531 );
xor ( n5534 , n5186 , n5252 );
nor ( n5535 , n1766 , n5479 );
and ( n5536 , n5534 , n5535 );
xor ( n5537 , n5534 , n5535 );
xor ( n5538 , n5190 , n5250 );
nor ( n5539 , n1598 , n5479 );
and ( n5540 , n5538 , n5539 );
xor ( n5541 , n5538 , n5539 );
xor ( n5542 , n5194 , n5248 );
nor ( n5543 , n1445 , n5479 );
and ( n5544 , n5542 , n5543 );
xor ( n5545 , n5542 , n5543 );
xor ( n5546 , n5198 , n5246 );
nor ( n5547 , n1303 , n5479 );
and ( n5548 , n5546 , n5547 );
xor ( n5549 , n5546 , n5547 );
xor ( n5550 , n5202 , n5244 );
nor ( n5551 , n1176 , n5479 );
and ( n5552 , n5550 , n5551 );
xor ( n5553 , n5550 , n5551 );
xor ( n5554 , n5206 , n5242 );
nor ( n5555 , n1062 , n5479 );
and ( n5556 , n5554 , n5555 );
xor ( n5557 , n5554 , n5555 );
xor ( n5558 , n5210 , n5240 );
nor ( n5559 , n958 , n5479 );
and ( n5560 , n5558 , n5559 );
xor ( n5561 , n5558 , n5559 );
xor ( n5562 , n5214 , n5238 );
nor ( n5563 , n868 , n5479 );
and ( n5564 , n5562 , n5563 );
xor ( n5565 , n5562 , n5563 );
xor ( n5566 , n5218 , n5236 );
nor ( n5567 , n796 , n5479 );
and ( n5568 , n5566 , n5567 );
xor ( n5569 , n5566 , n5567 );
xor ( n5570 , n5222 , n5234 );
nor ( n5571 , n733 , n5479 );
and ( n5572 , n5570 , n5571 );
xor ( n5573 , n5570 , n5571 );
xor ( n5574 , n5227 , n5232 );
nor ( n5575 , n684 , n5479 );
and ( n5576 , n5574 , n5575 );
xor ( n5577 , n5574 , n5575 );
xor ( n5578 , n5229 , n5230 );
buf ( n5579 , n5578 );
nor ( n5580 , n646 , n5479 );
and ( n5581 , n5579 , n5580 );
xor ( n5582 , n5579 , n5580 );
nor ( n5583 , n601 , n4788 );
buf ( n5584 , n5583 );
nor ( n5585 , n622 , n5479 );
and ( n5586 , n5584 , n5585 );
buf ( n5587 , n5586 );
and ( n5588 , n5582 , n5587 );
or ( n5589 , n5581 , n5588 );
and ( n5590 , n5577 , n5589 );
or ( n5591 , n5576 , n5590 );
and ( n5592 , n5573 , n5591 );
or ( n5593 , n5572 , n5592 );
and ( n5594 , n5569 , n5593 );
or ( n5595 , n5568 , n5594 );
and ( n5596 , n5565 , n5595 );
or ( n5597 , n5564 , n5596 );
and ( n5598 , n5561 , n5597 );
or ( n5599 , n5560 , n5598 );
and ( n5600 , n5557 , n5599 );
or ( n5601 , n5556 , n5600 );
and ( n5602 , n5553 , n5601 );
or ( n5603 , n5552 , n5602 );
and ( n5604 , n5549 , n5603 );
or ( n5605 , n5548 , n5604 );
and ( n5606 , n5545 , n5605 );
or ( n5607 , n5544 , n5606 );
and ( n5608 , n5541 , n5607 );
or ( n5609 , n5540 , n5608 );
and ( n5610 , n5537 , n5609 );
or ( n5611 , n5536 , n5610 );
and ( n5612 , n5533 , n5611 );
or ( n5613 , n5532 , n5612 );
and ( n5614 , n5529 , n5613 );
or ( n5615 , n5528 , n5614 );
and ( n5616 , n5525 , n5615 );
or ( n5617 , n5524 , n5616 );
and ( n5618 , n5521 , n5617 );
or ( n5619 , n5520 , n5618 );
and ( n5620 , n5517 , n5619 );
or ( n5621 , n5516 , n5620 );
and ( n5622 , n5513 , n5621 );
or ( n5623 , n5512 , n5622 );
and ( n5624 , n5509 , n5623 );
or ( n5625 , n5508 , n5624 );
and ( n5626 , n5505 , n5625 );
or ( n5627 , n5504 , n5626 );
and ( n5628 , n5501 , n5627 );
or ( n5629 , n5500 , n5628 );
and ( n5630 , n5497 , n5629 );
or ( n5631 , n5496 , n5630 );
and ( n5632 , n5493 , n5631 );
or ( n5633 , n5492 , n5632 );
and ( n5634 , n5489 , n5633 );
or ( n5635 , n5488 , n5634 );
and ( n5636 , n5485 , n5635 );
or ( n5637 , n5484 , n5636 );
xor ( n5638 , n5481 , n5637 );
and ( n5639 , n5422 , n5426 );
and ( n5640 , n5426 , n5462 );
and ( n5641 , n5422 , n5462 );
or ( n5642 , n5639 , n5640 , n5641 );
and ( n5643 , n5294 , n5417 );
and ( n5644 , n5417 , n5463 );
and ( n5645 , n5294 , n5463 );
or ( n5646 , n5643 , n5644 , n5645 );
xor ( n5647 , n5642 , n5646 );
and ( n5648 , n5298 , n5345 );
and ( n5649 , n5345 , n5416 );
and ( n5650 , n5298 , n5416 );
or ( n5651 , n5648 , n5649 , n5650 );
and ( n5652 , n5350 , n5376 );
and ( n5653 , n5376 , n5415 );
and ( n5654 , n5350 , n5415 );
or ( n5655 , n5652 , n5653 , n5654 );
and ( n5656 , n5311 , n5327 );
and ( n5657 , n5327 , n5343 );
and ( n5658 , n5311 , n5343 );
or ( n5659 , n5656 , n5657 , n5658 );
and ( n5660 , n5354 , n5358 );
and ( n5661 , n5358 , n5375 );
and ( n5662 , n5354 , n5375 );
or ( n5663 , n5660 , n5661 , n5662 );
xor ( n5664 , n5659 , n5663 );
and ( n5665 , n5332 , n5336 );
and ( n5666 , n5336 , n5342 );
and ( n5667 , n5332 , n5342 );
or ( n5668 , n5665 , n5666 , n5667 );
and ( n5669 , n5322 , n5323 );
and ( n5670 , n5323 , n5325 );
and ( n5671 , n5322 , n5325 );
or ( n5672 , n5669 , n5670 , n5671 );
and ( n5673 , n3182 , n940 );
and ( n5674 , n3545 , n840 );
xor ( n5675 , n5673 , n5674 );
and ( n5676 , n3801 , n771 );
xor ( n5677 , n5675 , n5676 );
xor ( n5678 , n5672 , n5677 );
and ( n5679 , n2462 , n1254 );
and ( n5680 , n2779 , n1134 );
xor ( n5681 , n5679 , n5680 );
and ( n5682 , n3024 , n1034 );
xor ( n5683 , n5681 , n5682 );
xor ( n5684 , n5678 , n5683 );
xor ( n5685 , n5668 , n5684 );
and ( n5686 , n5338 , n5339 );
and ( n5687 , n5339 , n5341 );
and ( n5688 , n5338 , n5341 );
or ( n5689 , n5686 , n5687 , n5688 );
and ( n5690 , n5364 , n5365 );
and ( n5691 , n5365 , n5367 );
and ( n5692 , n5364 , n5367 );
or ( n5693 , n5690 , n5691 , n5692 );
xor ( n5694 , n5689 , n5693 );
and ( n5695 , n1933 , n1738 );
and ( n5696 , n2120 , n1551 );
xor ( n5697 , n5695 , n5696 );
and ( n5698 , n2324 , n1424 );
xor ( n5699 , n5697 , n5698 );
xor ( n5700 , n5694 , n5699 );
xor ( n5701 , n5685 , n5700 );
xor ( n5702 , n5664 , n5701 );
xor ( n5703 , n5655 , n5702 );
and ( n5704 , n5381 , n5396 );
and ( n5705 , n5396 , n5414 );
and ( n5706 , n5381 , n5414 );
or ( n5707 , n5704 , n5705 , n5706 );
and ( n5708 , n5363 , n5368 );
and ( n5709 , n5368 , n5374 );
and ( n5710 , n5363 , n5374 );
or ( n5711 , n5708 , n5709 , n5710 );
and ( n5712 , n5385 , n5389 );
and ( n5713 , n5389 , n5395 );
and ( n5714 , n5385 , n5395 );
or ( n5715 , n5712 , n5713 , n5714 );
xor ( n5716 , n5711 , n5715 );
and ( n5717 , n5370 , n5371 );
and ( n5718 , n5371 , n5373 );
and ( n5719 , n5370 , n5373 );
or ( n5720 , n5717 , n5718 , n5719 );
and ( n5721 , n1383 , n2298 );
and ( n5722 , n1580 , n2100 );
xor ( n5723 , n5721 , n5722 );
and ( n5724 , n1694 , n1882 );
xor ( n5725 , n5723 , n5724 );
xor ( n5726 , n5720 , n5725 );
and ( n5727 , n1047 , n2981 );
and ( n5728 , n1164 , n2739 );
xor ( n5729 , n5727 , n5728 );
and ( n5730 , n1287 , n2544 );
xor ( n5731 , n5729 , n5730 );
xor ( n5732 , n5726 , n5731 );
xor ( n5733 , n5716 , n5732 );
xor ( n5734 , n5707 , n5733 );
and ( n5735 , n5401 , n5406 );
and ( n5736 , n5406 , n5413 );
and ( n5737 , n5401 , n5413 );
or ( n5738 , n5735 , n5736 , n5737 );
and ( n5739 , n5391 , n5392 );
and ( n5740 , n5392 , n5394 );
and ( n5741 , n5391 , n5394 );
or ( n5742 , n5739 , n5740 , n5741 );
and ( n5743 , n5402 , n5403 );
and ( n5744 , n5403 , n5405 );
and ( n5745 , n5402 , n5405 );
or ( n5746 , n5743 , n5744 , n5745 );
xor ( n5747 , n5742 , n5746 );
and ( n5748 , n783 , n3749 );
and ( n5749 , n856 , n3495 );
xor ( n5750 , n5748 , n5749 );
and ( n5751 , n925 , n3271 );
xor ( n5752 , n5750 , n5751 );
xor ( n5753 , n5747 , n5752 );
xor ( n5754 , n5738 , n5753 );
and ( n5755 , n5409 , n5410 );
and ( n5756 , n5410 , n5412 );
and ( n5757 , n5409 , n5412 );
or ( n5758 , n5755 , n5756 , n5757 );
and ( n5759 , n632 , n4730 );
and ( n5760 , n671 , n4403 );
xor ( n5761 , n5759 , n5760 );
and ( n5762 , n715 , n4102 );
xor ( n5763 , n5761 , n5762 );
xor ( n5764 , n5758 , n5763 );
buf ( n5765 , n441 );
and ( n5766 , n599 , n5765 );
and ( n5767 , n608 , n5408 );
xor ( n5768 , n5766 , n5767 );
and ( n5769 , n611 , n5103 );
xor ( n5770 , n5768 , n5769 );
xor ( n5771 , n5764 , n5770 );
xor ( n5772 , n5754 , n5771 );
xor ( n5773 , n5734 , n5772 );
xor ( n5774 , n5703 , n5773 );
xor ( n5775 , n5651 , n5774 );
and ( n5776 , n5302 , n5306 );
and ( n5777 , n5306 , n5344 );
and ( n5778 , n5302 , n5344 );
or ( n5779 , n5776 , n5777 , n5778 );
and ( n5780 , n5431 , n5456 );
and ( n5781 , n5456 , n5461 );
and ( n5782 , n5431 , n5461 );
or ( n5783 , n5780 , n5781 , n5782 );
xor ( n5784 , n5779 , n5783 );
and ( n5785 , n5435 , n5439 );
and ( n5786 , n5439 , n5455 );
and ( n5787 , n5435 , n5455 );
or ( n5788 , n5785 , n5786 , n5787 );
and ( n5789 , n5444 , n5448 );
and ( n5790 , n5448 , n5454 );
and ( n5791 , n5444 , n5454 );
or ( n5792 , n5789 , n5790 , n5791 );
and ( n5793 , n5315 , n5320 );
and ( n5794 , n5320 , n5326 );
and ( n5795 , n5315 , n5326 );
or ( n5796 , n5793 , n5794 , n5795 );
xor ( n5797 , n5792 , n5796 );
and ( n5798 , n5450 , n5451 );
and ( n5799 , n5451 , n5453 );
and ( n5800 , n5450 , n5453 );
or ( n5801 , n5798 , n5799 , n5800 );
and ( n5802 , n5316 , n5317 );
and ( n5803 , n5317 , n5319 );
and ( n5804 , n5316 , n5319 );
or ( n5805 , n5802 , n5803 , n5804 );
xor ( n5806 , n5801 , n5805 );
and ( n5807 , n4132 , n719 );
and ( n5808 , n4438 , n663 );
xor ( n5809 , n5807 , n5808 );
and ( n5810 , n4766 , n635 );
xor ( n5811 , n5809 , n5810 );
xor ( n5812 , n5806 , n5811 );
xor ( n5813 , n5797 , n5812 );
xor ( n5814 , n5788 , n5813 );
and ( n5815 , n5458 , n5460 );
and ( n5816 , n4959 , n606 );
and ( n5817 , n5459 , n615 );
xor ( n5818 , n5816 , n5817 );
buf ( n5819 , n441 );
and ( n5820 , n5819 , n612 );
xor ( n5821 , n5818 , n5820 );
xor ( n5822 , n5815 , n5821 );
xor ( n5823 , n5814 , n5822 );
xor ( n5824 , n5784 , n5823 );
xor ( n5825 , n5775 , n5824 );
xor ( n5826 , n5647 , n5825 );
and ( n5827 , n5285 , n5289 );
and ( n5828 , n5289 , n5464 );
and ( n5829 , n5285 , n5464 );
or ( n5830 , n5827 , n5828 , n5829 );
xor ( n5831 , n5826 , n5830 );
and ( n5832 , n5465 , n5469 );
and ( n5833 , n5470 , n5473 );
or ( n5834 , n5832 , n5833 );
xor ( n5835 , n5831 , n5834 );
buf ( n5836 , n5835 );
buf ( n5837 , n5836 );
not ( n5838 , n5837 );
buf ( n5839 , n527 );
not ( n5840 , n5839 );
nor ( n5841 , n5838 , n5840 );
xor ( n5842 , n5638 , n5841 );
xor ( n5843 , n5485 , n5635 );
nor ( n5844 , n5477 , n5840 );
and ( n5845 , n5843 , n5844 );
xor ( n5846 , n5843 , n5844 );
xor ( n5847 , n5489 , n5633 );
nor ( n5848 , n5126 , n5840 );
and ( n5849 , n5847 , n5848 );
xor ( n5850 , n5847 , n5848 );
xor ( n5851 , n5493 , n5631 );
nor ( n5852 , n4786 , n5840 );
and ( n5853 , n5851 , n5852 );
xor ( n5854 , n5851 , n5852 );
xor ( n5855 , n5497 , n5629 );
nor ( n5856 , n4458 , n5840 );
and ( n5857 , n5855 , n5856 );
xor ( n5858 , n5855 , n5856 );
xor ( n5859 , n5501 , n5627 );
nor ( n5860 , n4151 , n5840 );
and ( n5861 , n5859 , n5860 );
xor ( n5862 , n5859 , n5860 );
xor ( n5863 , n5505 , n5625 );
nor ( n5864 , n3853 , n5840 );
and ( n5865 , n5863 , n5864 );
xor ( n5866 , n5863 , n5864 );
xor ( n5867 , n5509 , n5623 );
nor ( n5868 , n3570 , n5840 );
and ( n5869 , n5867 , n5868 );
xor ( n5870 , n5867 , n5868 );
xor ( n5871 , n5513 , n5621 );
nor ( n5872 , n3300 , n5840 );
and ( n5873 , n5871 , n5872 );
xor ( n5874 , n5871 , n5872 );
xor ( n5875 , n5517 , n5619 );
nor ( n5876 , n3043 , n5840 );
and ( n5877 , n5875 , n5876 );
xor ( n5878 , n5875 , n5876 );
xor ( n5879 , n5521 , n5617 );
nor ( n5880 , n2797 , n5840 );
and ( n5881 , n5879 , n5880 );
xor ( n5882 , n5879 , n5880 );
xor ( n5883 , n5525 , n5615 );
nor ( n5884 , n2566 , n5840 );
and ( n5885 , n5883 , n5884 );
xor ( n5886 , n5883 , n5884 );
xor ( n5887 , n5529 , n5613 );
nor ( n5888 , n2343 , n5840 );
and ( n5889 , n5887 , n5888 );
xor ( n5890 , n5887 , n5888 );
xor ( n5891 , n5533 , n5611 );
nor ( n5892 , n2137 , n5840 );
and ( n5893 , n5891 , n5892 );
xor ( n5894 , n5891 , n5892 );
xor ( n5895 , n5537 , n5609 );
nor ( n5896 , n1945 , n5840 );
and ( n5897 , n5895 , n5896 );
xor ( n5898 , n5895 , n5896 );
xor ( n5899 , n5541 , n5607 );
nor ( n5900 , n1766 , n5840 );
and ( n5901 , n5899 , n5900 );
xor ( n5902 , n5899 , n5900 );
xor ( n5903 , n5545 , n5605 );
nor ( n5904 , n1598 , n5840 );
and ( n5905 , n5903 , n5904 );
xor ( n5906 , n5903 , n5904 );
xor ( n5907 , n5549 , n5603 );
nor ( n5908 , n1445 , n5840 );
and ( n5909 , n5907 , n5908 );
xor ( n5910 , n5907 , n5908 );
xor ( n5911 , n5553 , n5601 );
nor ( n5912 , n1303 , n5840 );
and ( n5913 , n5911 , n5912 );
xor ( n5914 , n5911 , n5912 );
xor ( n5915 , n5557 , n5599 );
nor ( n5916 , n1176 , n5840 );
and ( n5917 , n5915 , n5916 );
xor ( n5918 , n5915 , n5916 );
xor ( n5919 , n5561 , n5597 );
nor ( n5920 , n1062 , n5840 );
and ( n5921 , n5919 , n5920 );
xor ( n5922 , n5919 , n5920 );
xor ( n5923 , n5565 , n5595 );
nor ( n5924 , n958 , n5840 );
and ( n5925 , n5923 , n5924 );
xor ( n5926 , n5923 , n5924 );
xor ( n5927 , n5569 , n5593 );
nor ( n5928 , n868 , n5840 );
and ( n5929 , n5927 , n5928 );
xor ( n5930 , n5927 , n5928 );
xor ( n5931 , n5573 , n5591 );
nor ( n5932 , n796 , n5840 );
and ( n5933 , n5931 , n5932 );
xor ( n5934 , n5931 , n5932 );
xor ( n5935 , n5577 , n5589 );
nor ( n5936 , n733 , n5840 );
and ( n5937 , n5935 , n5936 );
xor ( n5938 , n5935 , n5936 );
xor ( n5939 , n5582 , n5587 );
nor ( n5940 , n684 , n5840 );
and ( n5941 , n5939 , n5940 );
xor ( n5942 , n5939 , n5940 );
xor ( n5943 , n5584 , n5585 );
buf ( n5944 , n5943 );
nor ( n5945 , n646 , n5840 );
and ( n5946 , n5944 , n5945 );
xor ( n5947 , n5944 , n5945 );
nor ( n5948 , n601 , n5128 );
buf ( n5949 , n5948 );
nor ( n5950 , n622 , n5840 );
and ( n5951 , n5949 , n5950 );
buf ( n5952 , n5951 );
and ( n5953 , n5947 , n5952 );
or ( n5954 , n5946 , n5953 );
and ( n5955 , n5942 , n5954 );
or ( n5956 , n5941 , n5955 );
and ( n5957 , n5938 , n5956 );
or ( n5958 , n5937 , n5957 );
and ( n5959 , n5934 , n5958 );
or ( n5960 , n5933 , n5959 );
and ( n5961 , n5930 , n5960 );
or ( n5962 , n5929 , n5961 );
and ( n5963 , n5926 , n5962 );
or ( n5964 , n5925 , n5963 );
and ( n5965 , n5922 , n5964 );
or ( n5966 , n5921 , n5965 );
and ( n5967 , n5918 , n5966 );
or ( n5968 , n5917 , n5967 );
and ( n5969 , n5914 , n5968 );
or ( n5970 , n5913 , n5969 );
and ( n5971 , n5910 , n5970 );
or ( n5972 , n5909 , n5971 );
and ( n5973 , n5906 , n5972 );
or ( n5974 , n5905 , n5973 );
and ( n5975 , n5902 , n5974 );
or ( n5976 , n5901 , n5975 );
and ( n5977 , n5898 , n5976 );
or ( n5978 , n5897 , n5977 );
and ( n5979 , n5894 , n5978 );
or ( n5980 , n5893 , n5979 );
and ( n5981 , n5890 , n5980 );
or ( n5982 , n5889 , n5981 );
and ( n5983 , n5886 , n5982 );
or ( n5984 , n5885 , n5983 );
and ( n5985 , n5882 , n5984 );
or ( n5986 , n5881 , n5985 );
and ( n5987 , n5878 , n5986 );
or ( n5988 , n5877 , n5987 );
and ( n5989 , n5874 , n5988 );
or ( n5990 , n5873 , n5989 );
and ( n5991 , n5870 , n5990 );
or ( n5992 , n5869 , n5991 );
and ( n5993 , n5866 , n5992 );
or ( n5994 , n5865 , n5993 );
and ( n5995 , n5862 , n5994 );
or ( n5996 , n5861 , n5995 );
and ( n5997 , n5858 , n5996 );
or ( n5998 , n5857 , n5997 );
and ( n5999 , n5854 , n5998 );
or ( n6000 , n5853 , n5999 );
and ( n6001 , n5850 , n6000 );
or ( n6002 , n5849 , n6001 );
and ( n6003 , n5846 , n6002 );
or ( n6004 , n5845 , n6003 );
xor ( n6005 , n5842 , n6004 );
and ( n6006 , n5779 , n5783 );
and ( n6007 , n5783 , n5823 );
and ( n6008 , n5779 , n5823 );
or ( n6009 , n6006 , n6007 , n6008 );
and ( n6010 , n5651 , n5774 );
and ( n6011 , n5774 , n5824 );
and ( n6012 , n5651 , n5824 );
or ( n6013 , n6010 , n6011 , n6012 );
xor ( n6014 , n6009 , n6013 );
and ( n6015 , n5655 , n5702 );
and ( n6016 , n5702 , n5773 );
and ( n6017 , n5655 , n5773 );
or ( n6018 , n6015 , n6016 , n6017 );
and ( n6019 , n5707 , n5733 );
and ( n6020 , n5733 , n5772 );
and ( n6021 , n5707 , n5772 );
or ( n6022 , n6019 , n6020 , n6021 );
and ( n6023 , n5668 , n5684 );
and ( n6024 , n5684 , n5700 );
and ( n6025 , n5668 , n5700 );
or ( n6026 , n6023 , n6024 , n6025 );
and ( n6027 , n5711 , n5715 );
and ( n6028 , n5715 , n5732 );
and ( n6029 , n5711 , n5732 );
or ( n6030 , n6027 , n6028 , n6029 );
xor ( n6031 , n6026 , n6030 );
and ( n6032 , n5689 , n5693 );
and ( n6033 , n5693 , n5699 );
and ( n6034 , n5689 , n5699 );
or ( n6035 , n6032 , n6033 , n6034 );
and ( n6036 , n5679 , n5680 );
and ( n6037 , n5680 , n5682 );
and ( n6038 , n5679 , n5682 );
or ( n6039 , n6036 , n6037 , n6038 );
and ( n6040 , n3182 , n1034 );
and ( n6041 , n3545 , n940 );
xor ( n6042 , n6040 , n6041 );
and ( n6043 , n3801 , n840 );
xor ( n6044 , n6042 , n6043 );
xor ( n6045 , n6039 , n6044 );
and ( n6046 , n2462 , n1424 );
and ( n6047 , n2779 , n1254 );
xor ( n6048 , n6046 , n6047 );
and ( n6049 , n3024 , n1134 );
xor ( n6050 , n6048 , n6049 );
xor ( n6051 , n6045 , n6050 );
xor ( n6052 , n6035 , n6051 );
and ( n6053 , n5695 , n5696 );
and ( n6054 , n5696 , n5698 );
and ( n6055 , n5695 , n5698 );
or ( n6056 , n6053 , n6054 , n6055 );
and ( n6057 , n5721 , n5722 );
and ( n6058 , n5722 , n5724 );
and ( n6059 , n5721 , n5724 );
or ( n6060 , n6057 , n6058 , n6059 );
xor ( n6061 , n6056 , n6060 );
buf ( n6062 , n1933 );
and ( n6063 , n2120 , n1738 );
xor ( n6064 , n6062 , n6063 );
and ( n6065 , n2324 , n1551 );
xor ( n6066 , n6064 , n6065 );
xor ( n6067 , n6061 , n6066 );
xor ( n6068 , n6052 , n6067 );
xor ( n6069 , n6031 , n6068 );
xor ( n6070 , n6022 , n6069 );
and ( n6071 , n5738 , n5753 );
and ( n6072 , n5753 , n5771 );
and ( n6073 , n5738 , n5771 );
or ( n6074 , n6071 , n6072 , n6073 );
and ( n6075 , n5720 , n5725 );
and ( n6076 , n5725 , n5731 );
and ( n6077 , n5720 , n5731 );
or ( n6078 , n6075 , n6076 , n6077 );
and ( n6079 , n5742 , n5746 );
and ( n6080 , n5746 , n5752 );
and ( n6081 , n5742 , n5752 );
or ( n6082 , n6079 , n6080 , n6081 );
xor ( n6083 , n6078 , n6082 );
and ( n6084 , n5727 , n5728 );
and ( n6085 , n5728 , n5730 );
and ( n6086 , n5727 , n5730 );
or ( n6087 , n6084 , n6085 , n6086 );
and ( n6088 , n1383 , n2544 );
and ( n6089 , n1580 , n2298 );
xor ( n6090 , n6088 , n6089 );
and ( n6091 , n1694 , n2100 );
xor ( n6092 , n6090 , n6091 );
xor ( n6093 , n6087 , n6092 );
and ( n6094 , n1047 , n3271 );
and ( n6095 , n1164 , n2981 );
xor ( n6096 , n6094 , n6095 );
and ( n6097 , n1287 , n2739 );
xor ( n6098 , n6096 , n6097 );
xor ( n6099 , n6093 , n6098 );
xor ( n6100 , n6083 , n6099 );
xor ( n6101 , n6074 , n6100 );
and ( n6102 , n5758 , n5763 );
and ( n6103 , n5763 , n5770 );
and ( n6104 , n5758 , n5770 );
or ( n6105 , n6102 , n6103 , n6104 );
and ( n6106 , n5748 , n5749 );
and ( n6107 , n5749 , n5751 );
and ( n6108 , n5748 , n5751 );
or ( n6109 , n6106 , n6107 , n6108 );
and ( n6110 , n5759 , n5760 );
and ( n6111 , n5760 , n5762 );
and ( n6112 , n5759 , n5762 );
or ( n6113 , n6110 , n6111 , n6112 );
xor ( n6114 , n6109 , n6113 );
and ( n6115 , n783 , n4102 );
and ( n6116 , n856 , n3749 );
xor ( n6117 , n6115 , n6116 );
and ( n6118 , n925 , n3495 );
xor ( n6119 , n6117 , n6118 );
xor ( n6120 , n6114 , n6119 );
xor ( n6121 , n6105 , n6120 );
and ( n6122 , n5766 , n5767 );
and ( n6123 , n5767 , n5769 );
and ( n6124 , n5766 , n5769 );
or ( n6125 , n6122 , n6123 , n6124 );
and ( n6126 , n632 , n5103 );
and ( n6127 , n671 , n4730 );
xor ( n6128 , n6126 , n6127 );
and ( n6129 , n715 , n4403 );
xor ( n6130 , n6128 , n6129 );
xor ( n6131 , n6125 , n6130 );
buf ( n6132 , n440 );
and ( n6133 , n599 , n6132 );
and ( n6134 , n608 , n5765 );
xor ( n6135 , n6133 , n6134 );
and ( n6136 , n611 , n5408 );
xor ( n6137 , n6135 , n6136 );
xor ( n6138 , n6131 , n6137 );
xor ( n6139 , n6121 , n6138 );
xor ( n6140 , n6101 , n6139 );
xor ( n6141 , n6070 , n6140 );
xor ( n6142 , n6018 , n6141 );
and ( n6143 , n5659 , n5663 );
and ( n6144 , n5663 , n5701 );
and ( n6145 , n5659 , n5701 );
or ( n6146 , n6143 , n6144 , n6145 );
and ( n6147 , n5788 , n5813 );
and ( n6148 , n5813 , n5822 );
and ( n6149 , n5788 , n5822 );
or ( n6150 , n6147 , n6148 , n6149 );
xor ( n6151 , n6146 , n6150 );
and ( n6152 , n5792 , n5796 );
and ( n6153 , n5796 , n5812 );
and ( n6154 , n5792 , n5812 );
or ( n6155 , n6152 , n6153 , n6154 );
and ( n6156 , n5801 , n5805 );
and ( n6157 , n5805 , n5811 );
and ( n6158 , n5801 , n5811 );
or ( n6159 , n6156 , n6157 , n6158 );
and ( n6160 , n5672 , n5677 );
and ( n6161 , n5677 , n5683 );
and ( n6162 , n5672 , n5683 );
or ( n6163 , n6160 , n6161 , n6162 );
xor ( n6164 , n6159 , n6163 );
and ( n6165 , n5807 , n5808 );
and ( n6166 , n5808 , n5810 );
and ( n6167 , n5807 , n5810 );
or ( n6168 , n6165 , n6166 , n6167 );
and ( n6169 , n5673 , n5674 );
and ( n6170 , n5674 , n5676 );
and ( n6171 , n5673 , n5676 );
or ( n6172 , n6169 , n6170 , n6171 );
xor ( n6173 , n6168 , n6172 );
and ( n6174 , n4132 , n771 );
and ( n6175 , n4438 , n719 );
xor ( n6176 , n6174 , n6175 );
and ( n6177 , n4766 , n663 );
xor ( n6178 , n6176 , n6177 );
xor ( n6179 , n6173 , n6178 );
xor ( n6180 , n6164 , n6179 );
xor ( n6181 , n6155 , n6180 );
and ( n6182 , n5815 , n5821 );
and ( n6183 , n5816 , n5817 );
and ( n6184 , n5817 , n5820 );
and ( n6185 , n5816 , n5820 );
or ( n6186 , n6183 , n6184 , n6185 );
buf ( n6187 , n440 );
and ( n6188 , n6187 , n612 );
xor ( n6189 , n6186 , n6188 );
and ( n6190 , n4959 , n635 );
and ( n6191 , n5459 , n606 );
xor ( n6192 , n6190 , n6191 );
and ( n6193 , n5819 , n615 );
xor ( n6194 , n6192 , n6193 );
xor ( n6195 , n6189 , n6194 );
xor ( n6196 , n6182 , n6195 );
xor ( n6197 , n6181 , n6196 );
xor ( n6198 , n6151 , n6197 );
xor ( n6199 , n6142 , n6198 );
xor ( n6200 , n6014 , n6199 );
and ( n6201 , n5642 , n5646 );
and ( n6202 , n5646 , n5825 );
and ( n6203 , n5642 , n5825 );
or ( n6204 , n6201 , n6202 , n6203 );
xor ( n6205 , n6200 , n6204 );
and ( n6206 , n5826 , n5830 );
and ( n6207 , n5831 , n5834 );
or ( n6208 , n6206 , n6207 );
xor ( n6209 , n6205 , n6208 );
buf ( n6210 , n6209 );
buf ( n6211 , n6210 );
not ( n6212 , n6211 );
buf ( n6213 , n528 );
not ( n6214 , n6213 );
nor ( n6215 , n6212 , n6214 );
xor ( n6216 , n6005 , n6215 );
xor ( n6217 , n5846 , n6002 );
nor ( n6218 , n5838 , n6214 );
and ( n6219 , n6217 , n6218 );
xor ( n6220 , n6217 , n6218 );
xor ( n6221 , n5850 , n6000 );
nor ( n6222 , n5477 , n6214 );
and ( n6223 , n6221 , n6222 );
xor ( n6224 , n6221 , n6222 );
xor ( n6225 , n5854 , n5998 );
nor ( n6226 , n5126 , n6214 );
and ( n6227 , n6225 , n6226 );
xor ( n6228 , n6225 , n6226 );
xor ( n6229 , n5858 , n5996 );
nor ( n6230 , n4786 , n6214 );
and ( n6231 , n6229 , n6230 );
xor ( n6232 , n6229 , n6230 );
xor ( n6233 , n5862 , n5994 );
nor ( n6234 , n4458 , n6214 );
and ( n6235 , n6233 , n6234 );
xor ( n6236 , n6233 , n6234 );
xor ( n6237 , n5866 , n5992 );
nor ( n6238 , n4151 , n6214 );
and ( n6239 , n6237 , n6238 );
xor ( n6240 , n6237 , n6238 );
xor ( n6241 , n5870 , n5990 );
nor ( n6242 , n3853 , n6214 );
and ( n6243 , n6241 , n6242 );
xor ( n6244 , n6241 , n6242 );
xor ( n6245 , n5874 , n5988 );
nor ( n6246 , n3570 , n6214 );
and ( n6247 , n6245 , n6246 );
xor ( n6248 , n6245 , n6246 );
xor ( n6249 , n5878 , n5986 );
nor ( n6250 , n3300 , n6214 );
and ( n6251 , n6249 , n6250 );
xor ( n6252 , n6249 , n6250 );
xor ( n6253 , n5882 , n5984 );
nor ( n6254 , n3043 , n6214 );
and ( n6255 , n6253 , n6254 );
xor ( n6256 , n6253 , n6254 );
xor ( n6257 , n5886 , n5982 );
nor ( n6258 , n2797 , n6214 );
and ( n6259 , n6257 , n6258 );
xor ( n6260 , n6257 , n6258 );
xor ( n6261 , n5890 , n5980 );
nor ( n6262 , n2566 , n6214 );
and ( n6263 , n6261 , n6262 );
xor ( n6264 , n6261 , n6262 );
xor ( n6265 , n5894 , n5978 );
nor ( n6266 , n2343 , n6214 );
and ( n6267 , n6265 , n6266 );
xor ( n6268 , n6265 , n6266 );
xor ( n6269 , n5898 , n5976 );
nor ( n6270 , n2137 , n6214 );
and ( n6271 , n6269 , n6270 );
xor ( n6272 , n6269 , n6270 );
xor ( n6273 , n5902 , n5974 );
nor ( n6274 , n1945 , n6214 );
and ( n6275 , n6273 , n6274 );
xor ( n6276 , n6273 , n6274 );
xor ( n6277 , n5906 , n5972 );
nor ( n6278 , n1766 , n6214 );
and ( n6279 , n6277 , n6278 );
xor ( n6280 , n6277 , n6278 );
xor ( n6281 , n5910 , n5970 );
nor ( n6282 , n1598 , n6214 );
and ( n6283 , n6281 , n6282 );
xor ( n6284 , n6281 , n6282 );
xor ( n6285 , n5914 , n5968 );
nor ( n6286 , n1445 , n6214 );
and ( n6287 , n6285 , n6286 );
xor ( n6288 , n6285 , n6286 );
xor ( n6289 , n5918 , n5966 );
nor ( n6290 , n1303 , n6214 );
and ( n6291 , n6289 , n6290 );
xor ( n6292 , n6289 , n6290 );
xor ( n6293 , n5922 , n5964 );
nor ( n6294 , n1176 , n6214 );
and ( n6295 , n6293 , n6294 );
xor ( n6296 , n6293 , n6294 );
xor ( n6297 , n5926 , n5962 );
nor ( n6298 , n1062 , n6214 );
and ( n6299 , n6297 , n6298 );
xor ( n6300 , n6297 , n6298 );
xor ( n6301 , n5930 , n5960 );
nor ( n6302 , n958 , n6214 );
and ( n6303 , n6301 , n6302 );
xor ( n6304 , n6301 , n6302 );
xor ( n6305 , n5934 , n5958 );
nor ( n6306 , n868 , n6214 );
and ( n6307 , n6305 , n6306 );
xor ( n6308 , n6305 , n6306 );
xor ( n6309 , n5938 , n5956 );
nor ( n6310 , n796 , n6214 );
and ( n6311 , n6309 , n6310 );
xor ( n6312 , n6309 , n6310 );
xor ( n6313 , n5942 , n5954 );
nor ( n6314 , n733 , n6214 );
and ( n6315 , n6313 , n6314 );
xor ( n6316 , n6313 , n6314 );
xor ( n6317 , n5947 , n5952 );
nor ( n6318 , n684 , n6214 );
and ( n6319 , n6317 , n6318 );
xor ( n6320 , n6317 , n6318 );
xor ( n6321 , n5949 , n5950 );
buf ( n6322 , n6321 );
nor ( n6323 , n646 , n6214 );
and ( n6324 , n6322 , n6323 );
xor ( n6325 , n6322 , n6323 );
nor ( n6326 , n601 , n5479 );
buf ( n6327 , n6326 );
nor ( n6328 , n622 , n6214 );
and ( n6329 , n6327 , n6328 );
buf ( n6330 , n6329 );
and ( n6331 , n6325 , n6330 );
or ( n6332 , n6324 , n6331 );
and ( n6333 , n6320 , n6332 );
or ( n6334 , n6319 , n6333 );
and ( n6335 , n6316 , n6334 );
or ( n6336 , n6315 , n6335 );
and ( n6337 , n6312 , n6336 );
or ( n6338 , n6311 , n6337 );
and ( n6339 , n6308 , n6338 );
or ( n6340 , n6307 , n6339 );
and ( n6341 , n6304 , n6340 );
or ( n6342 , n6303 , n6341 );
and ( n6343 , n6300 , n6342 );
or ( n6344 , n6299 , n6343 );
and ( n6345 , n6296 , n6344 );
or ( n6346 , n6295 , n6345 );
and ( n6347 , n6292 , n6346 );
or ( n6348 , n6291 , n6347 );
and ( n6349 , n6288 , n6348 );
or ( n6350 , n6287 , n6349 );
and ( n6351 , n6284 , n6350 );
or ( n6352 , n6283 , n6351 );
and ( n6353 , n6280 , n6352 );
or ( n6354 , n6279 , n6353 );
and ( n6355 , n6276 , n6354 );
or ( n6356 , n6275 , n6355 );
and ( n6357 , n6272 , n6356 );
or ( n6358 , n6271 , n6357 );
and ( n6359 , n6268 , n6358 );
or ( n6360 , n6267 , n6359 );
and ( n6361 , n6264 , n6360 );
or ( n6362 , n6263 , n6361 );
and ( n6363 , n6260 , n6362 );
or ( n6364 , n6259 , n6363 );
and ( n6365 , n6256 , n6364 );
or ( n6366 , n6255 , n6365 );
and ( n6367 , n6252 , n6366 );
or ( n6368 , n6251 , n6367 );
and ( n6369 , n6248 , n6368 );
or ( n6370 , n6247 , n6369 );
and ( n6371 , n6244 , n6370 );
or ( n6372 , n6243 , n6371 );
and ( n6373 , n6240 , n6372 );
or ( n6374 , n6239 , n6373 );
and ( n6375 , n6236 , n6374 );
or ( n6376 , n6235 , n6375 );
and ( n6377 , n6232 , n6376 );
or ( n6378 , n6231 , n6377 );
and ( n6379 , n6228 , n6378 );
or ( n6380 , n6227 , n6379 );
and ( n6381 , n6224 , n6380 );
or ( n6382 , n6223 , n6381 );
and ( n6383 , n6220 , n6382 );
or ( n6384 , n6219 , n6383 );
xor ( n6385 , n6216 , n6384 );
and ( n6386 , n6018 , n6141 );
and ( n6387 , n6141 , n6198 );
and ( n6388 , n6018 , n6198 );
or ( n6389 , n6386 , n6387 , n6388 );
and ( n6390 , n6022 , n6069 );
and ( n6391 , n6069 , n6140 );
and ( n6392 , n6022 , n6140 );
or ( n6393 , n6390 , n6391 , n6392 );
and ( n6394 , n6074 , n6100 );
and ( n6395 , n6100 , n6139 );
and ( n6396 , n6074 , n6139 );
or ( n6397 , n6394 , n6395 , n6396 );
and ( n6398 , n6035 , n6051 );
and ( n6399 , n6051 , n6067 );
and ( n6400 , n6035 , n6067 );
or ( n6401 , n6398 , n6399 , n6400 );
and ( n6402 , n6078 , n6082 );
and ( n6403 , n6082 , n6099 );
and ( n6404 , n6078 , n6099 );
or ( n6405 , n6402 , n6403 , n6404 );
xor ( n6406 , n6401 , n6405 );
and ( n6407 , n6056 , n6060 );
and ( n6408 , n6060 , n6066 );
and ( n6409 , n6056 , n6066 );
or ( n6410 , n6407 , n6408 , n6409 );
and ( n6411 , n6046 , n6047 );
and ( n6412 , n6047 , n6049 );
and ( n6413 , n6046 , n6049 );
or ( n6414 , n6411 , n6412 , n6413 );
and ( n6415 , n3182 , n1134 );
and ( n6416 , n3545 , n1034 );
xor ( n6417 , n6415 , n6416 );
and ( n6418 , n3801 , n940 );
xor ( n6419 , n6417 , n6418 );
xor ( n6420 , n6414 , n6419 );
and ( n6421 , n2462 , n1551 );
and ( n6422 , n2779 , n1424 );
xor ( n6423 , n6421 , n6422 );
and ( n6424 , n3024 , n1254 );
xor ( n6425 , n6423 , n6424 );
xor ( n6426 , n6420 , n6425 );
xor ( n6427 , n6410 , n6426 );
and ( n6428 , n6062 , n6063 );
and ( n6429 , n6063 , n6065 );
and ( n6430 , n6062 , n6065 );
or ( n6431 , n6428 , n6429 , n6430 );
and ( n6432 , n6088 , n6089 );
and ( n6433 , n6089 , n6091 );
and ( n6434 , n6088 , n6091 );
or ( n6435 , n6432 , n6433 , n6434 );
xor ( n6436 , n6431 , n6435 );
and ( n6437 , n2324 , n1738 );
buf ( n6438 , n6437 );
xor ( n6439 , n6436 , n6438 );
xor ( n6440 , n6427 , n6439 );
xor ( n6441 , n6406 , n6440 );
xor ( n6442 , n6397 , n6441 );
and ( n6443 , n6105 , n6120 );
and ( n6444 , n6120 , n6138 );
and ( n6445 , n6105 , n6138 );
or ( n6446 , n6443 , n6444 , n6445 );
and ( n6447 , n6087 , n6092 );
and ( n6448 , n6092 , n6098 );
and ( n6449 , n6087 , n6098 );
or ( n6450 , n6447 , n6448 , n6449 );
and ( n6451 , n6109 , n6113 );
and ( n6452 , n6113 , n6119 );
and ( n6453 , n6109 , n6119 );
or ( n6454 , n6451 , n6452 , n6453 );
xor ( n6455 , n6450 , n6454 );
and ( n6456 , n6094 , n6095 );
and ( n6457 , n6095 , n6097 );
and ( n6458 , n6094 , n6097 );
or ( n6459 , n6456 , n6457 , n6458 );
and ( n6460 , n1383 , n2739 );
and ( n6461 , n1580 , n2544 );
xor ( n6462 , n6460 , n6461 );
and ( n6463 , n1694 , n2298 );
xor ( n6464 , n6462 , n6463 );
xor ( n6465 , n6459 , n6464 );
and ( n6466 , n1047 , n3495 );
and ( n6467 , n1164 , n3271 );
xor ( n6468 , n6466 , n6467 );
and ( n6469 , n1287 , n2981 );
xor ( n6470 , n6468 , n6469 );
xor ( n6471 , n6465 , n6470 );
xor ( n6472 , n6455 , n6471 );
xor ( n6473 , n6446 , n6472 );
and ( n6474 , n6125 , n6130 );
and ( n6475 , n6130 , n6137 );
and ( n6476 , n6125 , n6137 );
or ( n6477 , n6474 , n6475 , n6476 );
and ( n6478 , n6115 , n6116 );
and ( n6479 , n6116 , n6118 );
and ( n6480 , n6115 , n6118 );
or ( n6481 , n6478 , n6479 , n6480 );
and ( n6482 , n6126 , n6127 );
and ( n6483 , n6127 , n6129 );
and ( n6484 , n6126 , n6129 );
or ( n6485 , n6482 , n6483 , n6484 );
xor ( n6486 , n6481 , n6485 );
and ( n6487 , n783 , n4403 );
and ( n6488 , n856 , n4102 );
xor ( n6489 , n6487 , n6488 );
and ( n6490 , n925 , n3749 );
xor ( n6491 , n6489 , n6490 );
xor ( n6492 , n6486 , n6491 );
xor ( n6493 , n6477 , n6492 );
and ( n6494 , n6133 , n6134 );
and ( n6495 , n6134 , n6136 );
and ( n6496 , n6133 , n6136 );
or ( n6497 , n6494 , n6495 , n6496 );
and ( n6498 , n632 , n5408 );
and ( n6499 , n671 , n5103 );
xor ( n6500 , n6498 , n6499 );
and ( n6501 , n715 , n4730 );
xor ( n6502 , n6500 , n6501 );
xor ( n6503 , n6497 , n6502 );
buf ( n6504 , n439 );
and ( n6505 , n599 , n6504 );
and ( n6506 , n608 , n6132 );
xor ( n6507 , n6505 , n6506 );
and ( n6508 , n611 , n5765 );
xor ( n6509 , n6507 , n6508 );
xor ( n6510 , n6503 , n6509 );
xor ( n6511 , n6493 , n6510 );
xor ( n6512 , n6473 , n6511 );
xor ( n6513 , n6442 , n6512 );
xor ( n6514 , n6393 , n6513 );
and ( n6515 , n6026 , n6030 );
and ( n6516 , n6030 , n6068 );
and ( n6517 , n6026 , n6068 );
or ( n6518 , n6515 , n6516 , n6517 );
and ( n6519 , n6155 , n6180 );
and ( n6520 , n6180 , n6196 );
and ( n6521 , n6155 , n6196 );
or ( n6522 , n6519 , n6520 , n6521 );
xor ( n6523 , n6518 , n6522 );
and ( n6524 , n6159 , n6163 );
and ( n6525 , n6163 , n6179 );
and ( n6526 , n6159 , n6179 );
or ( n6527 , n6524 , n6525 , n6526 );
and ( n6528 , n6168 , n6172 );
and ( n6529 , n6172 , n6178 );
and ( n6530 , n6168 , n6178 );
or ( n6531 , n6528 , n6529 , n6530 );
and ( n6532 , n6039 , n6044 );
and ( n6533 , n6044 , n6050 );
and ( n6534 , n6039 , n6050 );
or ( n6535 , n6532 , n6533 , n6534 );
xor ( n6536 , n6531 , n6535 );
and ( n6537 , n6174 , n6175 );
and ( n6538 , n6175 , n6177 );
and ( n6539 , n6174 , n6177 );
or ( n6540 , n6537 , n6538 , n6539 );
and ( n6541 , n6040 , n6041 );
and ( n6542 , n6041 , n6043 );
and ( n6543 , n6040 , n6043 );
or ( n6544 , n6541 , n6542 , n6543 );
xor ( n6545 , n6540 , n6544 );
and ( n6546 , n4132 , n840 );
and ( n6547 , n4438 , n771 );
xor ( n6548 , n6546 , n6547 );
and ( n6549 , n4766 , n719 );
xor ( n6550 , n6548 , n6549 );
xor ( n6551 , n6545 , n6550 );
xor ( n6552 , n6536 , n6551 );
xor ( n6553 , n6527 , n6552 );
and ( n6554 , n6186 , n6188 );
and ( n6555 , n6188 , n6194 );
and ( n6556 , n6186 , n6194 );
or ( n6557 , n6554 , n6555 , n6556 );
and ( n6558 , n6190 , n6191 );
and ( n6559 , n6191 , n6193 );
and ( n6560 , n6190 , n6193 );
or ( n6561 , n6558 , n6559 , n6560 );
and ( n6562 , n4959 , n663 );
and ( n6563 , n5459 , n635 );
xor ( n6564 , n6562 , n6563 );
and ( n6565 , n5819 , n606 );
xor ( n6566 , n6564 , n6565 );
xor ( n6567 , n6561 , n6566 );
and ( n6568 , n6187 , n615 );
buf ( n6569 , n439 );
and ( n6570 , n6569 , n612 );
xor ( n6571 , n6568 , n6570 );
xor ( n6572 , n6567 , n6571 );
xor ( n6573 , n6557 , n6572 );
xor ( n6574 , n6553 , n6573 );
xor ( n6575 , n6523 , n6574 );
xor ( n6576 , n6514 , n6575 );
xor ( n6577 , n6389 , n6576 );
and ( n6578 , n6182 , n6195 );
and ( n6579 , n6146 , n6150 );
and ( n6580 , n6150 , n6197 );
and ( n6581 , n6146 , n6197 );
or ( n6582 , n6579 , n6580 , n6581 );
xor ( n6583 , n6578 , n6582 );
xor ( n6584 , n6577 , n6583 );
and ( n6585 , n6009 , n6013 );
and ( n6586 , n6013 , n6199 );
and ( n6587 , n6009 , n6199 );
or ( n6588 , n6585 , n6586 , n6587 );
xor ( n6589 , n6584 , n6588 );
and ( n6590 , n6200 , n6204 );
and ( n6591 , n6205 , n6208 );
or ( n6592 , n6590 , n6591 );
xor ( n6593 , n6589 , n6592 );
buf ( n6594 , n6593 );
buf ( n6595 , n6594 );
not ( n6596 , n6595 );
buf ( n6597 , n529 );
not ( n6598 , n6597 );
nor ( n6599 , n6596 , n6598 );
xor ( n6600 , n6385 , n6599 );
xor ( n6601 , n6220 , n6382 );
nor ( n6602 , n6212 , n6598 );
and ( n6603 , n6601 , n6602 );
xor ( n6604 , n6601 , n6602 );
xor ( n6605 , n6224 , n6380 );
nor ( n6606 , n5838 , n6598 );
and ( n6607 , n6605 , n6606 );
xor ( n6608 , n6605 , n6606 );
xor ( n6609 , n6228 , n6378 );
nor ( n6610 , n5477 , n6598 );
and ( n6611 , n6609 , n6610 );
xor ( n6612 , n6609 , n6610 );
xor ( n6613 , n6232 , n6376 );
nor ( n6614 , n5126 , n6598 );
and ( n6615 , n6613 , n6614 );
xor ( n6616 , n6613 , n6614 );
xor ( n6617 , n6236 , n6374 );
nor ( n6618 , n4786 , n6598 );
and ( n6619 , n6617 , n6618 );
xor ( n6620 , n6617 , n6618 );
xor ( n6621 , n6240 , n6372 );
nor ( n6622 , n4458 , n6598 );
and ( n6623 , n6621 , n6622 );
xor ( n6624 , n6621 , n6622 );
xor ( n6625 , n6244 , n6370 );
nor ( n6626 , n4151 , n6598 );
and ( n6627 , n6625 , n6626 );
xor ( n6628 , n6625 , n6626 );
xor ( n6629 , n6248 , n6368 );
nor ( n6630 , n3853 , n6598 );
and ( n6631 , n6629 , n6630 );
xor ( n6632 , n6629 , n6630 );
xor ( n6633 , n6252 , n6366 );
nor ( n6634 , n3570 , n6598 );
and ( n6635 , n6633 , n6634 );
xor ( n6636 , n6633 , n6634 );
xor ( n6637 , n6256 , n6364 );
nor ( n6638 , n3300 , n6598 );
and ( n6639 , n6637 , n6638 );
xor ( n6640 , n6637 , n6638 );
xor ( n6641 , n6260 , n6362 );
nor ( n6642 , n3043 , n6598 );
and ( n6643 , n6641 , n6642 );
xor ( n6644 , n6641 , n6642 );
xor ( n6645 , n6264 , n6360 );
nor ( n6646 , n2797 , n6598 );
and ( n6647 , n6645 , n6646 );
xor ( n6648 , n6645 , n6646 );
xor ( n6649 , n6268 , n6358 );
nor ( n6650 , n2566 , n6598 );
and ( n6651 , n6649 , n6650 );
xor ( n6652 , n6649 , n6650 );
xor ( n6653 , n6272 , n6356 );
nor ( n6654 , n2343 , n6598 );
and ( n6655 , n6653 , n6654 );
xor ( n6656 , n6653 , n6654 );
xor ( n6657 , n6276 , n6354 );
nor ( n6658 , n2137 , n6598 );
and ( n6659 , n6657 , n6658 );
xor ( n6660 , n6657 , n6658 );
xor ( n6661 , n6280 , n6352 );
nor ( n6662 , n1945 , n6598 );
and ( n6663 , n6661 , n6662 );
xor ( n6664 , n6661 , n6662 );
xor ( n6665 , n6284 , n6350 );
nor ( n6666 , n1766 , n6598 );
and ( n6667 , n6665 , n6666 );
xor ( n6668 , n6665 , n6666 );
xor ( n6669 , n6288 , n6348 );
nor ( n6670 , n1598 , n6598 );
and ( n6671 , n6669 , n6670 );
xor ( n6672 , n6669 , n6670 );
xor ( n6673 , n6292 , n6346 );
nor ( n6674 , n1445 , n6598 );
and ( n6675 , n6673 , n6674 );
xor ( n6676 , n6673 , n6674 );
xor ( n6677 , n6296 , n6344 );
nor ( n6678 , n1303 , n6598 );
and ( n6679 , n6677 , n6678 );
xor ( n6680 , n6677 , n6678 );
xor ( n6681 , n6300 , n6342 );
nor ( n6682 , n1176 , n6598 );
and ( n6683 , n6681 , n6682 );
xor ( n6684 , n6681 , n6682 );
xor ( n6685 , n6304 , n6340 );
nor ( n6686 , n1062 , n6598 );
and ( n6687 , n6685 , n6686 );
xor ( n6688 , n6685 , n6686 );
xor ( n6689 , n6308 , n6338 );
nor ( n6690 , n958 , n6598 );
and ( n6691 , n6689 , n6690 );
xor ( n6692 , n6689 , n6690 );
xor ( n6693 , n6312 , n6336 );
nor ( n6694 , n868 , n6598 );
and ( n6695 , n6693 , n6694 );
xor ( n6696 , n6693 , n6694 );
xor ( n6697 , n6316 , n6334 );
nor ( n6698 , n796 , n6598 );
and ( n6699 , n6697 , n6698 );
xor ( n6700 , n6697 , n6698 );
xor ( n6701 , n6320 , n6332 );
nor ( n6702 , n733 , n6598 );
and ( n6703 , n6701 , n6702 );
xor ( n6704 , n6701 , n6702 );
xor ( n6705 , n6325 , n6330 );
nor ( n6706 , n684 , n6598 );
and ( n6707 , n6705 , n6706 );
xor ( n6708 , n6705 , n6706 );
xor ( n6709 , n6327 , n6328 );
buf ( n6710 , n6709 );
nor ( n6711 , n646 , n6598 );
and ( n6712 , n6710 , n6711 );
xor ( n6713 , n6710 , n6711 );
nor ( n6714 , n601 , n5840 );
buf ( n6715 , n6714 );
nor ( n6716 , n622 , n6598 );
and ( n6717 , n6715 , n6716 );
buf ( n6718 , n6717 );
and ( n6719 , n6713 , n6718 );
or ( n6720 , n6712 , n6719 );
and ( n6721 , n6708 , n6720 );
or ( n6722 , n6707 , n6721 );
and ( n6723 , n6704 , n6722 );
or ( n6724 , n6703 , n6723 );
and ( n6725 , n6700 , n6724 );
or ( n6726 , n6699 , n6725 );
and ( n6727 , n6696 , n6726 );
or ( n6728 , n6695 , n6727 );
and ( n6729 , n6692 , n6728 );
or ( n6730 , n6691 , n6729 );
and ( n6731 , n6688 , n6730 );
or ( n6732 , n6687 , n6731 );
and ( n6733 , n6684 , n6732 );
or ( n6734 , n6683 , n6733 );
and ( n6735 , n6680 , n6734 );
or ( n6736 , n6679 , n6735 );
and ( n6737 , n6676 , n6736 );
or ( n6738 , n6675 , n6737 );
and ( n6739 , n6672 , n6738 );
or ( n6740 , n6671 , n6739 );
and ( n6741 , n6668 , n6740 );
or ( n6742 , n6667 , n6741 );
and ( n6743 , n6664 , n6742 );
or ( n6744 , n6663 , n6743 );
and ( n6745 , n6660 , n6744 );
or ( n6746 , n6659 , n6745 );
and ( n6747 , n6656 , n6746 );
or ( n6748 , n6655 , n6747 );
and ( n6749 , n6652 , n6748 );
or ( n6750 , n6651 , n6749 );
and ( n6751 , n6648 , n6750 );
or ( n6752 , n6647 , n6751 );
and ( n6753 , n6644 , n6752 );
or ( n6754 , n6643 , n6753 );
and ( n6755 , n6640 , n6754 );
or ( n6756 , n6639 , n6755 );
and ( n6757 , n6636 , n6756 );
or ( n6758 , n6635 , n6757 );
and ( n6759 , n6632 , n6758 );
or ( n6760 , n6631 , n6759 );
and ( n6761 , n6628 , n6760 );
or ( n6762 , n6627 , n6761 );
and ( n6763 , n6624 , n6762 );
or ( n6764 , n6623 , n6763 );
and ( n6765 , n6620 , n6764 );
or ( n6766 , n6619 , n6765 );
and ( n6767 , n6616 , n6766 );
or ( n6768 , n6615 , n6767 );
and ( n6769 , n6612 , n6768 );
or ( n6770 , n6611 , n6769 );
and ( n6771 , n6608 , n6770 );
or ( n6772 , n6607 , n6771 );
and ( n6773 , n6604 , n6772 );
or ( n6774 , n6603 , n6773 );
xor ( n6775 , n6600 , n6774 );
and ( n6776 , n6578 , n6582 );
and ( n6777 , n6389 , n6576 );
and ( n6778 , n6576 , n6583 );
and ( n6779 , n6389 , n6583 );
or ( n6780 , n6777 , n6778 , n6779 );
xor ( n6781 , n6776 , n6780 );
and ( n6782 , n6393 , n6513 );
and ( n6783 , n6513 , n6575 );
and ( n6784 , n6393 , n6575 );
or ( n6785 , n6782 , n6783 , n6784 );
and ( n6786 , n6397 , n6441 );
and ( n6787 , n6441 , n6512 );
and ( n6788 , n6397 , n6512 );
or ( n6789 , n6786 , n6787 , n6788 );
and ( n6790 , n6401 , n6405 );
and ( n6791 , n6405 , n6440 );
and ( n6792 , n6401 , n6440 );
or ( n6793 , n6790 , n6791 , n6792 );
and ( n6794 , n6527 , n6552 );
and ( n6795 , n6552 , n6573 );
and ( n6796 , n6527 , n6573 );
or ( n6797 , n6794 , n6795 , n6796 );
xor ( n6798 , n6793 , n6797 );
and ( n6799 , n6531 , n6535 );
and ( n6800 , n6535 , n6551 );
and ( n6801 , n6531 , n6551 );
or ( n6802 , n6799 , n6800 , n6801 );
and ( n6803 , n6568 , n6570 );
and ( n6804 , n6561 , n6566 );
and ( n6805 , n6566 , n6571 );
and ( n6806 , n6561 , n6571 );
or ( n6807 , n6804 , n6805 , n6806 );
xor ( n6808 , n6803 , n6807 );
and ( n6809 , n6562 , n6563 );
and ( n6810 , n6563 , n6565 );
and ( n6811 , n6562 , n6565 );
or ( n6812 , n6809 , n6810 , n6811 );
and ( n6813 , n6187 , n606 );
and ( n6814 , n6569 , n615 );
xor ( n6815 , n6813 , n6814 );
buf ( n6816 , n438 );
and ( n6817 , n6816 , n612 );
xor ( n6818 , n6815 , n6817 );
xor ( n6819 , n6812 , n6818 );
and ( n6820 , n4959 , n719 );
and ( n6821 , n5459 , n663 );
xor ( n6822 , n6820 , n6821 );
and ( n6823 , n5819 , n635 );
xor ( n6824 , n6822 , n6823 );
xor ( n6825 , n6819 , n6824 );
xor ( n6826 , n6808 , n6825 );
xor ( n6827 , n6802 , n6826 );
and ( n6828 , n6540 , n6544 );
and ( n6829 , n6544 , n6550 );
and ( n6830 , n6540 , n6550 );
or ( n6831 , n6828 , n6829 , n6830 );
and ( n6832 , n6414 , n6419 );
and ( n6833 , n6419 , n6425 );
and ( n6834 , n6414 , n6425 );
or ( n6835 , n6832 , n6833 , n6834 );
xor ( n6836 , n6831 , n6835 );
and ( n6837 , n6546 , n6547 );
and ( n6838 , n6547 , n6549 );
and ( n6839 , n6546 , n6549 );
or ( n6840 , n6837 , n6838 , n6839 );
and ( n6841 , n6415 , n6416 );
and ( n6842 , n6416 , n6418 );
and ( n6843 , n6415 , n6418 );
or ( n6844 , n6841 , n6842 , n6843 );
xor ( n6845 , n6840 , n6844 );
and ( n6846 , n4132 , n940 );
and ( n6847 , n4438 , n840 );
xor ( n6848 , n6846 , n6847 );
and ( n6849 , n4766 , n771 );
xor ( n6850 , n6848 , n6849 );
xor ( n6851 , n6845 , n6850 );
xor ( n6852 , n6836 , n6851 );
xor ( n6853 , n6827 , n6852 );
xor ( n6854 , n6798 , n6853 );
xor ( n6855 , n6789 , n6854 );
and ( n6856 , n6446 , n6472 );
and ( n6857 , n6472 , n6511 );
and ( n6858 , n6446 , n6511 );
or ( n6859 , n6856 , n6857 , n6858 );
and ( n6860 , n6410 , n6426 );
and ( n6861 , n6426 , n6439 );
and ( n6862 , n6410 , n6439 );
or ( n6863 , n6860 , n6861 , n6862 );
and ( n6864 , n6450 , n6454 );
and ( n6865 , n6454 , n6471 );
and ( n6866 , n6450 , n6471 );
or ( n6867 , n6864 , n6865 , n6866 );
xor ( n6868 , n6863 , n6867 );
and ( n6869 , n6431 , n6435 );
and ( n6870 , n6435 , n6438 );
and ( n6871 , n6431 , n6438 );
or ( n6872 , n6869 , n6870 , n6871 );
and ( n6873 , n6421 , n6422 );
and ( n6874 , n6422 , n6424 );
and ( n6875 , n6421 , n6424 );
or ( n6876 , n6873 , n6874 , n6875 );
and ( n6877 , n3182 , n1254 );
and ( n6878 , n3545 , n1134 );
xor ( n6879 , n6877 , n6878 );
and ( n6880 , n3801 , n1034 );
xor ( n6881 , n6879 , n6880 );
xor ( n6882 , n6876 , n6881 );
and ( n6883 , n2462 , n1738 );
and ( n6884 , n2779 , n1551 );
xor ( n6885 , n6883 , n6884 );
and ( n6886 , n3024 , n1424 );
xor ( n6887 , n6885 , n6886 );
xor ( n6888 , n6882 , n6887 );
xor ( n6889 , n6872 , n6888 );
and ( n6890 , n1933 , n2100 );
and ( n6891 , n2120 , n1882 );
and ( n6892 , n6890 , n6891 );
and ( n6893 , n6891 , n6437 );
and ( n6894 , n6890 , n6437 );
or ( n6895 , n6892 , n6893 , n6894 );
and ( n6896 , n6460 , n6461 );
and ( n6897 , n6461 , n6463 );
and ( n6898 , n6460 , n6463 );
or ( n6899 , n6896 , n6897 , n6898 );
xor ( n6900 , n6895 , n6899 );
and ( n6901 , n1933 , n2298 );
buf ( n6902 , n2120 );
xor ( n6903 , n6901 , n6902 );
and ( n6904 , n2324 , n1882 );
xor ( n6905 , n6903 , n6904 );
xor ( n6906 , n6900 , n6905 );
xor ( n6907 , n6889 , n6906 );
xor ( n6908 , n6868 , n6907 );
xor ( n6909 , n6859 , n6908 );
and ( n6910 , n6477 , n6492 );
and ( n6911 , n6492 , n6510 );
and ( n6912 , n6477 , n6510 );
or ( n6913 , n6910 , n6911 , n6912 );
and ( n6914 , n6459 , n6464 );
and ( n6915 , n6464 , n6470 );
and ( n6916 , n6459 , n6470 );
or ( n6917 , n6914 , n6915 , n6916 );
and ( n6918 , n6481 , n6485 );
and ( n6919 , n6485 , n6491 );
and ( n6920 , n6481 , n6491 );
or ( n6921 , n6918 , n6919 , n6920 );
xor ( n6922 , n6917 , n6921 );
and ( n6923 , n6466 , n6467 );
and ( n6924 , n6467 , n6469 );
and ( n6925 , n6466 , n6469 );
or ( n6926 , n6923 , n6924 , n6925 );
and ( n6927 , n1383 , n2981 );
and ( n6928 , n1580 , n2739 );
xor ( n6929 , n6927 , n6928 );
and ( n6930 , n1694 , n2544 );
xor ( n6931 , n6929 , n6930 );
xor ( n6932 , n6926 , n6931 );
and ( n6933 , n1047 , n3749 );
and ( n6934 , n1164 , n3495 );
xor ( n6935 , n6933 , n6934 );
and ( n6936 , n1287 , n3271 );
xor ( n6937 , n6935 , n6936 );
xor ( n6938 , n6932 , n6937 );
xor ( n6939 , n6922 , n6938 );
xor ( n6940 , n6913 , n6939 );
and ( n6941 , n6497 , n6502 );
and ( n6942 , n6502 , n6509 );
and ( n6943 , n6497 , n6509 );
or ( n6944 , n6941 , n6942 , n6943 );
and ( n6945 , n6487 , n6488 );
and ( n6946 , n6488 , n6490 );
and ( n6947 , n6487 , n6490 );
or ( n6948 , n6945 , n6946 , n6947 );
and ( n6949 , n6498 , n6499 );
and ( n6950 , n6499 , n6501 );
and ( n6951 , n6498 , n6501 );
or ( n6952 , n6949 , n6950 , n6951 );
xor ( n6953 , n6948 , n6952 );
and ( n6954 , n783 , n4730 );
and ( n6955 , n856 , n4403 );
xor ( n6956 , n6954 , n6955 );
and ( n6957 , n925 , n4102 );
xor ( n6958 , n6956 , n6957 );
xor ( n6959 , n6953 , n6958 );
xor ( n6960 , n6944 , n6959 );
and ( n6961 , n6505 , n6506 );
and ( n6962 , n6506 , n6508 );
and ( n6963 , n6505 , n6508 );
or ( n6964 , n6961 , n6962 , n6963 );
and ( n6965 , n632 , n5765 );
and ( n6966 , n671 , n5408 );
xor ( n6967 , n6965 , n6966 );
and ( n6968 , n715 , n5103 );
xor ( n6969 , n6967 , n6968 );
xor ( n6970 , n6964 , n6969 );
buf ( n6971 , n438 );
and ( n6972 , n599 , n6971 );
and ( n6973 , n608 , n6504 );
xor ( n6974 , n6972 , n6973 );
and ( n6975 , n611 , n6132 );
xor ( n6976 , n6974 , n6975 );
xor ( n6977 , n6970 , n6976 );
xor ( n6978 , n6960 , n6977 );
xor ( n6979 , n6940 , n6978 );
xor ( n6980 , n6909 , n6979 );
xor ( n6981 , n6855 , n6980 );
xor ( n6982 , n6785 , n6981 );
and ( n6983 , n6557 , n6572 );
and ( n6984 , n6518 , n6522 );
and ( n6985 , n6522 , n6574 );
and ( n6986 , n6518 , n6574 );
or ( n6987 , n6984 , n6985 , n6986 );
xor ( n6988 , n6983 , n6987 );
xor ( n6989 , n6982 , n6988 );
xor ( n6990 , n6781 , n6989 );
and ( n6991 , n6584 , n6588 );
and ( n6992 , n6589 , n6592 );
or ( n6993 , n6991 , n6992 );
xor ( n6994 , n6990 , n6993 );
buf ( n6995 , n6994 );
buf ( n6996 , n6995 );
not ( n6997 , n6996 );
buf ( n6998 , n530 );
not ( n6999 , n6998 );
nor ( n7000 , n6997 , n6999 );
xor ( n7001 , n6775 , n7000 );
xor ( n7002 , n6604 , n6772 );
nor ( n7003 , n6596 , n6999 );
and ( n7004 , n7002 , n7003 );
xor ( n7005 , n7002 , n7003 );
xor ( n7006 , n6608 , n6770 );
nor ( n7007 , n6212 , n6999 );
and ( n7008 , n7006 , n7007 );
xor ( n7009 , n7006 , n7007 );
xor ( n7010 , n6612 , n6768 );
nor ( n7011 , n5838 , n6999 );
and ( n7012 , n7010 , n7011 );
xor ( n7013 , n7010 , n7011 );
xor ( n7014 , n6616 , n6766 );
nor ( n7015 , n5477 , n6999 );
and ( n7016 , n7014 , n7015 );
xor ( n7017 , n7014 , n7015 );
xor ( n7018 , n6620 , n6764 );
nor ( n7019 , n5126 , n6999 );
and ( n7020 , n7018 , n7019 );
xor ( n7021 , n7018 , n7019 );
xor ( n7022 , n6624 , n6762 );
nor ( n7023 , n4786 , n6999 );
and ( n7024 , n7022 , n7023 );
xor ( n7025 , n7022 , n7023 );
xor ( n7026 , n6628 , n6760 );
nor ( n7027 , n4458 , n6999 );
and ( n7028 , n7026 , n7027 );
xor ( n7029 , n7026 , n7027 );
xor ( n7030 , n6632 , n6758 );
nor ( n7031 , n4151 , n6999 );
and ( n7032 , n7030 , n7031 );
xor ( n7033 , n7030 , n7031 );
xor ( n7034 , n6636 , n6756 );
nor ( n7035 , n3853 , n6999 );
and ( n7036 , n7034 , n7035 );
xor ( n7037 , n7034 , n7035 );
xor ( n7038 , n6640 , n6754 );
nor ( n7039 , n3570 , n6999 );
and ( n7040 , n7038 , n7039 );
xor ( n7041 , n7038 , n7039 );
xor ( n7042 , n6644 , n6752 );
nor ( n7043 , n3300 , n6999 );
and ( n7044 , n7042 , n7043 );
xor ( n7045 , n7042 , n7043 );
xor ( n7046 , n6648 , n6750 );
nor ( n7047 , n3043 , n6999 );
and ( n7048 , n7046 , n7047 );
xor ( n7049 , n7046 , n7047 );
xor ( n7050 , n6652 , n6748 );
nor ( n7051 , n2797 , n6999 );
and ( n7052 , n7050 , n7051 );
xor ( n7053 , n7050 , n7051 );
xor ( n7054 , n6656 , n6746 );
nor ( n7055 , n2566 , n6999 );
and ( n7056 , n7054 , n7055 );
xor ( n7057 , n7054 , n7055 );
xor ( n7058 , n6660 , n6744 );
nor ( n7059 , n2343 , n6999 );
and ( n7060 , n7058 , n7059 );
xor ( n7061 , n7058 , n7059 );
xor ( n7062 , n6664 , n6742 );
nor ( n7063 , n2137 , n6999 );
and ( n7064 , n7062 , n7063 );
xor ( n7065 , n7062 , n7063 );
xor ( n7066 , n6668 , n6740 );
nor ( n7067 , n1945 , n6999 );
and ( n7068 , n7066 , n7067 );
xor ( n7069 , n7066 , n7067 );
xor ( n7070 , n6672 , n6738 );
nor ( n7071 , n1766 , n6999 );
and ( n7072 , n7070 , n7071 );
xor ( n7073 , n7070 , n7071 );
xor ( n7074 , n6676 , n6736 );
nor ( n7075 , n1598 , n6999 );
and ( n7076 , n7074 , n7075 );
xor ( n7077 , n7074 , n7075 );
xor ( n7078 , n6680 , n6734 );
nor ( n7079 , n1445 , n6999 );
and ( n7080 , n7078 , n7079 );
xor ( n7081 , n7078 , n7079 );
xor ( n7082 , n6684 , n6732 );
nor ( n7083 , n1303 , n6999 );
and ( n7084 , n7082 , n7083 );
xor ( n7085 , n7082 , n7083 );
xor ( n7086 , n6688 , n6730 );
nor ( n7087 , n1176 , n6999 );
and ( n7088 , n7086 , n7087 );
xor ( n7089 , n7086 , n7087 );
xor ( n7090 , n6692 , n6728 );
nor ( n7091 , n1062 , n6999 );
and ( n7092 , n7090 , n7091 );
xor ( n7093 , n7090 , n7091 );
xor ( n7094 , n6696 , n6726 );
nor ( n7095 , n958 , n6999 );
and ( n7096 , n7094 , n7095 );
xor ( n7097 , n7094 , n7095 );
xor ( n7098 , n6700 , n6724 );
nor ( n7099 , n868 , n6999 );
and ( n7100 , n7098 , n7099 );
xor ( n7101 , n7098 , n7099 );
xor ( n7102 , n6704 , n6722 );
nor ( n7103 , n796 , n6999 );
and ( n7104 , n7102 , n7103 );
xor ( n7105 , n7102 , n7103 );
xor ( n7106 , n6708 , n6720 );
nor ( n7107 , n733 , n6999 );
and ( n7108 , n7106 , n7107 );
xor ( n7109 , n7106 , n7107 );
xor ( n7110 , n6713 , n6718 );
nor ( n7111 , n684 , n6999 );
and ( n7112 , n7110 , n7111 );
xor ( n7113 , n7110 , n7111 );
xor ( n7114 , n6715 , n6716 );
buf ( n7115 , n7114 );
nor ( n7116 , n646 , n6999 );
and ( n7117 , n7115 , n7116 );
xor ( n7118 , n7115 , n7116 );
nor ( n7119 , n601 , n6214 );
buf ( n7120 , n7119 );
nor ( n7121 , n622 , n6999 );
and ( n7122 , n7120 , n7121 );
buf ( n7123 , n7122 );
and ( n7124 , n7118 , n7123 );
or ( n7125 , n7117 , n7124 );
and ( n7126 , n7113 , n7125 );
or ( n7127 , n7112 , n7126 );
and ( n7128 , n7109 , n7127 );
or ( n7129 , n7108 , n7128 );
and ( n7130 , n7105 , n7129 );
or ( n7131 , n7104 , n7130 );
and ( n7132 , n7101 , n7131 );
or ( n7133 , n7100 , n7132 );
and ( n7134 , n7097 , n7133 );
or ( n7135 , n7096 , n7134 );
and ( n7136 , n7093 , n7135 );
or ( n7137 , n7092 , n7136 );
and ( n7138 , n7089 , n7137 );
or ( n7139 , n7088 , n7138 );
and ( n7140 , n7085 , n7139 );
or ( n7141 , n7084 , n7140 );
and ( n7142 , n7081 , n7141 );
or ( n7143 , n7080 , n7142 );
and ( n7144 , n7077 , n7143 );
or ( n7145 , n7076 , n7144 );
and ( n7146 , n7073 , n7145 );
or ( n7147 , n7072 , n7146 );
and ( n7148 , n7069 , n7147 );
or ( n7149 , n7068 , n7148 );
and ( n7150 , n7065 , n7149 );
or ( n7151 , n7064 , n7150 );
and ( n7152 , n7061 , n7151 );
or ( n7153 , n7060 , n7152 );
and ( n7154 , n7057 , n7153 );
or ( n7155 , n7056 , n7154 );
and ( n7156 , n7053 , n7155 );
or ( n7157 , n7052 , n7156 );
and ( n7158 , n7049 , n7157 );
or ( n7159 , n7048 , n7158 );
and ( n7160 , n7045 , n7159 );
or ( n7161 , n7044 , n7160 );
and ( n7162 , n7041 , n7161 );
or ( n7163 , n7040 , n7162 );
and ( n7164 , n7037 , n7163 );
or ( n7165 , n7036 , n7164 );
and ( n7166 , n7033 , n7165 );
or ( n7167 , n7032 , n7166 );
and ( n7168 , n7029 , n7167 );
or ( n7169 , n7028 , n7168 );
and ( n7170 , n7025 , n7169 );
or ( n7171 , n7024 , n7170 );
and ( n7172 , n7021 , n7171 );
or ( n7173 , n7020 , n7172 );
and ( n7174 , n7017 , n7173 );
or ( n7175 , n7016 , n7174 );
and ( n7176 , n7013 , n7175 );
or ( n7177 , n7012 , n7176 );
and ( n7178 , n7009 , n7177 );
or ( n7179 , n7008 , n7178 );
and ( n7180 , n7005 , n7179 );
or ( n7181 , n7004 , n7180 );
xor ( n7182 , n7001 , n7181 );
and ( n7183 , n6983 , n6987 );
and ( n7184 , n6785 , n6981 );
and ( n7185 , n6981 , n6988 );
and ( n7186 , n6785 , n6988 );
or ( n7187 , n7184 , n7185 , n7186 );
xor ( n7188 , n7183 , n7187 );
and ( n7189 , n6789 , n6854 );
and ( n7190 , n6854 , n6980 );
and ( n7191 , n6789 , n6980 );
or ( n7192 , n7189 , n7190 , n7191 );
and ( n7193 , n6859 , n6908 );
and ( n7194 , n6908 , n6979 );
and ( n7195 , n6859 , n6979 );
or ( n7196 , n7193 , n7194 , n7195 );
and ( n7197 , n6913 , n6939 );
and ( n7198 , n6939 , n6978 );
and ( n7199 , n6913 , n6978 );
or ( n7200 , n7197 , n7198 , n7199 );
and ( n7201 , n6872 , n6888 );
and ( n7202 , n6888 , n6906 );
and ( n7203 , n6872 , n6906 );
or ( n7204 , n7201 , n7202 , n7203 );
and ( n7205 , n6917 , n6921 );
and ( n7206 , n6921 , n6938 );
and ( n7207 , n6917 , n6938 );
or ( n7208 , n7205 , n7206 , n7207 );
xor ( n7209 , n7204 , n7208 );
and ( n7210 , n6895 , n6899 );
and ( n7211 , n6899 , n6905 );
and ( n7212 , n6895 , n6905 );
or ( n7213 , n7210 , n7211 , n7212 );
and ( n7214 , n6883 , n6884 );
and ( n7215 , n6884 , n6886 );
and ( n7216 , n6883 , n6886 );
or ( n7217 , n7214 , n7215 , n7216 );
and ( n7218 , n3182 , n1424 );
and ( n7219 , n3545 , n1254 );
xor ( n7220 , n7218 , n7219 );
and ( n7221 , n3801 , n1134 );
xor ( n7222 , n7220 , n7221 );
xor ( n7223 , n7217 , n7222 );
and ( n7224 , n2462 , n1882 );
and ( n7225 , n2779 , n1738 );
xor ( n7226 , n7224 , n7225 );
and ( n7227 , n3024 , n1551 );
xor ( n7228 , n7226 , n7227 );
xor ( n7229 , n7223 , n7228 );
xor ( n7230 , n7213 , n7229 );
and ( n7231 , n6901 , n6902 );
and ( n7232 , n6902 , n6904 );
and ( n7233 , n6901 , n6904 );
or ( n7234 , n7231 , n7232 , n7233 );
and ( n7235 , n6927 , n6928 );
and ( n7236 , n6928 , n6930 );
and ( n7237 , n6927 , n6930 );
or ( n7238 , n7235 , n7236 , n7237 );
xor ( n7239 , n7234 , n7238 );
and ( n7240 , n1933 , n2544 );
and ( n7241 , n2120 , n2298 );
xor ( n7242 , n7240 , n7241 );
and ( n7243 , n2324 , n2100 );
xor ( n7244 , n7242 , n7243 );
xor ( n7245 , n7239 , n7244 );
xor ( n7246 , n7230 , n7245 );
xor ( n7247 , n7209 , n7246 );
xor ( n7248 , n7200 , n7247 );
and ( n7249 , n6944 , n6959 );
and ( n7250 , n6959 , n6977 );
and ( n7251 , n6944 , n6977 );
or ( n7252 , n7249 , n7250 , n7251 );
and ( n7253 , n6926 , n6931 );
and ( n7254 , n6931 , n6937 );
and ( n7255 , n6926 , n6937 );
or ( n7256 , n7253 , n7254 , n7255 );
and ( n7257 , n6948 , n6952 );
and ( n7258 , n6952 , n6958 );
and ( n7259 , n6948 , n6958 );
or ( n7260 , n7257 , n7258 , n7259 );
xor ( n7261 , n7256 , n7260 );
and ( n7262 , n6933 , n6934 );
and ( n7263 , n6934 , n6936 );
and ( n7264 , n6933 , n6936 );
or ( n7265 , n7262 , n7263 , n7264 );
and ( n7266 , n1383 , n3271 );
and ( n7267 , n1580 , n2981 );
xor ( n7268 , n7266 , n7267 );
and ( n7269 , n1694 , n2739 );
xor ( n7270 , n7268 , n7269 );
xor ( n7271 , n7265 , n7270 );
and ( n7272 , n1047 , n4102 );
and ( n7273 , n1164 , n3749 );
xor ( n7274 , n7272 , n7273 );
and ( n7275 , n1287 , n3495 );
xor ( n7276 , n7274 , n7275 );
xor ( n7277 , n7271 , n7276 );
xor ( n7278 , n7261 , n7277 );
xor ( n7279 , n7252 , n7278 );
and ( n7280 , n6964 , n6969 );
and ( n7281 , n6969 , n6976 );
and ( n7282 , n6964 , n6976 );
or ( n7283 , n7280 , n7281 , n7282 );
and ( n7284 , n6954 , n6955 );
and ( n7285 , n6955 , n6957 );
and ( n7286 , n6954 , n6957 );
or ( n7287 , n7284 , n7285 , n7286 );
and ( n7288 , n6965 , n6966 );
and ( n7289 , n6966 , n6968 );
and ( n7290 , n6965 , n6968 );
or ( n7291 , n7288 , n7289 , n7290 );
xor ( n7292 , n7287 , n7291 );
and ( n7293 , n783 , n5103 );
and ( n7294 , n856 , n4730 );
xor ( n7295 , n7293 , n7294 );
and ( n7296 , n925 , n4403 );
xor ( n7297 , n7295 , n7296 );
xor ( n7298 , n7292 , n7297 );
xor ( n7299 , n7283 , n7298 );
and ( n7300 , n6972 , n6973 );
and ( n7301 , n6973 , n6975 );
and ( n7302 , n6972 , n6975 );
or ( n7303 , n7300 , n7301 , n7302 );
and ( n7304 , n632 , n6132 );
and ( n7305 , n671 , n5765 );
xor ( n7306 , n7304 , n7305 );
and ( n7307 , n715 , n5408 );
xor ( n7308 , n7306 , n7307 );
xor ( n7309 , n7303 , n7308 );
buf ( n7310 , n437 );
and ( n7311 , n599 , n7310 );
and ( n7312 , n608 , n6971 );
xor ( n7313 , n7311 , n7312 );
and ( n7314 , n611 , n6504 );
xor ( n7315 , n7313 , n7314 );
xor ( n7316 , n7309 , n7315 );
xor ( n7317 , n7299 , n7316 );
xor ( n7318 , n7279 , n7317 );
xor ( n7319 , n7248 , n7318 );
xor ( n7320 , n7196 , n7319 );
and ( n7321 , n6802 , n6826 );
and ( n7322 , n6826 , n6852 );
and ( n7323 , n6802 , n6852 );
or ( n7324 , n7321 , n7322 , n7323 );
and ( n7325 , n6863 , n6867 );
and ( n7326 , n6867 , n6907 );
and ( n7327 , n6863 , n6907 );
or ( n7328 , n7325 , n7326 , n7327 );
xor ( n7329 , n7324 , n7328 );
and ( n7330 , n6831 , n6835 );
and ( n7331 , n6835 , n6851 );
and ( n7332 , n6831 , n6851 );
or ( n7333 , n7330 , n7331 , n7332 );
and ( n7334 , n6840 , n6844 );
and ( n7335 , n6844 , n6850 );
and ( n7336 , n6840 , n6850 );
or ( n7337 , n7334 , n7335 , n7336 );
and ( n7338 , n6876 , n6881 );
and ( n7339 , n6881 , n6887 );
and ( n7340 , n6876 , n6887 );
or ( n7341 , n7338 , n7339 , n7340 );
xor ( n7342 , n7337 , n7341 );
and ( n7343 , n6846 , n6847 );
and ( n7344 , n6847 , n6849 );
and ( n7345 , n6846 , n6849 );
or ( n7346 , n7343 , n7344 , n7345 );
and ( n7347 , n6877 , n6878 );
and ( n7348 , n6878 , n6880 );
and ( n7349 , n6877 , n6880 );
or ( n7350 , n7347 , n7348 , n7349 );
xor ( n7351 , n7346 , n7350 );
and ( n7352 , n4132 , n1034 );
and ( n7353 , n4438 , n940 );
xor ( n7354 , n7352 , n7353 );
and ( n7355 , n4766 , n840 );
xor ( n7356 , n7354 , n7355 );
xor ( n7357 , n7351 , n7356 );
xor ( n7358 , n7342 , n7357 );
xor ( n7359 , n7333 , n7358 );
and ( n7360 , n6812 , n6818 );
and ( n7361 , n6818 , n6824 );
and ( n7362 , n6812 , n6824 );
or ( n7363 , n7360 , n7361 , n7362 );
and ( n7364 , n6820 , n6821 );
and ( n7365 , n6821 , n6823 );
and ( n7366 , n6820 , n6823 );
or ( n7367 , n7364 , n7365 , n7366 );
and ( n7368 , n6187 , n635 );
and ( n7369 , n6569 , n606 );
xor ( n7370 , n7368 , n7369 );
and ( n7371 , n6816 , n615 );
xor ( n7372 , n7370 , n7371 );
xor ( n7373 , n7367 , n7372 );
and ( n7374 , n4959 , n771 );
and ( n7375 , n5459 , n719 );
xor ( n7376 , n7374 , n7375 );
and ( n7377 , n5819 , n663 );
xor ( n7378 , n7376 , n7377 );
xor ( n7379 , n7373 , n7378 );
xor ( n7380 , n7363 , n7379 );
and ( n7381 , n6813 , n6814 );
and ( n7382 , n6814 , n6817 );
and ( n7383 , n6813 , n6817 );
or ( n7384 , n7381 , n7382 , n7383 );
buf ( n7385 , n437 );
and ( n7386 , n7385 , n612 );
xor ( n7387 , n7384 , n7386 );
xor ( n7388 , n7380 , n7387 );
xor ( n7389 , n7359 , n7388 );
xor ( n7390 , n7329 , n7389 );
xor ( n7391 , n7320 , n7390 );
xor ( n7392 , n7192 , n7391 );
and ( n7393 , n6803 , n6807 );
and ( n7394 , n6807 , n6825 );
and ( n7395 , n6803 , n6825 );
or ( n7396 , n7393 , n7394 , n7395 );
and ( n7397 , n6793 , n6797 );
and ( n7398 , n6797 , n6853 );
and ( n7399 , n6793 , n6853 );
or ( n7400 , n7397 , n7398 , n7399 );
xor ( n7401 , n7396 , n7400 );
xor ( n7402 , n7392 , n7401 );
xor ( n7403 , n7188 , n7402 );
and ( n7404 , n6776 , n6780 );
and ( n7405 , n6780 , n6989 );
and ( n7406 , n6776 , n6989 );
or ( n7407 , n7404 , n7405 , n7406 );
xor ( n7408 , n7403 , n7407 );
and ( n7409 , n6990 , n6993 );
xor ( n7410 , n7408 , n7409 );
buf ( n7411 , n7410 );
buf ( n7412 , n7411 );
not ( n7413 , n7412 );
buf ( n7414 , n531 );
not ( n7415 , n7414 );
nor ( n7416 , n7413 , n7415 );
xor ( n7417 , n7182 , n7416 );
xor ( n7418 , n7005 , n7179 );
nor ( n7419 , n6997 , n7415 );
and ( n7420 , n7418 , n7419 );
xor ( n7421 , n7418 , n7419 );
xor ( n7422 , n7009 , n7177 );
nor ( n7423 , n6596 , n7415 );
and ( n7424 , n7422 , n7423 );
xor ( n7425 , n7422 , n7423 );
xor ( n7426 , n7013 , n7175 );
nor ( n7427 , n6212 , n7415 );
and ( n7428 , n7426 , n7427 );
xor ( n7429 , n7426 , n7427 );
xor ( n7430 , n7017 , n7173 );
nor ( n7431 , n5838 , n7415 );
and ( n7432 , n7430 , n7431 );
xor ( n7433 , n7430 , n7431 );
xor ( n7434 , n7021 , n7171 );
nor ( n7435 , n5477 , n7415 );
and ( n7436 , n7434 , n7435 );
xor ( n7437 , n7434 , n7435 );
xor ( n7438 , n7025 , n7169 );
nor ( n7439 , n5126 , n7415 );
and ( n7440 , n7438 , n7439 );
xor ( n7441 , n7438 , n7439 );
xor ( n7442 , n7029 , n7167 );
nor ( n7443 , n4786 , n7415 );
and ( n7444 , n7442 , n7443 );
xor ( n7445 , n7442 , n7443 );
xor ( n7446 , n7033 , n7165 );
nor ( n7447 , n4458 , n7415 );
and ( n7448 , n7446 , n7447 );
xor ( n7449 , n7446 , n7447 );
xor ( n7450 , n7037 , n7163 );
nor ( n7451 , n4151 , n7415 );
and ( n7452 , n7450 , n7451 );
xor ( n7453 , n7450 , n7451 );
xor ( n7454 , n7041 , n7161 );
nor ( n7455 , n3853 , n7415 );
and ( n7456 , n7454 , n7455 );
xor ( n7457 , n7454 , n7455 );
xor ( n7458 , n7045 , n7159 );
nor ( n7459 , n3570 , n7415 );
and ( n7460 , n7458 , n7459 );
xor ( n7461 , n7458 , n7459 );
xor ( n7462 , n7049 , n7157 );
nor ( n7463 , n3300 , n7415 );
and ( n7464 , n7462 , n7463 );
xor ( n7465 , n7462 , n7463 );
xor ( n7466 , n7053 , n7155 );
nor ( n7467 , n3043 , n7415 );
and ( n7468 , n7466 , n7467 );
xor ( n7469 , n7466 , n7467 );
xor ( n7470 , n7057 , n7153 );
nor ( n7471 , n2797 , n7415 );
and ( n7472 , n7470 , n7471 );
xor ( n7473 , n7470 , n7471 );
xor ( n7474 , n7061 , n7151 );
nor ( n7475 , n2566 , n7415 );
and ( n7476 , n7474 , n7475 );
xor ( n7477 , n7474 , n7475 );
xor ( n7478 , n7065 , n7149 );
nor ( n7479 , n2343 , n7415 );
and ( n7480 , n7478 , n7479 );
xor ( n7481 , n7478 , n7479 );
xor ( n7482 , n7069 , n7147 );
nor ( n7483 , n2137 , n7415 );
and ( n7484 , n7482 , n7483 );
xor ( n7485 , n7482 , n7483 );
xor ( n7486 , n7073 , n7145 );
nor ( n7487 , n1945 , n7415 );
and ( n7488 , n7486 , n7487 );
xor ( n7489 , n7486 , n7487 );
xor ( n7490 , n7077 , n7143 );
nor ( n7491 , n1766 , n7415 );
and ( n7492 , n7490 , n7491 );
xor ( n7493 , n7490 , n7491 );
xor ( n7494 , n7081 , n7141 );
nor ( n7495 , n1598 , n7415 );
and ( n7496 , n7494 , n7495 );
xor ( n7497 , n7494 , n7495 );
xor ( n7498 , n7085 , n7139 );
nor ( n7499 , n1445 , n7415 );
and ( n7500 , n7498 , n7499 );
xor ( n7501 , n7498 , n7499 );
xor ( n7502 , n7089 , n7137 );
nor ( n7503 , n1303 , n7415 );
and ( n7504 , n7502 , n7503 );
xor ( n7505 , n7502 , n7503 );
xor ( n7506 , n7093 , n7135 );
nor ( n7507 , n1176 , n7415 );
and ( n7508 , n7506 , n7507 );
xor ( n7509 , n7506 , n7507 );
xor ( n7510 , n7097 , n7133 );
nor ( n7511 , n1062 , n7415 );
and ( n7512 , n7510 , n7511 );
xor ( n7513 , n7510 , n7511 );
xor ( n7514 , n7101 , n7131 );
nor ( n7515 , n958 , n7415 );
and ( n7516 , n7514 , n7515 );
xor ( n7517 , n7514 , n7515 );
xor ( n7518 , n7105 , n7129 );
nor ( n7519 , n868 , n7415 );
and ( n7520 , n7518 , n7519 );
xor ( n7521 , n7518 , n7519 );
xor ( n7522 , n7109 , n7127 );
nor ( n7523 , n796 , n7415 );
and ( n7524 , n7522 , n7523 );
xor ( n7525 , n7522 , n7523 );
xor ( n7526 , n7113 , n7125 );
nor ( n7527 , n733 , n7415 );
and ( n7528 , n7526 , n7527 );
xor ( n7529 , n7526 , n7527 );
xor ( n7530 , n7118 , n7123 );
nor ( n7531 , n684 , n7415 );
and ( n7532 , n7530 , n7531 );
xor ( n7533 , n7530 , n7531 );
xor ( n7534 , n7120 , n7121 );
buf ( n7535 , n7534 );
nor ( n7536 , n646 , n7415 );
and ( n7537 , n7535 , n7536 );
xor ( n7538 , n7535 , n7536 );
nor ( n7539 , n601 , n6598 );
buf ( n7540 , n7539 );
nor ( n7541 , n622 , n7415 );
and ( n7542 , n7540 , n7541 );
buf ( n7543 , n7542 );
and ( n7544 , n7538 , n7543 );
or ( n7545 , n7537 , n7544 );
and ( n7546 , n7533 , n7545 );
or ( n7547 , n7532 , n7546 );
and ( n7548 , n7529 , n7547 );
or ( n7549 , n7528 , n7548 );
and ( n7550 , n7525 , n7549 );
or ( n7551 , n7524 , n7550 );
and ( n7552 , n7521 , n7551 );
or ( n7553 , n7520 , n7552 );
and ( n7554 , n7517 , n7553 );
or ( n7555 , n7516 , n7554 );
and ( n7556 , n7513 , n7555 );
or ( n7557 , n7512 , n7556 );
and ( n7558 , n7509 , n7557 );
or ( n7559 , n7508 , n7558 );
and ( n7560 , n7505 , n7559 );
or ( n7561 , n7504 , n7560 );
and ( n7562 , n7501 , n7561 );
or ( n7563 , n7500 , n7562 );
and ( n7564 , n7497 , n7563 );
or ( n7565 , n7496 , n7564 );
and ( n7566 , n7493 , n7565 );
or ( n7567 , n7492 , n7566 );
and ( n7568 , n7489 , n7567 );
or ( n7569 , n7488 , n7568 );
and ( n7570 , n7485 , n7569 );
or ( n7571 , n7484 , n7570 );
and ( n7572 , n7481 , n7571 );
or ( n7573 , n7480 , n7572 );
and ( n7574 , n7477 , n7573 );
or ( n7575 , n7476 , n7574 );
and ( n7576 , n7473 , n7575 );
or ( n7577 , n7472 , n7576 );
and ( n7578 , n7469 , n7577 );
or ( n7579 , n7468 , n7578 );
and ( n7580 , n7465 , n7579 );
or ( n7581 , n7464 , n7580 );
and ( n7582 , n7461 , n7581 );
or ( n7583 , n7460 , n7582 );
and ( n7584 , n7457 , n7583 );
or ( n7585 , n7456 , n7584 );
and ( n7586 , n7453 , n7585 );
or ( n7587 , n7452 , n7586 );
and ( n7588 , n7449 , n7587 );
or ( n7589 , n7448 , n7588 );
and ( n7590 , n7445 , n7589 );
or ( n7591 , n7444 , n7590 );
and ( n7592 , n7441 , n7591 );
or ( n7593 , n7440 , n7592 );
and ( n7594 , n7437 , n7593 );
or ( n7595 , n7436 , n7594 );
and ( n7596 , n7433 , n7595 );
or ( n7597 , n7432 , n7596 );
and ( n7598 , n7429 , n7597 );
or ( n7599 , n7428 , n7598 );
and ( n7600 , n7425 , n7599 );
or ( n7601 , n7424 , n7600 );
and ( n7602 , n7421 , n7601 );
or ( n7603 , n7420 , n7602 );
xor ( n7604 , n7417 , n7603 );
and ( n7605 , n7396 , n7400 );
and ( n7606 , n7192 , n7391 );
and ( n7607 , n7391 , n7401 );
and ( n7608 , n7192 , n7401 );
or ( n7609 , n7606 , n7607 , n7608 );
xor ( n7610 , n7605 , n7609 );
and ( n7611 , n7196 , n7319 );
and ( n7612 , n7319 , n7390 );
and ( n7613 , n7196 , n7390 );
or ( n7614 , n7611 , n7612 , n7613 );
and ( n7615 , n7200 , n7247 );
and ( n7616 , n7247 , n7318 );
and ( n7617 , n7200 , n7318 );
or ( n7618 , n7615 , n7616 , n7617 );
and ( n7619 , n7252 , n7278 );
and ( n7620 , n7278 , n7317 );
and ( n7621 , n7252 , n7317 );
or ( n7622 , n7619 , n7620 , n7621 );
and ( n7623 , n7283 , n7298 );
and ( n7624 , n7298 , n7316 );
and ( n7625 , n7283 , n7316 );
or ( n7626 , n7623 , n7624 , n7625 );
and ( n7627 , n7265 , n7270 );
and ( n7628 , n7270 , n7276 );
and ( n7629 , n7265 , n7276 );
or ( n7630 , n7627 , n7628 , n7629 );
and ( n7631 , n7287 , n7291 );
and ( n7632 , n7291 , n7297 );
and ( n7633 , n7287 , n7297 );
or ( n7634 , n7631 , n7632 , n7633 );
xor ( n7635 , n7630 , n7634 );
and ( n7636 , n7272 , n7273 );
and ( n7637 , n7273 , n7275 );
and ( n7638 , n7272 , n7275 );
or ( n7639 , n7636 , n7637 , n7638 );
and ( n7640 , n1383 , n3495 );
and ( n7641 , n1580 , n3271 );
xor ( n7642 , n7640 , n7641 );
and ( n7643 , n1694 , n2981 );
xor ( n7644 , n7642 , n7643 );
xor ( n7645 , n7639 , n7644 );
and ( n7646 , n1047 , n4403 );
and ( n7647 , n1164 , n4102 );
xor ( n7648 , n7646 , n7647 );
and ( n7649 , n1287 , n3749 );
xor ( n7650 , n7648 , n7649 );
xor ( n7651 , n7645 , n7650 );
xor ( n7652 , n7635 , n7651 );
xor ( n7653 , n7626 , n7652 );
and ( n7654 , n7303 , n7308 );
and ( n7655 , n7308 , n7315 );
and ( n7656 , n7303 , n7315 );
or ( n7657 , n7654 , n7655 , n7656 );
and ( n7658 , n7311 , n7312 );
and ( n7659 , n7312 , n7314 );
and ( n7660 , n7311 , n7314 );
or ( n7661 , n7658 , n7659 , n7660 );
buf ( n7662 , n436 );
and ( n7663 , n599 , n7662 );
and ( n7664 , n608 , n7310 );
xor ( n7665 , n7663 , n7664 );
and ( n7666 , n611 , n6971 );
xor ( n7667 , n7665 , n7666 );
xor ( n7668 , n7661 , n7667 );
and ( n7669 , n632 , n6504 );
and ( n7670 , n671 , n6132 );
xor ( n7671 , n7669 , n7670 );
and ( n7672 , n715 , n5765 );
xor ( n7673 , n7671 , n7672 );
xor ( n7674 , n7668 , n7673 );
xor ( n7675 , n7657 , n7674 );
and ( n7676 , n7293 , n7294 );
and ( n7677 , n7294 , n7296 );
and ( n7678 , n7293 , n7296 );
or ( n7679 , n7676 , n7677 , n7678 );
and ( n7680 , n7304 , n7305 );
and ( n7681 , n7305 , n7307 );
and ( n7682 , n7304 , n7307 );
or ( n7683 , n7680 , n7681 , n7682 );
xor ( n7684 , n7679 , n7683 );
and ( n7685 , n783 , n5408 );
and ( n7686 , n856 , n5103 );
xor ( n7687 , n7685 , n7686 );
and ( n7688 , n925 , n4730 );
xor ( n7689 , n7687 , n7688 );
xor ( n7690 , n7684 , n7689 );
xor ( n7691 , n7675 , n7690 );
xor ( n7692 , n7653 , n7691 );
xor ( n7693 , n7622 , n7692 );
and ( n7694 , n7213 , n7229 );
and ( n7695 , n7229 , n7245 );
and ( n7696 , n7213 , n7245 );
or ( n7697 , n7694 , n7695 , n7696 );
and ( n7698 , n7256 , n7260 );
and ( n7699 , n7260 , n7277 );
and ( n7700 , n7256 , n7277 );
or ( n7701 , n7698 , n7699 , n7700 );
xor ( n7702 , n7697 , n7701 );
and ( n7703 , n7234 , n7238 );
and ( n7704 , n7238 , n7244 );
and ( n7705 , n7234 , n7244 );
or ( n7706 , n7703 , n7704 , n7705 );
and ( n7707 , n7224 , n7225 );
and ( n7708 , n7225 , n7227 );
and ( n7709 , n7224 , n7227 );
or ( n7710 , n7707 , n7708 , n7709 );
and ( n7711 , n3182 , n1551 );
and ( n7712 , n3545 , n1424 );
xor ( n7713 , n7711 , n7712 );
and ( n7714 , n3801 , n1254 );
xor ( n7715 , n7713 , n7714 );
xor ( n7716 , n7710 , n7715 );
and ( n7717 , n2462 , n2100 );
and ( n7718 , n2779 , n1882 );
xor ( n7719 , n7717 , n7718 );
and ( n7720 , n3024 , n1738 );
xor ( n7721 , n7719 , n7720 );
xor ( n7722 , n7716 , n7721 );
xor ( n7723 , n7706 , n7722 );
and ( n7724 , n7240 , n7241 );
and ( n7725 , n7241 , n7243 );
and ( n7726 , n7240 , n7243 );
or ( n7727 , n7724 , n7725 , n7726 );
and ( n7728 , n7266 , n7267 );
and ( n7729 , n7267 , n7269 );
and ( n7730 , n7266 , n7269 );
or ( n7731 , n7728 , n7729 , n7730 );
xor ( n7732 , n7727 , n7731 );
and ( n7733 , n1933 , n2739 );
and ( n7734 , n2120 , n2544 );
xor ( n7735 , n7733 , n7734 );
buf ( n7736 , n2324 );
xor ( n7737 , n7735 , n7736 );
xor ( n7738 , n7732 , n7737 );
xor ( n7739 , n7723 , n7738 );
xor ( n7740 , n7702 , n7739 );
xor ( n7741 , n7693 , n7740 );
xor ( n7742 , n7618 , n7741 );
and ( n7743 , n7204 , n7208 );
and ( n7744 , n7208 , n7246 );
and ( n7745 , n7204 , n7246 );
or ( n7746 , n7743 , n7744 , n7745 );
and ( n7747 , n7333 , n7358 );
and ( n7748 , n7358 , n7388 );
and ( n7749 , n7333 , n7388 );
or ( n7750 , n7747 , n7748 , n7749 );
xor ( n7751 , n7746 , n7750 );
and ( n7752 , n7337 , n7341 );
and ( n7753 , n7341 , n7357 );
and ( n7754 , n7337 , n7357 );
or ( n7755 , n7752 , n7753 , n7754 );
and ( n7756 , n7346 , n7350 );
and ( n7757 , n7350 , n7356 );
and ( n7758 , n7346 , n7356 );
or ( n7759 , n7756 , n7757 , n7758 );
and ( n7760 , n7217 , n7222 );
and ( n7761 , n7222 , n7228 );
and ( n7762 , n7217 , n7228 );
or ( n7763 , n7760 , n7761 , n7762 );
xor ( n7764 , n7759 , n7763 );
and ( n7765 , n7352 , n7353 );
and ( n7766 , n7353 , n7355 );
and ( n7767 , n7352 , n7355 );
or ( n7768 , n7765 , n7766 , n7767 );
and ( n7769 , n7218 , n7219 );
and ( n7770 , n7219 , n7221 );
and ( n7771 , n7218 , n7221 );
or ( n7772 , n7769 , n7770 , n7771 );
xor ( n7773 , n7768 , n7772 );
and ( n7774 , n4132 , n1134 );
and ( n7775 , n4438 , n1034 );
xor ( n7776 , n7774 , n7775 );
and ( n7777 , n4766 , n940 );
xor ( n7778 , n7776 , n7777 );
xor ( n7779 , n7773 , n7778 );
xor ( n7780 , n7764 , n7779 );
xor ( n7781 , n7755 , n7780 );
and ( n7782 , n7367 , n7372 );
and ( n7783 , n7372 , n7378 );
and ( n7784 , n7367 , n7378 );
or ( n7785 , n7782 , n7783 , n7784 );
and ( n7786 , n7374 , n7375 );
and ( n7787 , n7375 , n7377 );
and ( n7788 , n7374 , n7377 );
or ( n7789 , n7786 , n7787 , n7788 );
and ( n7790 , n6187 , n663 );
and ( n7791 , n6569 , n635 );
xor ( n7792 , n7790 , n7791 );
and ( n7793 , n6816 , n606 );
xor ( n7794 , n7792 , n7793 );
xor ( n7795 , n7789 , n7794 );
and ( n7796 , n4959 , n840 );
and ( n7797 , n5459 , n771 );
xor ( n7798 , n7796 , n7797 );
and ( n7799 , n5819 , n719 );
xor ( n7800 , n7798 , n7799 );
xor ( n7801 , n7795 , n7800 );
xor ( n7802 , n7785 , n7801 );
and ( n7803 , n7368 , n7369 );
and ( n7804 , n7369 , n7371 );
and ( n7805 , n7368 , n7371 );
or ( n7806 , n7803 , n7804 , n7805 );
and ( n7807 , n7385 , n615 );
buf ( n7808 , n436 );
and ( n7809 , n7808 , n612 );
xor ( n7810 , n7807 , n7809 );
xor ( n7811 , n7806 , n7810 );
xor ( n7812 , n7802 , n7811 );
xor ( n7813 , n7781 , n7812 );
xor ( n7814 , n7751 , n7813 );
xor ( n7815 , n7742 , n7814 );
xor ( n7816 , n7614 , n7815 );
and ( n7817 , n7324 , n7328 );
and ( n7818 , n7328 , n7389 );
and ( n7819 , n7324 , n7389 );
or ( n7820 , n7817 , n7818 , n7819 );
and ( n7821 , n7384 , n7386 );
and ( n7822 , n7363 , n7379 );
and ( n7823 , n7379 , n7387 );
and ( n7824 , n7363 , n7387 );
or ( n7825 , n7822 , n7823 , n7824 );
xor ( n7826 , n7821 , n7825 );
xor ( n7827 , n7820 , n7826 );
xor ( n7828 , n7816 , n7827 );
xor ( n7829 , n7610 , n7828 );
and ( n7830 , n7183 , n7187 );
and ( n7831 , n7187 , n7402 );
and ( n7832 , n7183 , n7402 );
or ( n7833 , n7830 , n7831 , n7832 );
xor ( n7834 , n7829 , n7833 );
and ( n7835 , n7403 , n7407 );
and ( n7836 , n7408 , n7409 );
or ( n7837 , n7835 , n7836 );
xor ( n7838 , n7834 , n7837 );
buf ( n7839 , n7838 );
buf ( n7840 , n7839 );
not ( n7841 , n7840 );
buf ( n7842 , n532 );
not ( n7843 , n7842 );
nor ( n7844 , n7841 , n7843 );
xor ( n7845 , n7604 , n7844 );
xor ( n7846 , n7421 , n7601 );
nor ( n7847 , n7413 , n7843 );
and ( n7848 , n7846 , n7847 );
xor ( n7849 , n7846 , n7847 );
xor ( n7850 , n7425 , n7599 );
nor ( n7851 , n6997 , n7843 );
and ( n7852 , n7850 , n7851 );
xor ( n7853 , n7850 , n7851 );
xor ( n7854 , n7429 , n7597 );
nor ( n7855 , n6596 , n7843 );
and ( n7856 , n7854 , n7855 );
xor ( n7857 , n7854 , n7855 );
xor ( n7858 , n7433 , n7595 );
nor ( n7859 , n6212 , n7843 );
and ( n7860 , n7858 , n7859 );
xor ( n7861 , n7858 , n7859 );
xor ( n7862 , n7437 , n7593 );
nor ( n7863 , n5838 , n7843 );
and ( n7864 , n7862 , n7863 );
xor ( n7865 , n7862 , n7863 );
xor ( n7866 , n7441 , n7591 );
nor ( n7867 , n5477 , n7843 );
and ( n7868 , n7866 , n7867 );
xor ( n7869 , n7866 , n7867 );
xor ( n7870 , n7445 , n7589 );
nor ( n7871 , n5126 , n7843 );
and ( n7872 , n7870 , n7871 );
xor ( n7873 , n7870 , n7871 );
xor ( n7874 , n7449 , n7587 );
nor ( n7875 , n4786 , n7843 );
and ( n7876 , n7874 , n7875 );
xor ( n7877 , n7874 , n7875 );
xor ( n7878 , n7453 , n7585 );
nor ( n7879 , n4458 , n7843 );
and ( n7880 , n7878 , n7879 );
xor ( n7881 , n7878 , n7879 );
xor ( n7882 , n7457 , n7583 );
nor ( n7883 , n4151 , n7843 );
and ( n7884 , n7882 , n7883 );
xor ( n7885 , n7882 , n7883 );
xor ( n7886 , n7461 , n7581 );
nor ( n7887 , n3853 , n7843 );
and ( n7888 , n7886 , n7887 );
xor ( n7889 , n7886 , n7887 );
xor ( n7890 , n7465 , n7579 );
nor ( n7891 , n3570 , n7843 );
and ( n7892 , n7890 , n7891 );
xor ( n7893 , n7890 , n7891 );
xor ( n7894 , n7469 , n7577 );
nor ( n7895 , n3300 , n7843 );
and ( n7896 , n7894 , n7895 );
xor ( n7897 , n7894 , n7895 );
xor ( n7898 , n7473 , n7575 );
nor ( n7899 , n3043 , n7843 );
and ( n7900 , n7898 , n7899 );
xor ( n7901 , n7898 , n7899 );
xor ( n7902 , n7477 , n7573 );
nor ( n7903 , n2797 , n7843 );
and ( n7904 , n7902 , n7903 );
xor ( n7905 , n7902 , n7903 );
xor ( n7906 , n7481 , n7571 );
nor ( n7907 , n2566 , n7843 );
and ( n7908 , n7906 , n7907 );
xor ( n7909 , n7906 , n7907 );
xor ( n7910 , n7485 , n7569 );
nor ( n7911 , n2343 , n7843 );
and ( n7912 , n7910 , n7911 );
xor ( n7913 , n7910 , n7911 );
xor ( n7914 , n7489 , n7567 );
nor ( n7915 , n2137 , n7843 );
and ( n7916 , n7914 , n7915 );
xor ( n7917 , n7914 , n7915 );
xor ( n7918 , n7493 , n7565 );
nor ( n7919 , n1945 , n7843 );
and ( n7920 , n7918 , n7919 );
xor ( n7921 , n7918 , n7919 );
xor ( n7922 , n7497 , n7563 );
nor ( n7923 , n1766 , n7843 );
and ( n7924 , n7922 , n7923 );
xor ( n7925 , n7922 , n7923 );
xor ( n7926 , n7501 , n7561 );
nor ( n7927 , n1598 , n7843 );
and ( n7928 , n7926 , n7927 );
xor ( n7929 , n7926 , n7927 );
xor ( n7930 , n7505 , n7559 );
nor ( n7931 , n1445 , n7843 );
and ( n7932 , n7930 , n7931 );
xor ( n7933 , n7930 , n7931 );
xor ( n7934 , n7509 , n7557 );
nor ( n7935 , n1303 , n7843 );
and ( n7936 , n7934 , n7935 );
xor ( n7937 , n7934 , n7935 );
xor ( n7938 , n7513 , n7555 );
nor ( n7939 , n1176 , n7843 );
and ( n7940 , n7938 , n7939 );
xor ( n7941 , n7938 , n7939 );
xor ( n7942 , n7517 , n7553 );
nor ( n7943 , n1062 , n7843 );
and ( n7944 , n7942 , n7943 );
xor ( n7945 , n7942 , n7943 );
xor ( n7946 , n7521 , n7551 );
nor ( n7947 , n958 , n7843 );
and ( n7948 , n7946 , n7947 );
xor ( n7949 , n7946 , n7947 );
xor ( n7950 , n7525 , n7549 );
nor ( n7951 , n868 , n7843 );
and ( n7952 , n7950 , n7951 );
xor ( n7953 , n7950 , n7951 );
xor ( n7954 , n7529 , n7547 );
nor ( n7955 , n796 , n7843 );
and ( n7956 , n7954 , n7955 );
xor ( n7957 , n7954 , n7955 );
xor ( n7958 , n7533 , n7545 );
nor ( n7959 , n733 , n7843 );
and ( n7960 , n7958 , n7959 );
xor ( n7961 , n7958 , n7959 );
xor ( n7962 , n7538 , n7543 );
nor ( n7963 , n684 , n7843 );
and ( n7964 , n7962 , n7963 );
xor ( n7965 , n7962 , n7963 );
xor ( n7966 , n7540 , n7541 );
buf ( n7967 , n7966 );
nor ( n7968 , n646 , n7843 );
and ( n7969 , n7967 , n7968 );
xor ( n7970 , n7967 , n7968 );
nor ( n7971 , n601 , n6999 );
buf ( n7972 , n7971 );
nor ( n7973 , n622 , n7843 );
and ( n7974 , n7972 , n7973 );
buf ( n7975 , n7974 );
and ( n7976 , n7970 , n7975 );
or ( n7977 , n7969 , n7976 );
and ( n7978 , n7965 , n7977 );
or ( n7979 , n7964 , n7978 );
and ( n7980 , n7961 , n7979 );
or ( n7981 , n7960 , n7980 );
and ( n7982 , n7957 , n7981 );
or ( n7983 , n7956 , n7982 );
and ( n7984 , n7953 , n7983 );
or ( n7985 , n7952 , n7984 );
and ( n7986 , n7949 , n7985 );
or ( n7987 , n7948 , n7986 );
and ( n7988 , n7945 , n7987 );
or ( n7989 , n7944 , n7988 );
and ( n7990 , n7941 , n7989 );
or ( n7991 , n7940 , n7990 );
and ( n7992 , n7937 , n7991 );
or ( n7993 , n7936 , n7992 );
and ( n7994 , n7933 , n7993 );
or ( n7995 , n7932 , n7994 );
and ( n7996 , n7929 , n7995 );
or ( n7997 , n7928 , n7996 );
and ( n7998 , n7925 , n7997 );
or ( n7999 , n7924 , n7998 );
and ( n8000 , n7921 , n7999 );
or ( n8001 , n7920 , n8000 );
and ( n8002 , n7917 , n8001 );
or ( n8003 , n7916 , n8002 );
and ( n8004 , n7913 , n8003 );
or ( n8005 , n7912 , n8004 );
and ( n8006 , n7909 , n8005 );
or ( n8007 , n7908 , n8006 );
and ( n8008 , n7905 , n8007 );
or ( n8009 , n7904 , n8008 );
and ( n8010 , n7901 , n8009 );
or ( n8011 , n7900 , n8010 );
and ( n8012 , n7897 , n8011 );
or ( n8013 , n7896 , n8012 );
and ( n8014 , n7893 , n8013 );
or ( n8015 , n7892 , n8014 );
and ( n8016 , n7889 , n8015 );
or ( n8017 , n7888 , n8016 );
and ( n8018 , n7885 , n8017 );
or ( n8019 , n7884 , n8018 );
and ( n8020 , n7881 , n8019 );
or ( n8021 , n7880 , n8020 );
and ( n8022 , n7877 , n8021 );
or ( n8023 , n7876 , n8022 );
and ( n8024 , n7873 , n8023 );
or ( n8025 , n7872 , n8024 );
and ( n8026 , n7869 , n8025 );
or ( n8027 , n7868 , n8026 );
and ( n8028 , n7865 , n8027 );
or ( n8029 , n7864 , n8028 );
and ( n8030 , n7861 , n8029 );
or ( n8031 , n7860 , n8030 );
and ( n8032 , n7857 , n8031 );
or ( n8033 , n7856 , n8032 );
and ( n8034 , n7853 , n8033 );
or ( n8035 , n7852 , n8034 );
and ( n8036 , n7849 , n8035 );
or ( n8037 , n7848 , n8036 );
xor ( n8038 , n7845 , n8037 );
and ( n8039 , n7820 , n7826 );
and ( n8040 , n7614 , n7815 );
and ( n8041 , n7815 , n7827 );
and ( n8042 , n7614 , n7827 );
or ( n8043 , n8040 , n8041 , n8042 );
xor ( n8044 , n8039 , n8043 );
and ( n8045 , n7618 , n7741 );
and ( n8046 , n7741 , n7814 );
and ( n8047 , n7618 , n7814 );
or ( n8048 , n8045 , n8046 , n8047 );
and ( n8049 , n7622 , n7692 );
and ( n8050 , n7692 , n7740 );
and ( n8051 , n7622 , n7740 );
or ( n8052 , n8049 , n8050 , n8051 );
and ( n8053 , n7697 , n7701 );
and ( n8054 , n7701 , n7739 );
and ( n8055 , n7697 , n7739 );
or ( n8056 , n8053 , n8054 , n8055 );
and ( n8057 , n7755 , n7780 );
and ( n8058 , n7780 , n7812 );
and ( n8059 , n7755 , n7812 );
or ( n8060 , n8057 , n8058 , n8059 );
xor ( n8061 , n8056 , n8060 );
and ( n8062 , n7759 , n7763 );
and ( n8063 , n7763 , n7779 );
and ( n8064 , n7759 , n7779 );
or ( n8065 , n8062 , n8063 , n8064 );
and ( n8066 , n7789 , n7794 );
and ( n8067 , n7794 , n7800 );
and ( n8068 , n7789 , n7800 );
or ( n8069 , n8066 , n8067 , n8068 );
and ( n8070 , n7790 , n7791 );
and ( n8071 , n7791 , n7793 );
and ( n8072 , n7790 , n7793 );
or ( n8073 , n8070 , n8071 , n8072 );
and ( n8074 , n7807 , n7809 );
xor ( n8075 , n8073 , n8074 );
and ( n8076 , n7385 , n606 );
and ( n8077 , n7808 , n615 );
xor ( n8078 , n8076 , n8077 );
buf ( n8079 , n435 );
and ( n8080 , n8079 , n612 );
xor ( n8081 , n8078 , n8080 );
xor ( n8082 , n8075 , n8081 );
xor ( n8083 , n8069 , n8082 );
and ( n8084 , n7796 , n7797 );
and ( n8085 , n7797 , n7799 );
and ( n8086 , n7796 , n7799 );
or ( n8087 , n8084 , n8085 , n8086 );
and ( n8088 , n6187 , n719 );
and ( n8089 , n6569 , n663 );
xor ( n8090 , n8088 , n8089 );
and ( n8091 , n6816 , n635 );
xor ( n8092 , n8090 , n8091 );
xor ( n8093 , n8087 , n8092 );
and ( n8094 , n4959 , n940 );
and ( n8095 , n5459 , n840 );
xor ( n8096 , n8094 , n8095 );
and ( n8097 , n5819 , n771 );
xor ( n8098 , n8096 , n8097 );
xor ( n8099 , n8093 , n8098 );
xor ( n8100 , n8083 , n8099 );
xor ( n8101 , n8065 , n8100 );
and ( n8102 , n7710 , n7715 );
and ( n8103 , n7715 , n7721 );
and ( n8104 , n7710 , n7721 );
or ( n8105 , n8102 , n8103 , n8104 );
and ( n8106 , n7768 , n7772 );
and ( n8107 , n7772 , n7778 );
and ( n8108 , n7768 , n7778 );
or ( n8109 , n8106 , n8107 , n8108 );
xor ( n8110 , n8105 , n8109 );
and ( n8111 , n7774 , n7775 );
and ( n8112 , n7775 , n7777 );
and ( n8113 , n7774 , n7777 );
or ( n8114 , n8111 , n8112 , n8113 );
and ( n8115 , n7711 , n7712 );
and ( n8116 , n7712 , n7714 );
and ( n8117 , n7711 , n7714 );
or ( n8118 , n8115 , n8116 , n8117 );
xor ( n8119 , n8114 , n8118 );
and ( n8120 , n4132 , n1254 );
and ( n8121 , n4438 , n1134 );
xor ( n8122 , n8120 , n8121 );
and ( n8123 , n4766 , n1034 );
xor ( n8124 , n8122 , n8123 );
xor ( n8125 , n8119 , n8124 );
xor ( n8126 , n8110 , n8125 );
xor ( n8127 , n8101 , n8126 );
xor ( n8128 , n8061 , n8127 );
xor ( n8129 , n8052 , n8128 );
and ( n8130 , n7626 , n7652 );
and ( n8131 , n7652 , n7691 );
and ( n8132 , n7626 , n7691 );
or ( n8133 , n8130 , n8131 , n8132 );
and ( n8134 , n7630 , n7634 );
and ( n8135 , n7634 , n7651 );
and ( n8136 , n7630 , n7651 );
or ( n8137 , n8134 , n8135 , n8136 );
and ( n8138 , n7706 , n7722 );
and ( n8139 , n7722 , n7738 );
and ( n8140 , n7706 , n7738 );
or ( n8141 , n8138 , n8139 , n8140 );
xor ( n8142 , n8137 , n8141 );
and ( n8143 , n7727 , n7731 );
and ( n8144 , n7731 , n7737 );
and ( n8145 , n7727 , n7737 );
or ( n8146 , n8143 , n8144 , n8145 );
and ( n8147 , n7717 , n7718 );
and ( n8148 , n7718 , n7720 );
and ( n8149 , n7717 , n7720 );
or ( n8150 , n8147 , n8148 , n8149 );
and ( n8151 , n3182 , n1738 );
and ( n8152 , n3545 , n1551 );
xor ( n8153 , n8151 , n8152 );
and ( n8154 , n3801 , n1424 );
xor ( n8155 , n8153 , n8154 );
xor ( n8156 , n8150 , n8155 );
and ( n8157 , n2462 , n2298 );
and ( n8158 , n2779 , n2100 );
xor ( n8159 , n8157 , n8158 );
and ( n8160 , n3024 , n1882 );
xor ( n8161 , n8159 , n8160 );
xor ( n8162 , n8156 , n8161 );
xor ( n8163 , n8146 , n8162 );
and ( n8164 , n7733 , n7734 );
and ( n8165 , n7734 , n7736 );
and ( n8166 , n7733 , n7736 );
or ( n8167 , n8164 , n8165 , n8166 );
and ( n8168 , n7640 , n7641 );
and ( n8169 , n7641 , n7643 );
and ( n8170 , n7640 , n7643 );
or ( n8171 , n8168 , n8169 , n8170 );
xor ( n8172 , n8167 , n8171 );
and ( n8173 , n1933 , n2981 );
and ( n8174 , n2120 , n2739 );
xor ( n8175 , n8173 , n8174 );
and ( n8176 , n2324 , n2544 );
xor ( n8177 , n8175 , n8176 );
xor ( n8178 , n8172 , n8177 );
xor ( n8179 , n8163 , n8178 );
xor ( n8180 , n8142 , n8179 );
xor ( n8181 , n8133 , n8180 );
and ( n8182 , n7657 , n7674 );
and ( n8183 , n7674 , n7690 );
and ( n8184 , n7657 , n7690 );
or ( n8185 , n8182 , n8183 , n8184 );
and ( n8186 , n7679 , n7683 );
and ( n8187 , n7683 , n7689 );
and ( n8188 , n7679 , n7689 );
or ( n8189 , n8186 , n8187 , n8188 );
and ( n8190 , n7639 , n7644 );
and ( n8191 , n7644 , n7650 );
and ( n8192 , n7639 , n7650 );
or ( n8193 , n8190 , n8191 , n8192 );
xor ( n8194 , n8189 , n8193 );
and ( n8195 , n7646 , n7647 );
and ( n8196 , n7647 , n7649 );
and ( n8197 , n7646 , n7649 );
or ( n8198 , n8195 , n8196 , n8197 );
and ( n8199 , n1383 , n3749 );
and ( n8200 , n1580 , n3495 );
xor ( n8201 , n8199 , n8200 );
and ( n8202 , n1694 , n3271 );
xor ( n8203 , n8201 , n8202 );
xor ( n8204 , n8198 , n8203 );
and ( n8205 , n1047 , n4730 );
and ( n8206 , n1164 , n4403 );
xor ( n8207 , n8205 , n8206 );
and ( n8208 , n1287 , n4102 );
xor ( n8209 , n8207 , n8208 );
xor ( n8210 , n8204 , n8209 );
xor ( n8211 , n8194 , n8210 );
xor ( n8212 , n8185 , n8211 );
and ( n8213 , n7661 , n7667 );
and ( n8214 , n7667 , n7673 );
and ( n8215 , n7661 , n7673 );
or ( n8216 , n8213 , n8214 , n8215 );
and ( n8217 , n7669 , n7670 );
and ( n8218 , n7670 , n7672 );
and ( n8219 , n7669 , n7672 );
or ( n8220 , n8217 , n8218 , n8219 );
and ( n8221 , n7685 , n7686 );
and ( n8222 , n7686 , n7688 );
and ( n8223 , n7685 , n7688 );
or ( n8224 , n8221 , n8222 , n8223 );
xor ( n8225 , n8220 , n8224 );
and ( n8226 , n783 , n5765 );
and ( n8227 , n856 , n5408 );
xor ( n8228 , n8226 , n8227 );
and ( n8229 , n925 , n5103 );
xor ( n8230 , n8228 , n8229 );
xor ( n8231 , n8225 , n8230 );
xor ( n8232 , n8216 , n8231 );
and ( n8233 , n7663 , n7664 );
and ( n8234 , n7664 , n7666 );
and ( n8235 , n7663 , n7666 );
or ( n8236 , n8233 , n8234 , n8235 );
and ( n8237 , n632 , n6971 );
and ( n8238 , n671 , n6504 );
xor ( n8239 , n8237 , n8238 );
and ( n8240 , n715 , n6132 );
xor ( n8241 , n8239 , n8240 );
xor ( n8242 , n8236 , n8241 );
buf ( n8243 , n435 );
and ( n8244 , n599 , n8243 );
and ( n8245 , n608 , n7662 );
xor ( n8246 , n8244 , n8245 );
and ( n8247 , n611 , n7310 );
xor ( n8248 , n8246 , n8247 );
xor ( n8249 , n8242 , n8248 );
xor ( n8250 , n8232 , n8249 );
xor ( n8251 , n8212 , n8250 );
xor ( n8252 , n8181 , n8251 );
xor ( n8253 , n8129 , n8252 );
xor ( n8254 , n8048 , n8253 );
and ( n8255 , n7746 , n7750 );
and ( n8256 , n7750 , n7813 );
and ( n8257 , n7746 , n7813 );
or ( n8258 , n8255 , n8256 , n8257 );
and ( n8259 , n7821 , n7825 );
and ( n8260 , n7806 , n7810 );
and ( n8261 , n7785 , n7801 );
and ( n8262 , n7801 , n7811 );
and ( n8263 , n7785 , n7811 );
or ( n8264 , n8261 , n8262 , n8263 );
xor ( n8265 , n8260 , n8264 );
xor ( n8266 , n8259 , n8265 );
xor ( n8267 , n8258 , n8266 );
xor ( n8268 , n8254 , n8267 );
xor ( n8269 , n8044 , n8268 );
and ( n8270 , n7605 , n7609 );
and ( n8271 , n7609 , n7828 );
and ( n8272 , n7605 , n7828 );
or ( n8273 , n8270 , n8271 , n8272 );
xor ( n8274 , n8269 , n8273 );
and ( n8275 , n7829 , n7833 );
and ( n8276 , n7834 , n7837 );
or ( n8277 , n8275 , n8276 );
xor ( n8278 , n8274 , n8277 );
buf ( n8279 , n8278 );
buf ( n8280 , n8279 );
not ( n8281 , n8280 );
buf ( n8282 , n533 );
not ( n8283 , n8282 );
nor ( n8284 , n8281 , n8283 );
xor ( n8285 , n8038 , n8284 );
xor ( n8286 , n7849 , n8035 );
nor ( n8287 , n7841 , n8283 );
and ( n8288 , n8286 , n8287 );
xor ( n8289 , n8286 , n8287 );
xor ( n8290 , n7853 , n8033 );
nor ( n8291 , n7413 , n8283 );
and ( n8292 , n8290 , n8291 );
xor ( n8293 , n8290 , n8291 );
xor ( n8294 , n7857 , n8031 );
nor ( n8295 , n6997 , n8283 );
and ( n8296 , n8294 , n8295 );
xor ( n8297 , n8294 , n8295 );
xor ( n8298 , n7861 , n8029 );
nor ( n8299 , n6596 , n8283 );
and ( n8300 , n8298 , n8299 );
xor ( n8301 , n8298 , n8299 );
xor ( n8302 , n7865 , n8027 );
nor ( n8303 , n6212 , n8283 );
and ( n8304 , n8302 , n8303 );
xor ( n8305 , n8302 , n8303 );
xor ( n8306 , n7869 , n8025 );
nor ( n8307 , n5838 , n8283 );
and ( n8308 , n8306 , n8307 );
xor ( n8309 , n8306 , n8307 );
xor ( n8310 , n7873 , n8023 );
nor ( n8311 , n5477 , n8283 );
and ( n8312 , n8310 , n8311 );
xor ( n8313 , n8310 , n8311 );
xor ( n8314 , n7877 , n8021 );
nor ( n8315 , n5126 , n8283 );
and ( n8316 , n8314 , n8315 );
xor ( n8317 , n8314 , n8315 );
xor ( n8318 , n7881 , n8019 );
nor ( n8319 , n4786 , n8283 );
and ( n8320 , n8318 , n8319 );
xor ( n8321 , n8318 , n8319 );
xor ( n8322 , n7885 , n8017 );
nor ( n8323 , n4458 , n8283 );
and ( n8324 , n8322 , n8323 );
xor ( n8325 , n8322 , n8323 );
xor ( n8326 , n7889 , n8015 );
nor ( n8327 , n4151 , n8283 );
and ( n8328 , n8326 , n8327 );
xor ( n8329 , n8326 , n8327 );
xor ( n8330 , n7893 , n8013 );
nor ( n8331 , n3853 , n8283 );
and ( n8332 , n8330 , n8331 );
xor ( n8333 , n8330 , n8331 );
xor ( n8334 , n7897 , n8011 );
nor ( n8335 , n3570 , n8283 );
and ( n8336 , n8334 , n8335 );
xor ( n8337 , n8334 , n8335 );
xor ( n8338 , n7901 , n8009 );
nor ( n8339 , n3300 , n8283 );
and ( n8340 , n8338 , n8339 );
xor ( n8341 , n8338 , n8339 );
xor ( n8342 , n7905 , n8007 );
nor ( n8343 , n3043 , n8283 );
and ( n8344 , n8342 , n8343 );
xor ( n8345 , n8342 , n8343 );
xor ( n8346 , n7909 , n8005 );
nor ( n8347 , n2797 , n8283 );
and ( n8348 , n8346 , n8347 );
xor ( n8349 , n8346 , n8347 );
xor ( n8350 , n7913 , n8003 );
nor ( n8351 , n2566 , n8283 );
and ( n8352 , n8350 , n8351 );
xor ( n8353 , n8350 , n8351 );
xor ( n8354 , n7917 , n8001 );
nor ( n8355 , n2343 , n8283 );
and ( n8356 , n8354 , n8355 );
xor ( n8357 , n8354 , n8355 );
xor ( n8358 , n7921 , n7999 );
nor ( n8359 , n2137 , n8283 );
and ( n8360 , n8358 , n8359 );
xor ( n8361 , n8358 , n8359 );
xor ( n8362 , n7925 , n7997 );
nor ( n8363 , n1945 , n8283 );
and ( n8364 , n8362 , n8363 );
xor ( n8365 , n8362 , n8363 );
xor ( n8366 , n7929 , n7995 );
nor ( n8367 , n1766 , n8283 );
and ( n8368 , n8366 , n8367 );
xor ( n8369 , n8366 , n8367 );
xor ( n8370 , n7933 , n7993 );
nor ( n8371 , n1598 , n8283 );
and ( n8372 , n8370 , n8371 );
xor ( n8373 , n8370 , n8371 );
xor ( n8374 , n7937 , n7991 );
nor ( n8375 , n1445 , n8283 );
and ( n8376 , n8374 , n8375 );
xor ( n8377 , n8374 , n8375 );
xor ( n8378 , n7941 , n7989 );
nor ( n8379 , n1303 , n8283 );
and ( n8380 , n8378 , n8379 );
xor ( n8381 , n8378 , n8379 );
xor ( n8382 , n7945 , n7987 );
nor ( n8383 , n1176 , n8283 );
and ( n8384 , n8382 , n8383 );
xor ( n8385 , n8382 , n8383 );
xor ( n8386 , n7949 , n7985 );
nor ( n8387 , n1062 , n8283 );
and ( n8388 , n8386 , n8387 );
xor ( n8389 , n8386 , n8387 );
xor ( n8390 , n7953 , n7983 );
nor ( n8391 , n958 , n8283 );
and ( n8392 , n8390 , n8391 );
xor ( n8393 , n8390 , n8391 );
xor ( n8394 , n7957 , n7981 );
nor ( n8395 , n868 , n8283 );
and ( n8396 , n8394 , n8395 );
xor ( n8397 , n8394 , n8395 );
xor ( n8398 , n7961 , n7979 );
nor ( n8399 , n796 , n8283 );
and ( n8400 , n8398 , n8399 );
xor ( n8401 , n8398 , n8399 );
xor ( n8402 , n7965 , n7977 );
nor ( n8403 , n733 , n8283 );
and ( n8404 , n8402 , n8403 );
xor ( n8405 , n8402 , n8403 );
xor ( n8406 , n7970 , n7975 );
nor ( n8407 , n684 , n8283 );
and ( n8408 , n8406 , n8407 );
xor ( n8409 , n8406 , n8407 );
xor ( n8410 , n7972 , n7973 );
buf ( n8411 , n8410 );
nor ( n8412 , n646 , n8283 );
and ( n8413 , n8411 , n8412 );
xor ( n8414 , n8411 , n8412 );
nor ( n8415 , n601 , n7415 );
buf ( n8416 , n8415 );
nor ( n8417 , n622 , n8283 );
and ( n8418 , n8416 , n8417 );
buf ( n8419 , n8418 );
and ( n8420 , n8414 , n8419 );
or ( n8421 , n8413 , n8420 );
and ( n8422 , n8409 , n8421 );
or ( n8423 , n8408 , n8422 );
and ( n8424 , n8405 , n8423 );
or ( n8425 , n8404 , n8424 );
and ( n8426 , n8401 , n8425 );
or ( n8427 , n8400 , n8426 );
and ( n8428 , n8397 , n8427 );
or ( n8429 , n8396 , n8428 );
and ( n8430 , n8393 , n8429 );
or ( n8431 , n8392 , n8430 );
and ( n8432 , n8389 , n8431 );
or ( n8433 , n8388 , n8432 );
and ( n8434 , n8385 , n8433 );
or ( n8435 , n8384 , n8434 );
and ( n8436 , n8381 , n8435 );
or ( n8437 , n8380 , n8436 );
and ( n8438 , n8377 , n8437 );
or ( n8439 , n8376 , n8438 );
and ( n8440 , n8373 , n8439 );
or ( n8441 , n8372 , n8440 );
and ( n8442 , n8369 , n8441 );
or ( n8443 , n8368 , n8442 );
and ( n8444 , n8365 , n8443 );
or ( n8445 , n8364 , n8444 );
and ( n8446 , n8361 , n8445 );
or ( n8447 , n8360 , n8446 );
and ( n8448 , n8357 , n8447 );
or ( n8449 , n8356 , n8448 );
and ( n8450 , n8353 , n8449 );
or ( n8451 , n8352 , n8450 );
and ( n8452 , n8349 , n8451 );
or ( n8453 , n8348 , n8452 );
and ( n8454 , n8345 , n8453 );
or ( n8455 , n8344 , n8454 );
and ( n8456 , n8341 , n8455 );
or ( n8457 , n8340 , n8456 );
and ( n8458 , n8337 , n8457 );
or ( n8459 , n8336 , n8458 );
and ( n8460 , n8333 , n8459 );
or ( n8461 , n8332 , n8460 );
and ( n8462 , n8329 , n8461 );
or ( n8463 , n8328 , n8462 );
and ( n8464 , n8325 , n8463 );
or ( n8465 , n8324 , n8464 );
and ( n8466 , n8321 , n8465 );
or ( n8467 , n8320 , n8466 );
and ( n8468 , n8317 , n8467 );
or ( n8469 , n8316 , n8468 );
and ( n8470 , n8313 , n8469 );
or ( n8471 , n8312 , n8470 );
and ( n8472 , n8309 , n8471 );
or ( n8473 , n8308 , n8472 );
and ( n8474 , n8305 , n8473 );
or ( n8475 , n8304 , n8474 );
and ( n8476 , n8301 , n8475 );
or ( n8477 , n8300 , n8476 );
and ( n8478 , n8297 , n8477 );
or ( n8479 , n8296 , n8478 );
and ( n8480 , n8293 , n8479 );
or ( n8481 , n8292 , n8480 );
and ( n8482 , n8289 , n8481 );
or ( n8483 , n8288 , n8482 );
xor ( n8484 , n8285 , n8483 );
and ( n8485 , n8258 , n8266 );
and ( n8486 , n8048 , n8253 );
and ( n8487 , n8253 , n8267 );
and ( n8488 , n8048 , n8267 );
or ( n8489 , n8486 , n8487 , n8488 );
xor ( n8490 , n8485 , n8489 );
and ( n8491 , n8052 , n8128 );
and ( n8492 , n8128 , n8252 );
and ( n8493 , n8052 , n8252 );
or ( n8494 , n8491 , n8492 , n8493 );
and ( n8495 , n8133 , n8180 );
and ( n8496 , n8180 , n8251 );
and ( n8497 , n8133 , n8251 );
or ( n8498 , n8495 , n8496 , n8497 );
and ( n8499 , n8065 , n8100 );
and ( n8500 , n8100 , n8126 );
and ( n8501 , n8065 , n8126 );
or ( n8502 , n8499 , n8500 , n8501 );
and ( n8503 , n8137 , n8141 );
and ( n8504 , n8141 , n8179 );
and ( n8505 , n8137 , n8179 );
or ( n8506 , n8503 , n8504 , n8505 );
xor ( n8507 , n8502 , n8506 );
and ( n8508 , n8105 , n8109 );
and ( n8509 , n8109 , n8125 );
and ( n8510 , n8105 , n8125 );
or ( n8511 , n8508 , n8509 , n8510 );
and ( n8512 , n8087 , n8092 );
and ( n8513 , n8092 , n8098 );
and ( n8514 , n8087 , n8098 );
or ( n8515 , n8512 , n8513 , n8514 );
and ( n8516 , n8076 , n8077 );
and ( n8517 , n8077 , n8080 );
and ( n8518 , n8076 , n8080 );
or ( n8519 , n8516 , n8517 , n8518 );
and ( n8520 , n8088 , n8089 );
and ( n8521 , n8089 , n8091 );
and ( n8522 , n8088 , n8091 );
or ( n8523 , n8520 , n8521 , n8522 );
xor ( n8524 , n8519 , n8523 );
and ( n8525 , n7385 , n635 );
and ( n8526 , n7808 , n606 );
xor ( n8527 , n8525 , n8526 );
and ( n8528 , n8079 , n615 );
xor ( n8529 , n8527 , n8528 );
xor ( n8530 , n8524 , n8529 );
xor ( n8531 , n8515 , n8530 );
and ( n8532 , n8094 , n8095 );
and ( n8533 , n8095 , n8097 );
and ( n8534 , n8094 , n8097 );
or ( n8535 , n8532 , n8533 , n8534 );
and ( n8536 , n6187 , n771 );
and ( n8537 , n6569 , n719 );
xor ( n8538 , n8536 , n8537 );
and ( n8539 , n6816 , n663 );
xor ( n8540 , n8538 , n8539 );
xor ( n8541 , n8535 , n8540 );
and ( n8542 , n4959 , n1034 );
and ( n8543 , n5459 , n940 );
xor ( n8544 , n8542 , n8543 );
and ( n8545 , n5819 , n840 );
xor ( n8546 , n8544 , n8545 );
xor ( n8547 , n8541 , n8546 );
xor ( n8548 , n8531 , n8547 );
xor ( n8549 , n8511 , n8548 );
and ( n8550 , n8114 , n8118 );
and ( n8551 , n8118 , n8124 );
and ( n8552 , n8114 , n8124 );
or ( n8553 , n8550 , n8551 , n8552 );
and ( n8554 , n8150 , n8155 );
and ( n8555 , n8155 , n8161 );
and ( n8556 , n8150 , n8161 );
or ( n8557 , n8554 , n8555 , n8556 );
xor ( n8558 , n8553 , n8557 );
and ( n8559 , n8120 , n8121 );
and ( n8560 , n8121 , n8123 );
and ( n8561 , n8120 , n8123 );
or ( n8562 , n8559 , n8560 , n8561 );
and ( n8563 , n8151 , n8152 );
and ( n8564 , n8152 , n8154 );
and ( n8565 , n8151 , n8154 );
or ( n8566 , n8563 , n8564 , n8565 );
xor ( n8567 , n8562 , n8566 );
and ( n8568 , n4132 , n1424 );
and ( n8569 , n4438 , n1254 );
xor ( n8570 , n8568 , n8569 );
and ( n8571 , n4766 , n1134 );
xor ( n8572 , n8570 , n8571 );
xor ( n8573 , n8567 , n8572 );
xor ( n8574 , n8558 , n8573 );
xor ( n8575 , n8549 , n8574 );
xor ( n8576 , n8507 , n8575 );
xor ( n8577 , n8498 , n8576 );
and ( n8578 , n8185 , n8211 );
and ( n8579 , n8211 , n8250 );
and ( n8580 , n8185 , n8250 );
or ( n8581 , n8578 , n8579 , n8580 );
and ( n8582 , n8146 , n8162 );
and ( n8583 , n8162 , n8178 );
and ( n8584 , n8146 , n8178 );
or ( n8585 , n8582 , n8583 , n8584 );
and ( n8586 , n8189 , n8193 );
and ( n8587 , n8193 , n8210 );
and ( n8588 , n8189 , n8210 );
or ( n8589 , n8586 , n8587 , n8588 );
xor ( n8590 , n8585 , n8589 );
and ( n8591 , n8167 , n8171 );
and ( n8592 , n8171 , n8177 );
and ( n8593 , n8167 , n8177 );
or ( n8594 , n8591 , n8592 , n8593 );
and ( n8595 , n8157 , n8158 );
and ( n8596 , n8158 , n8160 );
and ( n8597 , n8157 , n8160 );
or ( n8598 , n8595 , n8596 , n8597 );
and ( n8599 , n3182 , n1882 );
and ( n8600 , n3545 , n1738 );
xor ( n8601 , n8599 , n8600 );
and ( n8602 , n3801 , n1551 );
xor ( n8603 , n8601 , n8602 );
xor ( n8604 , n8598 , n8603 );
buf ( n8605 , n2462 );
and ( n8606 , n2779 , n2298 );
xor ( n8607 , n8605 , n8606 );
and ( n8608 , n3024 , n2100 );
xor ( n8609 , n8607 , n8608 );
xor ( n8610 , n8604 , n8609 );
xor ( n8611 , n8594 , n8610 );
and ( n8612 , n8173 , n8174 );
and ( n8613 , n8174 , n8176 );
and ( n8614 , n8173 , n8176 );
or ( n8615 , n8612 , n8613 , n8614 );
and ( n8616 , n8199 , n8200 );
and ( n8617 , n8200 , n8202 );
and ( n8618 , n8199 , n8202 );
or ( n8619 , n8616 , n8617 , n8618 );
xor ( n8620 , n8615 , n8619 );
and ( n8621 , n1933 , n3271 );
and ( n8622 , n2120 , n2981 );
xor ( n8623 , n8621 , n8622 );
and ( n8624 , n2324 , n2739 );
xor ( n8625 , n8623 , n8624 );
xor ( n8626 , n8620 , n8625 );
xor ( n8627 , n8611 , n8626 );
xor ( n8628 , n8590 , n8627 );
xor ( n8629 , n8581 , n8628 );
and ( n8630 , n8216 , n8231 );
and ( n8631 , n8231 , n8249 );
and ( n8632 , n8216 , n8249 );
or ( n8633 , n8630 , n8631 , n8632 );
and ( n8634 , n8198 , n8203 );
and ( n8635 , n8203 , n8209 );
and ( n8636 , n8198 , n8209 );
or ( n8637 , n8634 , n8635 , n8636 );
and ( n8638 , n8220 , n8224 );
and ( n8639 , n8224 , n8230 );
and ( n8640 , n8220 , n8230 );
or ( n8641 , n8638 , n8639 , n8640 );
xor ( n8642 , n8637 , n8641 );
and ( n8643 , n8205 , n8206 );
and ( n8644 , n8206 , n8208 );
and ( n8645 , n8205 , n8208 );
or ( n8646 , n8643 , n8644 , n8645 );
and ( n8647 , n1383 , n4102 );
and ( n8648 , n1580 , n3749 );
xor ( n8649 , n8647 , n8648 );
and ( n8650 , n1694 , n3495 );
xor ( n8651 , n8649 , n8650 );
xor ( n8652 , n8646 , n8651 );
and ( n8653 , n1047 , n5103 );
and ( n8654 , n1164 , n4730 );
xor ( n8655 , n8653 , n8654 );
and ( n8656 , n1287 , n4403 );
xor ( n8657 , n8655 , n8656 );
xor ( n8658 , n8652 , n8657 );
xor ( n8659 , n8642 , n8658 );
xor ( n8660 , n8633 , n8659 );
and ( n8661 , n8236 , n8241 );
and ( n8662 , n8241 , n8248 );
and ( n8663 , n8236 , n8248 );
or ( n8664 , n8661 , n8662 , n8663 );
and ( n8665 , n8244 , n8245 );
and ( n8666 , n8245 , n8247 );
and ( n8667 , n8244 , n8247 );
or ( n8668 , n8665 , n8666 , n8667 );
buf ( n8669 , n434 );
and ( n8670 , n599 , n8669 );
and ( n8671 , n608 , n8243 );
xor ( n8672 , n8670 , n8671 );
and ( n8673 , n611 , n7662 );
xor ( n8674 , n8672 , n8673 );
xor ( n8675 , n8668 , n8674 );
and ( n8676 , n632 , n7310 );
and ( n8677 , n671 , n6971 );
xor ( n8678 , n8676 , n8677 );
and ( n8679 , n715 , n6504 );
xor ( n8680 , n8678 , n8679 );
xor ( n8681 , n8675 , n8680 );
xor ( n8682 , n8664 , n8681 );
and ( n8683 , n8226 , n8227 );
and ( n8684 , n8227 , n8229 );
and ( n8685 , n8226 , n8229 );
or ( n8686 , n8683 , n8684 , n8685 );
and ( n8687 , n8237 , n8238 );
and ( n8688 , n8238 , n8240 );
and ( n8689 , n8237 , n8240 );
or ( n8690 , n8687 , n8688 , n8689 );
xor ( n8691 , n8686 , n8690 );
and ( n8692 , n783 , n6132 );
and ( n8693 , n856 , n5765 );
xor ( n8694 , n8692 , n8693 );
and ( n8695 , n925 , n5408 );
xor ( n8696 , n8694 , n8695 );
xor ( n8697 , n8691 , n8696 );
xor ( n8698 , n8682 , n8697 );
xor ( n8699 , n8660 , n8698 );
xor ( n8700 , n8629 , n8699 );
xor ( n8701 , n8577 , n8700 );
xor ( n8702 , n8494 , n8701 );
and ( n8703 , n8056 , n8060 );
and ( n8704 , n8060 , n8127 );
and ( n8705 , n8056 , n8127 );
or ( n8706 , n8703 , n8704 , n8705 );
and ( n8707 , n8259 , n8265 );
xor ( n8708 , n8706 , n8707 );
and ( n8709 , n8260 , n8264 );
and ( n8710 , n8069 , n8082 );
and ( n8711 , n8082 , n8099 );
and ( n8712 , n8069 , n8099 );
or ( n8713 , n8710 , n8711 , n8712 );
and ( n8714 , n8073 , n8074 );
and ( n8715 , n8074 , n8081 );
and ( n8716 , n8073 , n8081 );
or ( n8717 , n8714 , n8715 , n8716 );
buf ( n8718 , n434 );
and ( n8719 , n8718 , n612 );
xor ( n8720 , n8717 , n8719 );
xor ( n8721 , n8713 , n8720 );
xor ( n8722 , n8709 , n8721 );
xor ( n8723 , n8708 , n8722 );
xor ( n8724 , n8702 , n8723 );
xor ( n8725 , n8490 , n8724 );
and ( n8726 , n8039 , n8043 );
and ( n8727 , n8043 , n8268 );
and ( n8728 , n8039 , n8268 );
or ( n8729 , n8726 , n8727 , n8728 );
xor ( n8730 , n8725 , n8729 );
and ( n8731 , n8269 , n8273 );
and ( n8732 , n8274 , n8277 );
or ( n8733 , n8731 , n8732 );
xor ( n8734 , n8730 , n8733 );
buf ( n8735 , n8734 );
buf ( n8736 , n8735 );
not ( n8737 , n8736 );
buf ( n8738 , n534 );
not ( n8739 , n8738 );
nor ( n8740 , n8737 , n8739 );
xor ( n8741 , n8484 , n8740 );
xor ( n8742 , n8289 , n8481 );
nor ( n8743 , n8281 , n8739 );
and ( n8744 , n8742 , n8743 );
xor ( n8745 , n8742 , n8743 );
xor ( n8746 , n8293 , n8479 );
nor ( n8747 , n7841 , n8739 );
and ( n8748 , n8746 , n8747 );
xor ( n8749 , n8746 , n8747 );
xor ( n8750 , n8297 , n8477 );
nor ( n8751 , n7413 , n8739 );
and ( n8752 , n8750 , n8751 );
xor ( n8753 , n8750 , n8751 );
xor ( n8754 , n8301 , n8475 );
nor ( n8755 , n6997 , n8739 );
and ( n8756 , n8754 , n8755 );
xor ( n8757 , n8754 , n8755 );
xor ( n8758 , n8305 , n8473 );
nor ( n8759 , n6596 , n8739 );
and ( n8760 , n8758 , n8759 );
xor ( n8761 , n8758 , n8759 );
xor ( n8762 , n8309 , n8471 );
nor ( n8763 , n6212 , n8739 );
and ( n8764 , n8762 , n8763 );
xor ( n8765 , n8762 , n8763 );
xor ( n8766 , n8313 , n8469 );
nor ( n8767 , n5838 , n8739 );
and ( n8768 , n8766 , n8767 );
xor ( n8769 , n8766 , n8767 );
xor ( n8770 , n8317 , n8467 );
nor ( n8771 , n5477 , n8739 );
and ( n8772 , n8770 , n8771 );
xor ( n8773 , n8770 , n8771 );
xor ( n8774 , n8321 , n8465 );
nor ( n8775 , n5126 , n8739 );
and ( n8776 , n8774 , n8775 );
xor ( n8777 , n8774 , n8775 );
xor ( n8778 , n8325 , n8463 );
nor ( n8779 , n4786 , n8739 );
and ( n8780 , n8778 , n8779 );
xor ( n8781 , n8778 , n8779 );
xor ( n8782 , n8329 , n8461 );
nor ( n8783 , n4458 , n8739 );
and ( n8784 , n8782 , n8783 );
xor ( n8785 , n8782 , n8783 );
xor ( n8786 , n8333 , n8459 );
nor ( n8787 , n4151 , n8739 );
and ( n8788 , n8786 , n8787 );
xor ( n8789 , n8786 , n8787 );
xor ( n8790 , n8337 , n8457 );
nor ( n8791 , n3853 , n8739 );
and ( n8792 , n8790 , n8791 );
xor ( n8793 , n8790 , n8791 );
xor ( n8794 , n8341 , n8455 );
nor ( n8795 , n3570 , n8739 );
and ( n8796 , n8794 , n8795 );
xor ( n8797 , n8794 , n8795 );
xor ( n8798 , n8345 , n8453 );
nor ( n8799 , n3300 , n8739 );
and ( n8800 , n8798 , n8799 );
xor ( n8801 , n8798 , n8799 );
xor ( n8802 , n8349 , n8451 );
nor ( n8803 , n3043 , n8739 );
and ( n8804 , n8802 , n8803 );
xor ( n8805 , n8802 , n8803 );
xor ( n8806 , n8353 , n8449 );
nor ( n8807 , n2797 , n8739 );
and ( n8808 , n8806 , n8807 );
xor ( n8809 , n8806 , n8807 );
xor ( n8810 , n8357 , n8447 );
nor ( n8811 , n2566 , n8739 );
and ( n8812 , n8810 , n8811 );
xor ( n8813 , n8810 , n8811 );
xor ( n8814 , n8361 , n8445 );
nor ( n8815 , n2343 , n8739 );
and ( n8816 , n8814 , n8815 );
xor ( n8817 , n8814 , n8815 );
xor ( n8818 , n8365 , n8443 );
nor ( n8819 , n2137 , n8739 );
and ( n8820 , n8818 , n8819 );
xor ( n8821 , n8818 , n8819 );
xor ( n8822 , n8369 , n8441 );
nor ( n8823 , n1945 , n8739 );
and ( n8824 , n8822 , n8823 );
xor ( n8825 , n8822 , n8823 );
xor ( n8826 , n8373 , n8439 );
nor ( n8827 , n1766 , n8739 );
and ( n8828 , n8826 , n8827 );
xor ( n8829 , n8826 , n8827 );
xor ( n8830 , n8377 , n8437 );
nor ( n8831 , n1598 , n8739 );
and ( n8832 , n8830 , n8831 );
xor ( n8833 , n8830 , n8831 );
xor ( n8834 , n8381 , n8435 );
nor ( n8835 , n1445 , n8739 );
and ( n8836 , n8834 , n8835 );
xor ( n8837 , n8834 , n8835 );
xor ( n8838 , n8385 , n8433 );
nor ( n8839 , n1303 , n8739 );
and ( n8840 , n8838 , n8839 );
xor ( n8841 , n8838 , n8839 );
xor ( n8842 , n8389 , n8431 );
nor ( n8843 , n1176 , n8739 );
and ( n8844 , n8842 , n8843 );
xor ( n8845 , n8842 , n8843 );
xor ( n8846 , n8393 , n8429 );
nor ( n8847 , n1062 , n8739 );
and ( n8848 , n8846 , n8847 );
xor ( n8849 , n8846 , n8847 );
xor ( n8850 , n8397 , n8427 );
nor ( n8851 , n958 , n8739 );
and ( n8852 , n8850 , n8851 );
xor ( n8853 , n8850 , n8851 );
xor ( n8854 , n8401 , n8425 );
nor ( n8855 , n868 , n8739 );
and ( n8856 , n8854 , n8855 );
xor ( n8857 , n8854 , n8855 );
xor ( n8858 , n8405 , n8423 );
nor ( n8859 , n796 , n8739 );
and ( n8860 , n8858 , n8859 );
xor ( n8861 , n8858 , n8859 );
xor ( n8862 , n8409 , n8421 );
nor ( n8863 , n733 , n8739 );
and ( n8864 , n8862 , n8863 );
xor ( n8865 , n8862 , n8863 );
xor ( n8866 , n8414 , n8419 );
nor ( n8867 , n684 , n8739 );
and ( n8868 , n8866 , n8867 );
xor ( n8869 , n8866 , n8867 );
xor ( n8870 , n8416 , n8417 );
buf ( n8871 , n8870 );
nor ( n8872 , n646 , n8739 );
and ( n8873 , n8871 , n8872 );
xor ( n8874 , n8871 , n8872 );
nor ( n8875 , n601 , n7843 );
buf ( n8876 , n8875 );
nor ( n8877 , n622 , n8739 );
and ( n8878 , n8876 , n8877 );
buf ( n8879 , n8878 );
and ( n8880 , n8874 , n8879 );
or ( n8881 , n8873 , n8880 );
and ( n8882 , n8869 , n8881 );
or ( n8883 , n8868 , n8882 );
and ( n8884 , n8865 , n8883 );
or ( n8885 , n8864 , n8884 );
and ( n8886 , n8861 , n8885 );
or ( n8887 , n8860 , n8886 );
and ( n8888 , n8857 , n8887 );
or ( n8889 , n8856 , n8888 );
and ( n8890 , n8853 , n8889 );
or ( n8891 , n8852 , n8890 );
and ( n8892 , n8849 , n8891 );
or ( n8893 , n8848 , n8892 );
and ( n8894 , n8845 , n8893 );
or ( n8895 , n8844 , n8894 );
and ( n8896 , n8841 , n8895 );
or ( n8897 , n8840 , n8896 );
and ( n8898 , n8837 , n8897 );
or ( n8899 , n8836 , n8898 );
and ( n8900 , n8833 , n8899 );
or ( n8901 , n8832 , n8900 );
and ( n8902 , n8829 , n8901 );
or ( n8903 , n8828 , n8902 );
and ( n8904 , n8825 , n8903 );
or ( n8905 , n8824 , n8904 );
and ( n8906 , n8821 , n8905 );
or ( n8907 , n8820 , n8906 );
and ( n8908 , n8817 , n8907 );
or ( n8909 , n8816 , n8908 );
and ( n8910 , n8813 , n8909 );
or ( n8911 , n8812 , n8910 );
and ( n8912 , n8809 , n8911 );
or ( n8913 , n8808 , n8912 );
and ( n8914 , n8805 , n8913 );
or ( n8915 , n8804 , n8914 );
and ( n8916 , n8801 , n8915 );
or ( n8917 , n8800 , n8916 );
and ( n8918 , n8797 , n8917 );
or ( n8919 , n8796 , n8918 );
and ( n8920 , n8793 , n8919 );
or ( n8921 , n8792 , n8920 );
and ( n8922 , n8789 , n8921 );
or ( n8923 , n8788 , n8922 );
and ( n8924 , n8785 , n8923 );
or ( n8925 , n8784 , n8924 );
and ( n8926 , n8781 , n8925 );
or ( n8927 , n8780 , n8926 );
and ( n8928 , n8777 , n8927 );
or ( n8929 , n8776 , n8928 );
and ( n8930 , n8773 , n8929 );
or ( n8931 , n8772 , n8930 );
and ( n8932 , n8769 , n8931 );
or ( n8933 , n8768 , n8932 );
and ( n8934 , n8765 , n8933 );
or ( n8935 , n8764 , n8934 );
and ( n8936 , n8761 , n8935 );
or ( n8937 , n8760 , n8936 );
and ( n8938 , n8757 , n8937 );
or ( n8939 , n8756 , n8938 );
and ( n8940 , n8753 , n8939 );
or ( n8941 , n8752 , n8940 );
and ( n8942 , n8749 , n8941 );
or ( n8943 , n8748 , n8942 );
and ( n8944 , n8745 , n8943 );
or ( n8945 , n8744 , n8944 );
xor ( n8946 , n8741 , n8945 );
buf ( n8947 , n8946 );
buf ( n8948 , n8947 );
not ( n8949 , n8948 );
buf ( n8950 , n535 );
not ( n8951 , n8950 );
and ( n8952 , n8951 , n8948 );
nor ( n8953 , n8949 , n8952 );
buf ( n8954 , n497 );
not ( n8955 , n8954 );
nor ( n8956 , n601 , n8955 );
buf ( n8957 , n8956 );
nor ( n8958 , n622 , n652 );
xor ( n8959 , n8957 , n8958 );
buf ( n8960 , n8959 );
nor ( n8961 , n646 , n624 );
xor ( n8962 , n8960 , n8961 );
and ( n8963 , n605 , n625 );
buf ( n8964 , n8963 );
xor ( n8965 , n8962 , n8964 );
nor ( n8966 , n684 , n648 );
xor ( n8967 , n8965 , n8966 );
and ( n8968 , n627 , n649 );
and ( n8969 , n650 , n657 );
or ( n8970 , n8968 , n8969 );
xor ( n8971 , n8967 , n8970 );
nor ( n8972 , n733 , n686 );
xor ( n8973 , n8971 , n8972 );
and ( n8974 , n658 , n687 );
and ( n8975 , n688 , n700 );
or ( n8976 , n8974 , n8975 );
xor ( n8977 , n8973 , n8976 );
nor ( n8978 , n796 , n735 );
xor ( n8979 , n8977 , n8978 );
and ( n8980 , n701 , n736 );
and ( n8981 , n737 , n755 );
or ( n8982 , n8980 , n8981 );
xor ( n8983 , n8979 , n8982 );
nor ( n8984 , n868 , n798 );
xor ( n8985 , n8983 , n8984 );
and ( n8986 , n756 , n799 );
and ( n8987 , n800 , n824 );
or ( n8988 , n8986 , n8987 );
xor ( n8989 , n8985 , n8988 );
nor ( n8990 , n958 , n870 );
xor ( n8991 , n8989 , n8990 );
and ( n8992 , n825 , n871 );
and ( n8993 , n872 , n902 );
or ( n8994 , n8992 , n8993 );
xor ( n8995 , n8991 , n8994 );
nor ( n8996 , n1062 , n960 );
xor ( n8997 , n8995 , n8996 );
and ( n8998 , n903 , n961 );
and ( n8999 , n962 , n998 );
or ( n9000 , n8998 , n8999 );
xor ( n9001 , n8997 , n9000 );
nor ( n9002 , n1176 , n1064 );
xor ( n9003 , n9001 , n9002 );
and ( n9004 , n999 , n1065 );
and ( n9005 , n1066 , n1108 );
or ( n9006 , n9004 , n9005 );
xor ( n9007 , n9003 , n9006 );
nor ( n9008 , n1303 , n1178 );
xor ( n9009 , n9007 , n9008 );
and ( n9010 , n1109 , n1179 );
and ( n9011 , n1180 , n1228 );
or ( n9012 , n9010 , n9011 );
xor ( n9013 , n9009 , n9012 );
nor ( n9014 , n1445 , n1305 );
xor ( n9015 , n9013 , n9014 );
and ( n9016 , n1229 , n1306 );
and ( n9017 , n1307 , n1361 );
or ( n9018 , n9016 , n9017 );
xor ( n9019 , n9015 , n9018 );
nor ( n9020 , n1598 , n1447 );
xor ( n9021 , n9019 , n9020 );
and ( n9022 , n1362 , n1448 );
and ( n9023 , n1449 , n1509 );
or ( n9024 , n9022 , n9023 );
xor ( n9025 , n9021 , n9024 );
nor ( n9026 , n1766 , n1600 );
xor ( n9027 , n9025 , n9026 );
and ( n9028 , n1510 , n1601 );
and ( n9029 , n1602 , n1668 );
or ( n9030 , n9028 , n9029 );
xor ( n9031 , n9027 , n9030 );
nor ( n9032 , n1945 , n1768 );
xor ( n9033 , n9031 , n9032 );
and ( n9034 , n1669 , n1769 );
and ( n9035 , n1770 , n1842 );
or ( n9036 , n9034 , n9035 );
xor ( n9037 , n9033 , n9036 );
nor ( n9038 , n2137 , n1947 );
xor ( n9039 , n9037 , n9038 );
and ( n9040 , n1843 , n1948 );
and ( n9041 , n1949 , n2027 );
or ( n9042 , n9040 , n9041 );
xor ( n9043 , n9039 , n9042 );
nor ( n9044 , n2343 , n2139 );
xor ( n9045 , n9043 , n9044 );
and ( n9046 , n2028 , n2140 );
and ( n9047 , n2141 , n2225 );
or ( n9048 , n9046 , n9047 );
xor ( n9049 , n9045 , n9048 );
nor ( n9050 , n2566 , n2345 );
xor ( n9051 , n9049 , n9050 );
and ( n9052 , n2226 , n2346 );
and ( n9053 , n2347 , n2437 );
or ( n9054 , n9052 , n9053 );
xor ( n9055 , n9051 , n9054 );
nor ( n9056 , n2797 , n2568 );
xor ( n9057 , n9055 , n9056 );
and ( n9058 , n2438 , n2569 );
and ( n9059 , n2570 , n2666 );
or ( n9060 , n9058 , n9059 );
xor ( n9061 , n9057 , n9060 );
nor ( n9062 , n3043 , n2799 );
xor ( n9063 , n9061 , n9062 );
and ( n9064 , n2667 , n2800 );
and ( n9065 , n2801 , n2903 );
or ( n9066 , n9064 , n9065 );
xor ( n9067 , n9063 , n9066 );
nor ( n9068 , n3300 , n3045 );
xor ( n9069 , n9067 , n9068 );
and ( n9070 , n2904 , n3046 );
and ( n9071 , n3047 , n3155 );
or ( n9072 , n9070 , n9071 );
xor ( n9073 , n9069 , n9072 );
nor ( n9074 , n3570 , n3302 );
xor ( n9075 , n9073 , n9074 );
and ( n9076 , n3156 , n3303 );
and ( n9077 , n3304 , n3418 );
or ( n9078 , n9076 , n9077 );
xor ( n9079 , n9075 , n9078 );
nor ( n9080 , n3853 , n3572 );
xor ( n9081 , n9079 , n9080 );
and ( n9082 , n3419 , n3573 );
and ( n9083 , n3574 , n3694 );
or ( n9084 , n9082 , n9083 );
xor ( n9085 , n9081 , n9084 );
nor ( n9086 , n4151 , n3855 );
xor ( n9087 , n9085 , n9086 );
and ( n9088 , n3695 , n3856 );
and ( n9089 , n3857 , n3983 );
or ( n9090 , n9088 , n9089 );
xor ( n9091 , n9087 , n9090 );
nor ( n9092 , n4458 , n4153 );
xor ( n9093 , n9091 , n9092 );
and ( n9094 , n3984 , n4154 );
and ( n9095 , n4155 , n4287 );
or ( n9096 , n9094 , n9095 );
xor ( n9097 , n9093 , n9096 );
nor ( n9098 , n4786 , n4460 );
xor ( n9099 , n9097 , n9098 );
and ( n9100 , n4288 , n4461 );
and ( n9101 , n4462 , n4600 );
or ( n9102 , n9100 , n9101 );
xor ( n9103 , n9099 , n9102 );
nor ( n9104 , n5126 , n4788 );
xor ( n9105 , n9103 , n9104 );
and ( n9106 , n4601 , n4789 );
and ( n9107 , n4790 , n4934 );
or ( n9108 , n9106 , n9107 );
xor ( n9109 , n9105 , n9108 );
nor ( n9110 , n5477 , n5128 );
xor ( n9111 , n9109 , n9110 );
and ( n9112 , n4935 , n5129 );
and ( n9113 , n5130 , n5280 );
or ( n9114 , n9112 , n9113 );
xor ( n9115 , n9111 , n9114 );
nor ( n9116 , n5838 , n5479 );
xor ( n9117 , n9115 , n9116 );
and ( n9118 , n5281 , n5480 );
and ( n9119 , n5481 , n5637 );
or ( n9120 , n9118 , n9119 );
xor ( n9121 , n9117 , n9120 );
nor ( n9122 , n6212 , n5840 );
xor ( n9123 , n9121 , n9122 );
and ( n9124 , n5638 , n5841 );
and ( n9125 , n5842 , n6004 );
or ( n9126 , n9124 , n9125 );
xor ( n9127 , n9123 , n9126 );
nor ( n9128 , n6596 , n6214 );
xor ( n9129 , n9127 , n9128 );
and ( n9130 , n6005 , n6215 );
and ( n9131 , n6216 , n6384 );
or ( n9132 , n9130 , n9131 );
xor ( n9133 , n9129 , n9132 );
nor ( n9134 , n6997 , n6598 );
xor ( n9135 , n9133 , n9134 );
and ( n9136 , n6385 , n6599 );
and ( n9137 , n6600 , n6774 );
or ( n9138 , n9136 , n9137 );
xor ( n9139 , n9135 , n9138 );
nor ( n9140 , n7413 , n6999 );
xor ( n9141 , n9139 , n9140 );
and ( n9142 , n6775 , n7000 );
and ( n9143 , n7001 , n7181 );
or ( n9144 , n9142 , n9143 );
xor ( n9145 , n9141 , n9144 );
nor ( n9146 , n7841 , n7415 );
xor ( n9147 , n9145 , n9146 );
and ( n9148 , n7182 , n7416 );
and ( n9149 , n7417 , n7603 );
or ( n9150 , n9148 , n9149 );
xor ( n9151 , n9147 , n9150 );
nor ( n9152 , n8281 , n7843 );
xor ( n9153 , n9151 , n9152 );
and ( n9154 , n7604 , n7844 );
and ( n9155 , n7845 , n8037 );
or ( n9156 , n9154 , n9155 );
xor ( n9157 , n9153 , n9156 );
nor ( n9158 , n8737 , n8283 );
xor ( n9159 , n9157 , n9158 );
and ( n9160 , n8038 , n8284 );
and ( n9161 , n8285 , n8483 );
or ( n9162 , n9160 , n9161 );
xor ( n9163 , n9159 , n9162 );
and ( n9164 , n8706 , n8707 );
and ( n9165 , n8707 , n8722 );
and ( n9166 , n8706 , n8722 );
or ( n9167 , n9164 , n9165 , n9166 );
and ( n9168 , n8494 , n8701 );
and ( n9169 , n8701 , n8723 );
and ( n9170 , n8494 , n8723 );
or ( n9171 , n9168 , n9169 , n9170 );
xor ( n9172 , n9167 , n9171 );
and ( n9173 , n8498 , n8576 );
and ( n9174 , n8576 , n8700 );
and ( n9175 , n8498 , n8700 );
or ( n9176 , n9173 , n9174 , n9175 );
and ( n9177 , n8581 , n8628 );
and ( n9178 , n8628 , n8699 );
and ( n9179 , n8581 , n8699 );
or ( n9180 , n9177 , n9178 , n9179 );
and ( n9181 , n8511 , n8548 );
and ( n9182 , n8548 , n8574 );
and ( n9183 , n8511 , n8574 );
or ( n9184 , n9181 , n9182 , n9183 );
and ( n9185 , n8585 , n8589 );
and ( n9186 , n8589 , n8627 );
and ( n9187 , n8585 , n8627 );
or ( n9188 , n9185 , n9186 , n9187 );
xor ( n9189 , n9184 , n9188 );
and ( n9190 , n8553 , n8557 );
and ( n9191 , n8557 , n8573 );
and ( n9192 , n8553 , n8573 );
or ( n9193 , n9190 , n9191 , n9192 );
and ( n9194 , n8535 , n8540 );
and ( n9195 , n8540 , n8546 );
and ( n9196 , n8535 , n8546 );
or ( n9197 , n9194 , n9195 , n9196 );
and ( n9198 , n8525 , n8526 );
and ( n9199 , n8526 , n8528 );
and ( n9200 , n8525 , n8528 );
or ( n9201 , n9198 , n9199 , n9200 );
and ( n9202 , n8536 , n8537 );
and ( n9203 , n8537 , n8539 );
and ( n9204 , n8536 , n8539 );
or ( n9205 , n9202 , n9203 , n9204 );
xor ( n9206 , n9201 , n9205 );
and ( n9207 , n7385 , n663 );
and ( n9208 , n7808 , n635 );
xor ( n9209 , n9207 , n9208 );
and ( n9210 , n8079 , n606 );
xor ( n9211 , n9209 , n9210 );
xor ( n9212 , n9206 , n9211 );
xor ( n9213 , n9197 , n9212 );
and ( n9214 , n8542 , n8543 );
and ( n9215 , n8543 , n8545 );
and ( n9216 , n8542 , n8545 );
or ( n9217 , n9214 , n9215 , n9216 );
and ( n9218 , n6187 , n840 );
and ( n9219 , n6569 , n771 );
xor ( n9220 , n9218 , n9219 );
and ( n9221 , n6816 , n719 );
xor ( n9222 , n9220 , n9221 );
xor ( n9223 , n9217 , n9222 );
and ( n9224 , n4959 , n1134 );
and ( n9225 , n5459 , n1034 );
xor ( n9226 , n9224 , n9225 );
and ( n9227 , n5819 , n940 );
xor ( n9228 , n9226 , n9227 );
xor ( n9229 , n9223 , n9228 );
xor ( n9230 , n9213 , n9229 );
xor ( n9231 , n9193 , n9230 );
and ( n9232 , n8562 , n8566 );
and ( n9233 , n8566 , n8572 );
and ( n9234 , n8562 , n8572 );
or ( n9235 , n9232 , n9233 , n9234 );
and ( n9236 , n8598 , n8603 );
and ( n9237 , n8603 , n8609 );
and ( n9238 , n8598 , n8609 );
or ( n9239 , n9236 , n9237 , n9238 );
xor ( n9240 , n9235 , n9239 );
and ( n9241 , n8568 , n8569 );
and ( n9242 , n8569 , n8571 );
and ( n9243 , n8568 , n8571 );
or ( n9244 , n9241 , n9242 , n9243 );
and ( n9245 , n8599 , n8600 );
and ( n9246 , n8600 , n8602 );
and ( n9247 , n8599 , n8602 );
or ( n9248 , n9245 , n9246 , n9247 );
xor ( n9249 , n9244 , n9248 );
and ( n9250 , n4132 , n1551 );
and ( n9251 , n4438 , n1424 );
xor ( n9252 , n9250 , n9251 );
and ( n9253 , n4766 , n1254 );
xor ( n9254 , n9252 , n9253 );
xor ( n9255 , n9249 , n9254 );
xor ( n9256 , n9240 , n9255 );
xor ( n9257 , n9231 , n9256 );
xor ( n9258 , n9189 , n9257 );
xor ( n9259 , n9180 , n9258 );
and ( n9260 , n8633 , n8659 );
and ( n9261 , n8659 , n8698 );
and ( n9262 , n8633 , n8698 );
or ( n9263 , n9260 , n9261 , n9262 );
and ( n9264 , n8637 , n8641 );
and ( n9265 , n8641 , n8658 );
and ( n9266 , n8637 , n8658 );
or ( n9267 , n9264 , n9265 , n9266 );
and ( n9268 , n8594 , n8610 );
and ( n9269 , n8610 , n8626 );
and ( n9270 , n8594 , n8626 );
or ( n9271 , n9268 , n9269 , n9270 );
xor ( n9272 , n9267 , n9271 );
and ( n9273 , n8615 , n8619 );
and ( n9274 , n8619 , n8625 );
and ( n9275 , n8615 , n8625 );
or ( n9276 , n9273 , n9274 , n9275 );
and ( n9277 , n8647 , n8648 );
and ( n9278 , n8648 , n8650 );
and ( n9279 , n8647 , n8650 );
or ( n9280 , n9277 , n9278 , n9279 );
and ( n9281 , n8621 , n8622 );
and ( n9282 , n8622 , n8624 );
and ( n9283 , n8621 , n8624 );
or ( n9284 , n9281 , n9282 , n9283 );
xor ( n9285 , n9280 , n9284 );
and ( n9286 , n1933 , n3495 );
and ( n9287 , n2120 , n3271 );
xor ( n9288 , n9286 , n9287 );
and ( n9289 , n2324 , n2981 );
xor ( n9290 , n9288 , n9289 );
xor ( n9291 , n9285 , n9290 );
xor ( n9292 , n9276 , n9291 );
and ( n9293 , n8605 , n8606 );
and ( n9294 , n8606 , n8608 );
and ( n9295 , n8605 , n8608 );
or ( n9296 , n9293 , n9294 , n9295 );
and ( n9297 , n3182 , n2100 );
and ( n9298 , n3545 , n1882 );
xor ( n9299 , n9297 , n9298 );
and ( n9300 , n3801 , n1738 );
xor ( n9301 , n9299 , n9300 );
xor ( n9302 , n9296 , n9301 );
and ( n9303 , n3024 , n2298 );
buf ( n9304 , n9303 );
xor ( n9305 , n9302 , n9304 );
xor ( n9306 , n9292 , n9305 );
xor ( n9307 , n9272 , n9306 );
xor ( n9308 , n9263 , n9307 );
and ( n9309 , n8664 , n8681 );
and ( n9310 , n8681 , n8697 );
and ( n9311 , n8664 , n8697 );
or ( n9312 , n9309 , n9310 , n9311 );
and ( n9313 , n8646 , n8651 );
and ( n9314 , n8651 , n8657 );
and ( n9315 , n8646 , n8657 );
or ( n9316 , n9313 , n9314 , n9315 );
and ( n9317 , n8686 , n8690 );
and ( n9318 , n8690 , n8696 );
and ( n9319 , n8686 , n8696 );
or ( n9320 , n9317 , n9318 , n9319 );
xor ( n9321 , n9316 , n9320 );
and ( n9322 , n8653 , n8654 );
and ( n9323 , n8654 , n8656 );
and ( n9324 , n8653 , n8656 );
or ( n9325 , n9322 , n9323 , n9324 );
and ( n9326 , n1383 , n4403 );
and ( n9327 , n1580 , n4102 );
xor ( n9328 , n9326 , n9327 );
and ( n9329 , n1694 , n3749 );
xor ( n9330 , n9328 , n9329 );
xor ( n9331 , n9325 , n9330 );
and ( n9332 , n1047 , n5408 );
and ( n9333 , n1164 , n5103 );
xor ( n9334 , n9332 , n9333 );
and ( n9335 , n1287 , n4730 );
xor ( n9336 , n9334 , n9335 );
xor ( n9337 , n9331 , n9336 );
xor ( n9338 , n9321 , n9337 );
xor ( n9339 , n9312 , n9338 );
and ( n9340 , n8668 , n8674 );
and ( n9341 , n8674 , n8680 );
and ( n9342 , n8668 , n8680 );
or ( n9343 , n9340 , n9341 , n9342 );
and ( n9344 , n8670 , n8671 );
and ( n9345 , n8671 , n8673 );
and ( n9346 , n8670 , n8673 );
or ( n9347 , n9344 , n9345 , n9346 );
buf ( n9348 , n433 );
and ( n9349 , n599 , n9348 );
and ( n9350 , n608 , n8669 );
xor ( n9351 , n9349 , n9350 );
and ( n9352 , n611 , n8243 );
xor ( n9353 , n9351 , n9352 );
xor ( n9354 , n9347 , n9353 );
and ( n9355 , n632 , n7662 );
and ( n9356 , n671 , n7310 );
xor ( n9357 , n9355 , n9356 );
and ( n9358 , n715 , n6971 );
xor ( n9359 , n9357 , n9358 );
xor ( n9360 , n9354 , n9359 );
xor ( n9361 , n9343 , n9360 );
and ( n9362 , n8692 , n8693 );
and ( n9363 , n8693 , n8695 );
and ( n9364 , n8692 , n8695 );
or ( n9365 , n9362 , n9363 , n9364 );
and ( n9366 , n8676 , n8677 );
and ( n9367 , n8677 , n8679 );
and ( n9368 , n8676 , n8679 );
or ( n9369 , n9366 , n9367 , n9368 );
xor ( n9370 , n9365 , n9369 );
and ( n9371 , n783 , n6504 );
and ( n9372 , n856 , n6132 );
xor ( n9373 , n9371 , n9372 );
and ( n9374 , n925 , n5765 );
xor ( n9375 , n9373 , n9374 );
xor ( n9376 , n9370 , n9375 );
xor ( n9377 , n9361 , n9376 );
xor ( n9378 , n9339 , n9377 );
xor ( n9379 , n9308 , n9378 );
xor ( n9380 , n9259 , n9379 );
xor ( n9381 , n9176 , n9380 );
and ( n9382 , n8502 , n8506 );
and ( n9383 , n8506 , n8575 );
and ( n9384 , n8502 , n8575 );
or ( n9385 , n9382 , n9383 , n9384 );
and ( n9386 , n8709 , n8721 );
xor ( n9387 , n9385 , n9386 );
and ( n9388 , n8713 , n8720 );
and ( n9389 , n8515 , n8530 );
and ( n9390 , n8530 , n8547 );
and ( n9391 , n8515 , n8547 );
or ( n9392 , n9389 , n9390 , n9391 );
and ( n9393 , n8717 , n8719 );
xor ( n9394 , n9392 , n9393 );
and ( n9395 , n8519 , n8523 );
and ( n9396 , n8523 , n8529 );
and ( n9397 , n8519 , n8529 );
or ( n9398 , n9395 , n9396 , n9397 );
and ( n9399 , n8718 , n615 );
buf ( n9400 , n433 );
and ( n9401 , n9400 , n612 );
xor ( n9402 , n9399 , n9401 );
xor ( n9403 , n9398 , n9402 );
xor ( n9404 , n9394 , n9403 );
xor ( n9405 , n9388 , n9404 );
xor ( n9406 , n9387 , n9405 );
xor ( n9407 , n9381 , n9406 );
xor ( n9408 , n9172 , n9407 );
and ( n9409 , n8485 , n8489 );
and ( n9410 , n8489 , n8724 );
and ( n9411 , n8485 , n8724 );
or ( n9412 , n9409 , n9410 , n9411 );
xor ( n9413 , n9408 , n9412 );
and ( n9414 , n8725 , n8729 );
and ( n9415 , n8730 , n8733 );
or ( n9416 , n9414 , n9415 );
xor ( n9417 , n9413 , n9416 );
buf ( n9418 , n9417 );
buf ( n9419 , n9418 );
not ( n9420 , n9419 );
nor ( n9421 , n9420 , n8739 );
xor ( n9422 , n9163 , n9421 );
and ( n9423 , n8484 , n8740 );
and ( n9424 , n8741 , n8945 );
or ( n9425 , n9423 , n9424 );
xor ( n9426 , n9422 , n9425 );
buf ( n9427 , n9426 );
buf ( n9428 , n9427 );
not ( n9429 , n9428 );
buf ( n9430 , n536 );
not ( n9431 , n9430 );
nor ( n9432 , n9429 , n9431 );
xor ( n9433 , n8953 , n9432 );
xor ( n9434 , n8745 , n8943 );
buf ( n9435 , n9434 );
buf ( n9436 , n9435 );
not ( n9437 , n9436 );
and ( n9438 , n8951 , n9436 );
nor ( n9439 , n9437 , n9438 );
nor ( n9440 , n8949 , n9431 );
and ( n9441 , n9439 , n9440 );
xor ( n9442 , n9439 , n9440 );
xor ( n9443 , n8749 , n8941 );
buf ( n9444 , n9443 );
buf ( n9445 , n9444 );
not ( n9446 , n9445 );
and ( n9447 , n8951 , n9445 );
nor ( n9448 , n9446 , n9447 );
nor ( n9449 , n9437 , n9431 );
and ( n9450 , n9448 , n9449 );
xor ( n9451 , n9448 , n9449 );
xor ( n9452 , n8753 , n8939 );
buf ( n9453 , n9452 );
buf ( n9454 , n9453 );
not ( n9455 , n9454 );
and ( n9456 , n8951 , n9454 );
nor ( n9457 , n9455 , n9456 );
nor ( n9458 , n9446 , n9431 );
and ( n9459 , n9457 , n9458 );
xor ( n9460 , n9457 , n9458 );
xor ( n9461 , n8757 , n8937 );
buf ( n9462 , n9461 );
buf ( n9463 , n9462 );
not ( n9464 , n9463 );
and ( n9465 , n8951 , n9463 );
nor ( n9466 , n9464 , n9465 );
nor ( n9467 , n9455 , n9431 );
and ( n9468 , n9466 , n9467 );
xor ( n9469 , n9466 , n9467 );
xor ( n9470 , n8761 , n8935 );
buf ( n9471 , n9470 );
buf ( n9472 , n9471 );
not ( n9473 , n9472 );
and ( n9474 , n8951 , n9472 );
nor ( n9475 , n9473 , n9474 );
nor ( n9476 , n9464 , n9431 );
and ( n9477 , n9475 , n9476 );
xor ( n9478 , n9475 , n9476 );
xor ( n9479 , n8765 , n8933 );
buf ( n9480 , n9479 );
buf ( n9481 , n9480 );
not ( n9482 , n9481 );
and ( n9483 , n8951 , n9481 );
nor ( n9484 , n9482 , n9483 );
nor ( n9485 , n9473 , n9431 );
and ( n9486 , n9484 , n9485 );
xor ( n9487 , n9484 , n9485 );
xor ( n9488 , n8769 , n8931 );
buf ( n9489 , n9488 );
buf ( n9490 , n9489 );
not ( n9491 , n9490 );
and ( n9492 , n8951 , n9490 );
nor ( n9493 , n9491 , n9492 );
nor ( n9494 , n9482 , n9431 );
and ( n9495 , n9493 , n9494 );
xor ( n9496 , n9493 , n9494 );
xor ( n9497 , n8773 , n8929 );
buf ( n9498 , n9497 );
buf ( n9499 , n9498 );
not ( n9500 , n9499 );
and ( n9501 , n8951 , n9499 );
nor ( n9502 , n9500 , n9501 );
nor ( n9503 , n9491 , n9431 );
and ( n9504 , n9502 , n9503 );
xor ( n9505 , n9502 , n9503 );
xor ( n9506 , n8777 , n8927 );
buf ( n9507 , n9506 );
buf ( n9508 , n9507 );
not ( n9509 , n9508 );
and ( n9510 , n8951 , n9508 );
nor ( n9511 , n9509 , n9510 );
nor ( n9512 , n9500 , n9431 );
and ( n9513 , n9511 , n9512 );
xor ( n9514 , n9511 , n9512 );
xor ( n9515 , n8781 , n8925 );
buf ( n9516 , n9515 );
buf ( n9517 , n9516 );
not ( n9518 , n9517 );
and ( n9519 , n8951 , n9517 );
nor ( n9520 , n9518 , n9519 );
nor ( n9521 , n9509 , n9431 );
and ( n9522 , n9520 , n9521 );
xor ( n9523 , n9520 , n9521 );
xor ( n9524 , n8785 , n8923 );
buf ( n9525 , n9524 );
buf ( n9526 , n9525 );
not ( n9527 , n9526 );
and ( n9528 , n8951 , n9526 );
nor ( n9529 , n9527 , n9528 );
nor ( n9530 , n9518 , n9431 );
and ( n9531 , n9529 , n9530 );
xor ( n9532 , n9529 , n9530 );
xor ( n9533 , n8789 , n8921 );
buf ( n9534 , n9533 );
buf ( n9535 , n9534 );
not ( n9536 , n9535 );
and ( n9537 , n8951 , n9535 );
nor ( n9538 , n9536 , n9537 );
nor ( n9539 , n9527 , n9431 );
and ( n9540 , n9538 , n9539 );
xor ( n9541 , n9538 , n9539 );
xor ( n9542 , n8793 , n8919 );
buf ( n9543 , n9542 );
buf ( n9544 , n9543 );
not ( n9545 , n9544 );
and ( n9546 , n8951 , n9544 );
nor ( n9547 , n9545 , n9546 );
nor ( n9548 , n9536 , n9431 );
and ( n9549 , n9547 , n9548 );
xor ( n9550 , n9547 , n9548 );
xor ( n9551 , n8797 , n8917 );
buf ( n9552 , n9551 );
buf ( n9553 , n9552 );
not ( n9554 , n9553 );
and ( n9555 , n8951 , n9553 );
nor ( n9556 , n9554 , n9555 );
nor ( n9557 , n9545 , n9431 );
and ( n9558 , n9556 , n9557 );
xor ( n9559 , n9556 , n9557 );
xor ( n9560 , n8801 , n8915 );
buf ( n9561 , n9560 );
buf ( n9562 , n9561 );
not ( n9563 , n9562 );
and ( n9564 , n8951 , n9562 );
nor ( n9565 , n9563 , n9564 );
nor ( n9566 , n9554 , n9431 );
and ( n9567 , n9565 , n9566 );
xor ( n9568 , n9565 , n9566 );
xor ( n9569 , n8805 , n8913 );
buf ( n9570 , n9569 );
buf ( n9571 , n9570 );
not ( n9572 , n9571 );
and ( n9573 , n8951 , n9571 );
nor ( n9574 , n9572 , n9573 );
nor ( n9575 , n9563 , n9431 );
and ( n9576 , n9574 , n9575 );
xor ( n9577 , n9574 , n9575 );
xor ( n9578 , n8809 , n8911 );
buf ( n9579 , n9578 );
buf ( n9580 , n9579 );
not ( n9581 , n9580 );
and ( n9582 , n8951 , n9580 );
nor ( n9583 , n9581 , n9582 );
nor ( n9584 , n9572 , n9431 );
and ( n9585 , n9583 , n9584 );
xor ( n9586 , n9583 , n9584 );
xor ( n9587 , n8813 , n8909 );
buf ( n9588 , n9587 );
buf ( n9589 , n9588 );
not ( n9590 , n9589 );
and ( n9591 , n8951 , n9589 );
nor ( n9592 , n9590 , n9591 );
nor ( n9593 , n9581 , n9431 );
and ( n9594 , n9592 , n9593 );
xor ( n9595 , n9592 , n9593 );
xor ( n9596 , n8817 , n8907 );
buf ( n9597 , n9596 );
buf ( n9598 , n9597 );
not ( n9599 , n9598 );
and ( n9600 , n8951 , n9598 );
nor ( n9601 , n9599 , n9600 );
nor ( n9602 , n9590 , n9431 );
and ( n9603 , n9601 , n9602 );
xor ( n9604 , n9601 , n9602 );
xor ( n9605 , n8821 , n8905 );
buf ( n9606 , n9605 );
buf ( n9607 , n9606 );
not ( n9608 , n9607 );
and ( n9609 , n8951 , n9607 );
nor ( n9610 , n9608 , n9609 );
nor ( n9611 , n9599 , n9431 );
and ( n9612 , n9610 , n9611 );
xor ( n9613 , n9610 , n9611 );
xor ( n9614 , n8825 , n8903 );
buf ( n9615 , n9614 );
buf ( n9616 , n9615 );
not ( n9617 , n9616 );
and ( n9618 , n8951 , n9616 );
nor ( n9619 , n9617 , n9618 );
nor ( n9620 , n9608 , n9431 );
and ( n9621 , n9619 , n9620 );
xor ( n9622 , n9619 , n9620 );
xor ( n9623 , n8829 , n8901 );
buf ( n9624 , n9623 );
buf ( n9625 , n9624 );
not ( n9626 , n9625 );
and ( n9627 , n8951 , n9625 );
nor ( n9628 , n9626 , n9627 );
nor ( n9629 , n9617 , n9431 );
and ( n9630 , n9628 , n9629 );
xor ( n9631 , n9628 , n9629 );
xor ( n9632 , n8833 , n8899 );
buf ( n9633 , n9632 );
buf ( n9634 , n9633 );
not ( n9635 , n9634 );
and ( n9636 , n8951 , n9634 );
nor ( n9637 , n9635 , n9636 );
nor ( n9638 , n9626 , n9431 );
and ( n9639 , n9637 , n9638 );
xor ( n9640 , n9637 , n9638 );
xor ( n9641 , n8837 , n8897 );
buf ( n9642 , n9641 );
buf ( n9643 , n9642 );
not ( n9644 , n9643 );
and ( n9645 , n8951 , n9643 );
nor ( n9646 , n9644 , n9645 );
nor ( n9647 , n9635 , n9431 );
and ( n9648 , n9646 , n9647 );
xor ( n9649 , n9646 , n9647 );
xor ( n9650 , n8841 , n8895 );
buf ( n9651 , n9650 );
buf ( n9652 , n9651 );
not ( n9653 , n9652 );
and ( n9654 , n8951 , n9652 );
nor ( n9655 , n9653 , n9654 );
nor ( n9656 , n9644 , n9431 );
and ( n9657 , n9655 , n9656 );
xor ( n9658 , n9655 , n9656 );
xor ( n9659 , n8845 , n8893 );
buf ( n9660 , n9659 );
buf ( n9661 , n9660 );
not ( n9662 , n9661 );
and ( n9663 , n8951 , n9661 );
nor ( n9664 , n9662 , n9663 );
nor ( n9665 , n9653 , n9431 );
and ( n9666 , n9664 , n9665 );
xor ( n9667 , n9664 , n9665 );
xor ( n9668 , n8849 , n8891 );
buf ( n9669 , n9668 );
buf ( n9670 , n9669 );
not ( n9671 , n9670 );
and ( n9672 , n8951 , n9670 );
nor ( n9673 , n9671 , n9672 );
nor ( n9674 , n9662 , n9431 );
and ( n9675 , n9673 , n9674 );
xor ( n9676 , n9673 , n9674 );
xor ( n9677 , n8853 , n8889 );
buf ( n9678 , n9677 );
buf ( n9679 , n9678 );
not ( n9680 , n9679 );
and ( n9681 , n8951 , n9679 );
nor ( n9682 , n9680 , n9681 );
nor ( n9683 , n9671 , n9431 );
and ( n9684 , n9682 , n9683 );
xor ( n9685 , n9682 , n9683 );
xor ( n9686 , n8857 , n8887 );
buf ( n9687 , n9686 );
buf ( n9688 , n9687 );
not ( n9689 , n9688 );
and ( n9690 , n8951 , n9688 );
nor ( n9691 , n9689 , n9690 );
nor ( n9692 , n9680 , n9431 );
and ( n9693 , n9691 , n9692 );
xor ( n9694 , n9691 , n9692 );
xor ( n9695 , n8861 , n8885 );
buf ( n9696 , n9695 );
buf ( n9697 , n9696 );
not ( n9698 , n9697 );
and ( n9699 , n8951 , n9697 );
nor ( n9700 , n9698 , n9699 );
nor ( n9701 , n9689 , n9431 );
and ( n9702 , n9700 , n9701 );
xor ( n9703 , n9700 , n9701 );
xor ( n9704 , n8865 , n8883 );
buf ( n9705 , n9704 );
buf ( n9706 , n9705 );
not ( n9707 , n9706 );
and ( n9708 , n8951 , n9706 );
nor ( n9709 , n9707 , n9708 );
nor ( n9710 , n9698 , n9431 );
and ( n9711 , n9709 , n9710 );
xor ( n9712 , n9709 , n9710 );
xor ( n9713 , n8869 , n8881 );
buf ( n9714 , n9713 );
buf ( n9715 , n9714 );
not ( n9716 , n9715 );
and ( n9717 , n8951 , n9715 );
nor ( n9718 , n9716 , n9717 );
nor ( n9719 , n9707 , n9431 );
and ( n9720 , n9718 , n9719 );
xor ( n9721 , n9718 , n9719 );
xor ( n9722 , n8874 , n8879 );
buf ( n9723 , n9722 );
buf ( n9724 , n9723 );
not ( n9725 , n9724 );
and ( n9726 , n8951 , n9724 );
nor ( n9727 , n9725 , n9726 );
nor ( n9728 , n9716 , n9431 );
and ( n9729 , n9727 , n9728 );
xor ( n9730 , n9727 , n9728 );
xor ( n9731 , n8876 , n8877 );
buf ( n9732 , n9731 );
buf ( n9733 , n9732 );
not ( n9734 , n9733 );
and ( n9735 , n8951 , n9733 );
nor ( n9736 , n9734 , n9735 );
nor ( n9737 , n9725 , n9431 );
and ( n9738 , n9736 , n9737 );
xor ( n9739 , n9736 , n9737 );
nor ( n9740 , n601 , n8283 );
buf ( n9741 , n9740 );
buf ( n9742 , n9741 );
not ( n9743 , n9742 );
and ( n9744 , n8951 , n9742 );
nor ( n9745 , n9743 , n9744 );
nor ( n9746 , n9734 , n9431 );
and ( n9747 , n9745 , n9746 );
xor ( n9748 , n9745 , n9746 );
nor ( n9749 , n601 , n8739 );
buf ( n9750 , n9749 );
buf ( n9751 , n9750 );
not ( n9752 , n9751 );
and ( n9753 , n8951 , n9751 );
nor ( n9754 , n9752 , n9753 );
nor ( n9755 , n9743 , n9431 );
and ( n9756 , n9754 , n9755 );
and ( n9757 , n9748 , n9756 );
or ( n9758 , n9747 , n9757 );
and ( n9759 , n9739 , n9758 );
or ( n9760 , n9738 , n9759 );
and ( n9761 , n9730 , n9760 );
or ( n9762 , n9729 , n9761 );
and ( n9763 , n9721 , n9762 );
or ( n9764 , n9720 , n9763 );
and ( n9765 , n9712 , n9764 );
or ( n9766 , n9711 , n9765 );
and ( n9767 , n9703 , n9766 );
or ( n9768 , n9702 , n9767 );
and ( n9769 , n9694 , n9768 );
or ( n9770 , n9693 , n9769 );
and ( n9771 , n9685 , n9770 );
or ( n9772 , n9684 , n9771 );
and ( n9773 , n9676 , n9772 );
or ( n9774 , n9675 , n9773 );
and ( n9775 , n9667 , n9774 );
or ( n9776 , n9666 , n9775 );
and ( n9777 , n9658 , n9776 );
or ( n9778 , n9657 , n9777 );
and ( n9779 , n9649 , n9778 );
or ( n9780 , n9648 , n9779 );
and ( n9781 , n9640 , n9780 );
or ( n9782 , n9639 , n9781 );
and ( n9783 , n9631 , n9782 );
or ( n9784 , n9630 , n9783 );
and ( n9785 , n9622 , n9784 );
or ( n9786 , n9621 , n9785 );
and ( n9787 , n9613 , n9786 );
or ( n9788 , n9612 , n9787 );
and ( n9789 , n9604 , n9788 );
or ( n9790 , n9603 , n9789 );
and ( n9791 , n9595 , n9790 );
or ( n9792 , n9594 , n9791 );
and ( n9793 , n9586 , n9792 );
or ( n9794 , n9585 , n9793 );
and ( n9795 , n9577 , n9794 );
or ( n9796 , n9576 , n9795 );
and ( n9797 , n9568 , n9796 );
or ( n9798 , n9567 , n9797 );
and ( n9799 , n9559 , n9798 );
or ( n9800 , n9558 , n9799 );
and ( n9801 , n9550 , n9800 );
or ( n9802 , n9549 , n9801 );
and ( n9803 , n9541 , n9802 );
or ( n9804 , n9540 , n9803 );
and ( n9805 , n9532 , n9804 );
or ( n9806 , n9531 , n9805 );
and ( n9807 , n9523 , n9806 );
or ( n9808 , n9522 , n9807 );
and ( n9809 , n9514 , n9808 );
or ( n9810 , n9513 , n9809 );
and ( n9811 , n9505 , n9810 );
or ( n9812 , n9504 , n9811 );
and ( n9813 , n9496 , n9812 );
or ( n9814 , n9495 , n9813 );
and ( n9815 , n9487 , n9814 );
or ( n9816 , n9486 , n9815 );
and ( n9817 , n9478 , n9816 );
or ( n9818 , n9477 , n9817 );
and ( n9819 , n9469 , n9818 );
or ( n9820 , n9468 , n9819 );
and ( n9821 , n9460 , n9820 );
or ( n9822 , n9459 , n9821 );
and ( n9823 , n9451 , n9822 );
or ( n9824 , n9450 , n9823 );
and ( n9825 , n9442 , n9824 );
or ( n9826 , n9441 , n9825 );
xor ( n9827 , n9433 , n9826 );
buf ( n9828 , n496 );
not ( n9829 , n9828 );
nor ( n9830 , n601 , n9829 );
buf ( n9831 , n9830 );
nor ( n9832 , n622 , n603 );
xor ( n9833 , n9831 , n9832 );
buf ( n9834 , n9833 );
nor ( n9835 , n646 , n652 );
xor ( n9836 , n9834 , n9835 );
and ( n9837 , n8957 , n8958 );
buf ( n9838 , n9837 );
xor ( n9839 , n9836 , n9838 );
nor ( n9840 , n684 , n624 );
xor ( n9841 , n9839 , n9840 );
and ( n9842 , n8960 , n8961 );
and ( n9843 , n8962 , n8964 );
or ( n9844 , n9842 , n9843 );
xor ( n9845 , n9841 , n9844 );
nor ( n9846 , n733 , n648 );
xor ( n9847 , n9845 , n9846 );
and ( n9848 , n8965 , n8966 );
and ( n9849 , n8967 , n8970 );
or ( n9850 , n9848 , n9849 );
xor ( n9851 , n9847 , n9850 );
nor ( n9852 , n796 , n686 );
xor ( n9853 , n9851 , n9852 );
and ( n9854 , n8971 , n8972 );
and ( n9855 , n8973 , n8976 );
or ( n9856 , n9854 , n9855 );
xor ( n9857 , n9853 , n9856 );
nor ( n9858 , n868 , n735 );
xor ( n9859 , n9857 , n9858 );
and ( n9860 , n8977 , n8978 );
and ( n9861 , n8979 , n8982 );
or ( n9862 , n9860 , n9861 );
xor ( n9863 , n9859 , n9862 );
nor ( n9864 , n958 , n798 );
xor ( n9865 , n9863 , n9864 );
and ( n9866 , n8983 , n8984 );
and ( n9867 , n8985 , n8988 );
or ( n9868 , n9866 , n9867 );
xor ( n9869 , n9865 , n9868 );
nor ( n9870 , n1062 , n870 );
xor ( n9871 , n9869 , n9870 );
and ( n9872 , n8989 , n8990 );
and ( n9873 , n8991 , n8994 );
or ( n9874 , n9872 , n9873 );
xor ( n9875 , n9871 , n9874 );
nor ( n9876 , n1176 , n960 );
xor ( n9877 , n9875 , n9876 );
and ( n9878 , n8995 , n8996 );
and ( n9879 , n8997 , n9000 );
or ( n9880 , n9878 , n9879 );
xor ( n9881 , n9877 , n9880 );
nor ( n9882 , n1303 , n1064 );
xor ( n9883 , n9881 , n9882 );
and ( n9884 , n9001 , n9002 );
and ( n9885 , n9003 , n9006 );
or ( n9886 , n9884 , n9885 );
xor ( n9887 , n9883 , n9886 );
nor ( n9888 , n1445 , n1178 );
xor ( n9889 , n9887 , n9888 );
and ( n9890 , n9007 , n9008 );
and ( n9891 , n9009 , n9012 );
or ( n9892 , n9890 , n9891 );
xor ( n9893 , n9889 , n9892 );
nor ( n9894 , n1598 , n1305 );
xor ( n9895 , n9893 , n9894 );
and ( n9896 , n9013 , n9014 );
and ( n9897 , n9015 , n9018 );
or ( n9898 , n9896 , n9897 );
xor ( n9899 , n9895 , n9898 );
nor ( n9900 , n1766 , n1447 );
xor ( n9901 , n9899 , n9900 );
and ( n9902 , n9019 , n9020 );
and ( n9903 , n9021 , n9024 );
or ( n9904 , n9902 , n9903 );
xor ( n9905 , n9901 , n9904 );
nor ( n9906 , n1945 , n1600 );
xor ( n9907 , n9905 , n9906 );
and ( n9908 , n9025 , n9026 );
and ( n9909 , n9027 , n9030 );
or ( n9910 , n9908 , n9909 );
xor ( n9911 , n9907 , n9910 );
nor ( n9912 , n2137 , n1768 );
xor ( n9913 , n9911 , n9912 );
and ( n9914 , n9031 , n9032 );
and ( n9915 , n9033 , n9036 );
or ( n9916 , n9914 , n9915 );
xor ( n9917 , n9913 , n9916 );
nor ( n9918 , n2343 , n1947 );
xor ( n9919 , n9917 , n9918 );
and ( n9920 , n9037 , n9038 );
and ( n9921 , n9039 , n9042 );
or ( n9922 , n9920 , n9921 );
xor ( n9923 , n9919 , n9922 );
nor ( n9924 , n2566 , n2139 );
xor ( n9925 , n9923 , n9924 );
and ( n9926 , n9043 , n9044 );
and ( n9927 , n9045 , n9048 );
or ( n9928 , n9926 , n9927 );
xor ( n9929 , n9925 , n9928 );
nor ( n9930 , n2797 , n2345 );
xor ( n9931 , n9929 , n9930 );
and ( n9932 , n9049 , n9050 );
and ( n9933 , n9051 , n9054 );
or ( n9934 , n9932 , n9933 );
xor ( n9935 , n9931 , n9934 );
nor ( n9936 , n3043 , n2568 );
xor ( n9937 , n9935 , n9936 );
and ( n9938 , n9055 , n9056 );
and ( n9939 , n9057 , n9060 );
or ( n9940 , n9938 , n9939 );
xor ( n9941 , n9937 , n9940 );
nor ( n9942 , n3300 , n2799 );
xor ( n9943 , n9941 , n9942 );
and ( n9944 , n9061 , n9062 );
and ( n9945 , n9063 , n9066 );
or ( n9946 , n9944 , n9945 );
xor ( n9947 , n9943 , n9946 );
nor ( n9948 , n3570 , n3045 );
xor ( n9949 , n9947 , n9948 );
and ( n9950 , n9067 , n9068 );
and ( n9951 , n9069 , n9072 );
or ( n9952 , n9950 , n9951 );
xor ( n9953 , n9949 , n9952 );
nor ( n9954 , n3853 , n3302 );
xor ( n9955 , n9953 , n9954 );
and ( n9956 , n9073 , n9074 );
and ( n9957 , n9075 , n9078 );
or ( n9958 , n9956 , n9957 );
xor ( n9959 , n9955 , n9958 );
nor ( n9960 , n4151 , n3572 );
xor ( n9961 , n9959 , n9960 );
and ( n9962 , n9079 , n9080 );
and ( n9963 , n9081 , n9084 );
or ( n9964 , n9962 , n9963 );
xor ( n9965 , n9961 , n9964 );
nor ( n9966 , n4458 , n3855 );
xor ( n9967 , n9965 , n9966 );
and ( n9968 , n9085 , n9086 );
and ( n9969 , n9087 , n9090 );
or ( n9970 , n9968 , n9969 );
xor ( n9971 , n9967 , n9970 );
nor ( n9972 , n4786 , n4153 );
xor ( n9973 , n9971 , n9972 );
and ( n9974 , n9091 , n9092 );
and ( n9975 , n9093 , n9096 );
or ( n9976 , n9974 , n9975 );
xor ( n9977 , n9973 , n9976 );
nor ( n9978 , n5126 , n4460 );
xor ( n9979 , n9977 , n9978 );
and ( n9980 , n9097 , n9098 );
and ( n9981 , n9099 , n9102 );
or ( n9982 , n9980 , n9981 );
xor ( n9983 , n9979 , n9982 );
nor ( n9984 , n5477 , n4788 );
xor ( n9985 , n9983 , n9984 );
and ( n9986 , n9103 , n9104 );
and ( n9987 , n9105 , n9108 );
or ( n9988 , n9986 , n9987 );
xor ( n9989 , n9985 , n9988 );
nor ( n9990 , n5838 , n5128 );
xor ( n9991 , n9989 , n9990 );
and ( n9992 , n9109 , n9110 );
and ( n9993 , n9111 , n9114 );
or ( n9994 , n9992 , n9993 );
xor ( n9995 , n9991 , n9994 );
nor ( n9996 , n6212 , n5479 );
xor ( n9997 , n9995 , n9996 );
and ( n9998 , n9115 , n9116 );
and ( n9999 , n9117 , n9120 );
or ( n10000 , n9998 , n9999 );
xor ( n10001 , n9997 , n10000 );
nor ( n10002 , n6596 , n5840 );
xor ( n10003 , n10001 , n10002 );
and ( n10004 , n9121 , n9122 );
and ( n10005 , n9123 , n9126 );
or ( n10006 , n10004 , n10005 );
xor ( n10007 , n10003 , n10006 );
nor ( n10008 , n6997 , n6214 );
xor ( n10009 , n10007 , n10008 );
and ( n10010 , n9127 , n9128 );
and ( n10011 , n9129 , n9132 );
or ( n10012 , n10010 , n10011 );
xor ( n10013 , n10009 , n10012 );
nor ( n10014 , n7413 , n6598 );
xor ( n10015 , n10013 , n10014 );
and ( n10016 , n9133 , n9134 );
and ( n10017 , n9135 , n9138 );
or ( n10018 , n10016 , n10017 );
xor ( n10019 , n10015 , n10018 );
nor ( n10020 , n7841 , n6999 );
xor ( n10021 , n10019 , n10020 );
and ( n10022 , n9139 , n9140 );
and ( n10023 , n9141 , n9144 );
or ( n10024 , n10022 , n10023 );
xor ( n10025 , n10021 , n10024 );
nor ( n10026 , n8281 , n7415 );
xor ( n10027 , n10025 , n10026 );
and ( n10028 , n9145 , n9146 );
and ( n10029 , n9147 , n9150 );
or ( n10030 , n10028 , n10029 );
xor ( n10031 , n10027 , n10030 );
nor ( n10032 , n8737 , n7843 );
xor ( n10033 , n10031 , n10032 );
and ( n10034 , n9151 , n9152 );
and ( n10035 , n9153 , n9156 );
or ( n10036 , n10034 , n10035 );
xor ( n10037 , n10033 , n10036 );
nor ( n10038 , n9420 , n8283 );
xor ( n10039 , n10037 , n10038 );
and ( n10040 , n9157 , n9158 );
and ( n10041 , n9159 , n9162 );
or ( n10042 , n10040 , n10041 );
xor ( n10043 , n10039 , n10042 );
and ( n10044 , n9385 , n9386 );
and ( n10045 , n9386 , n9405 );
and ( n10046 , n9385 , n9405 );
or ( n10047 , n10044 , n10045 , n10046 );
and ( n10048 , n9176 , n9380 );
and ( n10049 , n9380 , n9406 );
and ( n10050 , n9176 , n9406 );
or ( n10051 , n10048 , n10049 , n10050 );
xor ( n10052 , n10047 , n10051 );
and ( n10053 , n9180 , n9258 );
and ( n10054 , n9258 , n9379 );
and ( n10055 , n9180 , n9379 );
or ( n10056 , n10053 , n10054 , n10055 );
and ( n10057 , n9263 , n9307 );
and ( n10058 , n9307 , n9378 );
and ( n10059 , n9263 , n9378 );
or ( n10060 , n10057 , n10058 , n10059 );
and ( n10061 , n9193 , n9230 );
and ( n10062 , n9230 , n9256 );
and ( n10063 , n9193 , n9256 );
or ( n10064 , n10061 , n10062 , n10063 );
and ( n10065 , n9267 , n9271 );
and ( n10066 , n9271 , n9306 );
and ( n10067 , n9267 , n9306 );
or ( n10068 , n10065 , n10066 , n10067 );
xor ( n10069 , n10064 , n10068 );
and ( n10070 , n9235 , n9239 );
and ( n10071 , n9239 , n9255 );
and ( n10072 , n9235 , n9255 );
or ( n10073 , n10070 , n10071 , n10072 );
and ( n10074 , n9217 , n9222 );
and ( n10075 , n9222 , n9228 );
and ( n10076 , n9217 , n9228 );
or ( n10077 , n10074 , n10075 , n10076 );
and ( n10078 , n9207 , n9208 );
and ( n10079 , n9208 , n9210 );
and ( n10080 , n9207 , n9210 );
or ( n10081 , n10078 , n10079 , n10080 );
and ( n10082 , n9218 , n9219 );
and ( n10083 , n9219 , n9221 );
and ( n10084 , n9218 , n9221 );
or ( n10085 , n10082 , n10083 , n10084 );
xor ( n10086 , n10081 , n10085 );
and ( n10087 , n7385 , n719 );
and ( n10088 , n7808 , n663 );
xor ( n10089 , n10087 , n10088 );
and ( n10090 , n8079 , n635 );
xor ( n10091 , n10089 , n10090 );
xor ( n10092 , n10086 , n10091 );
xor ( n10093 , n10077 , n10092 );
and ( n10094 , n9224 , n9225 );
and ( n10095 , n9225 , n9227 );
and ( n10096 , n9224 , n9227 );
or ( n10097 , n10094 , n10095 , n10096 );
and ( n10098 , n6187 , n940 );
and ( n10099 , n6569 , n840 );
xor ( n10100 , n10098 , n10099 );
and ( n10101 , n6816 , n771 );
xor ( n10102 , n10100 , n10101 );
xor ( n10103 , n10097 , n10102 );
and ( n10104 , n4959 , n1254 );
and ( n10105 , n5459 , n1134 );
xor ( n10106 , n10104 , n10105 );
and ( n10107 , n5819 , n1034 );
xor ( n10108 , n10106 , n10107 );
xor ( n10109 , n10103 , n10108 );
xor ( n10110 , n10093 , n10109 );
xor ( n10111 , n10073 , n10110 );
and ( n10112 , n9244 , n9248 );
and ( n10113 , n9248 , n9254 );
and ( n10114 , n9244 , n9254 );
or ( n10115 , n10112 , n10113 , n10114 );
and ( n10116 , n9296 , n9301 );
and ( n10117 , n9301 , n9304 );
and ( n10118 , n9296 , n9304 );
or ( n10119 , n10116 , n10117 , n10118 );
xor ( n10120 , n10115 , n10119 );
and ( n10121 , n9250 , n9251 );
and ( n10122 , n9251 , n9253 );
and ( n10123 , n9250 , n9253 );
or ( n10124 , n10121 , n10122 , n10123 );
and ( n10125 , n9297 , n9298 );
and ( n10126 , n9298 , n9300 );
and ( n10127 , n9297 , n9300 );
or ( n10128 , n10125 , n10126 , n10127 );
xor ( n10129 , n10124 , n10128 );
and ( n10130 , n4132 , n1738 );
and ( n10131 , n4438 , n1551 );
xor ( n10132 , n10130 , n10131 );
and ( n10133 , n4766 , n1424 );
xor ( n10134 , n10132 , n10133 );
xor ( n10135 , n10129 , n10134 );
xor ( n10136 , n10120 , n10135 );
xor ( n10137 , n10111 , n10136 );
xor ( n10138 , n10069 , n10137 );
xor ( n10139 , n10060 , n10138 );
and ( n10140 , n9312 , n9338 );
and ( n10141 , n9338 , n9377 );
and ( n10142 , n9312 , n9377 );
or ( n10143 , n10140 , n10141 , n10142 );
and ( n10144 , n9276 , n9291 );
and ( n10145 , n9291 , n9305 );
and ( n10146 , n9276 , n9305 );
or ( n10147 , n10144 , n10145 , n10146 );
and ( n10148 , n9316 , n9320 );
and ( n10149 , n9320 , n9337 );
and ( n10150 , n9316 , n9337 );
or ( n10151 , n10148 , n10149 , n10150 );
xor ( n10152 , n10147 , n10151 );
and ( n10153 , n9280 , n9284 );
and ( n10154 , n9284 , n9290 );
and ( n10155 , n9280 , n9290 );
or ( n10156 , n10153 , n10154 , n10155 );
and ( n10157 , n9326 , n9327 );
and ( n10158 , n9327 , n9329 );
and ( n10159 , n9326 , n9329 );
or ( n10160 , n10157 , n10158 , n10159 );
and ( n10161 , n9286 , n9287 );
and ( n10162 , n9287 , n9289 );
and ( n10163 , n9286 , n9289 );
or ( n10164 , n10161 , n10162 , n10163 );
xor ( n10165 , n10160 , n10164 );
and ( n10166 , n1933 , n3749 );
and ( n10167 , n2120 , n3495 );
xor ( n10168 , n10166 , n10167 );
and ( n10169 , n2324 , n3271 );
xor ( n10170 , n10168 , n10169 );
xor ( n10171 , n10165 , n10170 );
xor ( n10172 , n10156 , n10171 );
and ( n10173 , n2462 , n2739 );
and ( n10174 , n2779 , n2544 );
and ( n10175 , n10173 , n10174 );
and ( n10176 , n10174 , n9303 );
and ( n10177 , n10173 , n9303 );
or ( n10178 , n10175 , n10176 , n10177 );
and ( n10179 , n3182 , n2298 );
and ( n10180 , n3545 , n2100 );
xor ( n10181 , n10179 , n10180 );
and ( n10182 , n3801 , n1882 );
xor ( n10183 , n10181 , n10182 );
xor ( n10184 , n10178 , n10183 );
and ( n10185 , n2462 , n2981 );
buf ( n10186 , n2779 );
xor ( n10187 , n10185 , n10186 );
and ( n10188 , n3024 , n2544 );
xor ( n10189 , n10187 , n10188 );
xor ( n10190 , n10184 , n10189 );
xor ( n10191 , n10172 , n10190 );
xor ( n10192 , n10152 , n10191 );
xor ( n10193 , n10143 , n10192 );
and ( n10194 , n9343 , n9360 );
and ( n10195 , n9360 , n9376 );
and ( n10196 , n9343 , n9376 );
or ( n10197 , n10194 , n10195 , n10196 );
and ( n10198 , n9365 , n9369 );
and ( n10199 , n9369 , n9375 );
and ( n10200 , n9365 , n9375 );
or ( n10201 , n10198 , n10199 , n10200 );
and ( n10202 , n9325 , n9330 );
and ( n10203 , n9330 , n9336 );
and ( n10204 , n9325 , n9336 );
or ( n10205 , n10202 , n10203 , n10204 );
xor ( n10206 , n10201 , n10205 );
and ( n10207 , n9332 , n9333 );
and ( n10208 , n9333 , n9335 );
and ( n10209 , n9332 , n9335 );
or ( n10210 , n10207 , n10208 , n10209 );
and ( n10211 , n1383 , n4730 );
and ( n10212 , n1580 , n4403 );
xor ( n10213 , n10211 , n10212 );
and ( n10214 , n1694 , n4102 );
xor ( n10215 , n10213 , n10214 );
xor ( n10216 , n10210 , n10215 );
and ( n10217 , n1047 , n5765 );
and ( n10218 , n1164 , n5408 );
xor ( n10219 , n10217 , n10218 );
and ( n10220 , n1287 , n5103 );
xor ( n10221 , n10219 , n10220 );
xor ( n10222 , n10216 , n10221 );
xor ( n10223 , n10206 , n10222 );
xor ( n10224 , n10197 , n10223 );
and ( n10225 , n9347 , n9353 );
and ( n10226 , n9353 , n9359 );
and ( n10227 , n9347 , n9359 );
or ( n10228 , n10225 , n10226 , n10227 );
and ( n10229 , n9349 , n9350 );
and ( n10230 , n9350 , n9352 );
and ( n10231 , n9349 , n9352 );
or ( n10232 , n10229 , n10230 , n10231 );
and ( n10233 , n632 , n8243 );
and ( n10234 , n671 , n7662 );
xor ( n10235 , n10233 , n10234 );
and ( n10236 , n715 , n7310 );
xor ( n10237 , n10235 , n10236 );
xor ( n10238 , n10232 , n10237 );
buf ( n10239 , n432 );
and ( n10240 , n599 , n10239 );
and ( n10241 , n608 , n9348 );
xor ( n10242 , n10240 , n10241 );
and ( n10243 , n611 , n8669 );
xor ( n10244 , n10242 , n10243 );
xor ( n10245 , n10238 , n10244 );
xor ( n10246 , n10228 , n10245 );
and ( n10247 , n9355 , n9356 );
and ( n10248 , n9356 , n9358 );
and ( n10249 , n9355 , n9358 );
or ( n10250 , n10247 , n10248 , n10249 );
and ( n10251 , n9371 , n9372 );
and ( n10252 , n9372 , n9374 );
and ( n10253 , n9371 , n9374 );
or ( n10254 , n10251 , n10252 , n10253 );
xor ( n10255 , n10250 , n10254 );
and ( n10256 , n783 , n6971 );
and ( n10257 , n856 , n6504 );
xor ( n10258 , n10256 , n10257 );
and ( n10259 , n925 , n6132 );
xor ( n10260 , n10258 , n10259 );
xor ( n10261 , n10255 , n10260 );
xor ( n10262 , n10246 , n10261 );
xor ( n10263 , n10224 , n10262 );
xor ( n10264 , n10193 , n10263 );
xor ( n10265 , n10139 , n10264 );
xor ( n10266 , n10056 , n10265 );
and ( n10267 , n9184 , n9188 );
and ( n10268 , n9188 , n9257 );
and ( n10269 , n9184 , n9257 );
or ( n10270 , n10267 , n10268 , n10269 );
and ( n10271 , n9388 , n9404 );
xor ( n10272 , n10270 , n10271 );
and ( n10273 , n9392 , n9393 );
and ( n10274 , n9393 , n9403 );
and ( n10275 , n9392 , n9403 );
or ( n10276 , n10273 , n10274 , n10275 );
and ( n10277 , n9197 , n9212 );
and ( n10278 , n9212 , n9229 );
and ( n10279 , n9197 , n9229 );
or ( n10280 , n10277 , n10278 , n10279 );
and ( n10281 , n9398 , n9402 );
xor ( n10282 , n10280 , n10281 );
and ( n10283 , n9201 , n9205 );
and ( n10284 , n9205 , n9211 );
and ( n10285 , n9201 , n9211 );
or ( n10286 , n10283 , n10284 , n10285 );
and ( n10287 , n9399 , n9401 );
and ( n10288 , n8718 , n606 );
and ( n10289 , n9400 , n615 );
xor ( n10290 , n10288 , n10289 );
buf ( n10291 , n432 );
and ( n10292 , n10291 , n612 );
xor ( n10293 , n10290 , n10292 );
xor ( n10294 , n10287 , n10293 );
xor ( n10295 , n10286 , n10294 );
xor ( n10296 , n10282 , n10295 );
xor ( n10297 , n10276 , n10296 );
xor ( n10298 , n10272 , n10297 );
xor ( n10299 , n10266 , n10298 );
xor ( n10300 , n10052 , n10299 );
and ( n10301 , n9167 , n9171 );
and ( n10302 , n9171 , n9407 );
and ( n10303 , n9167 , n9407 );
or ( n10304 , n10301 , n10302 , n10303 );
xor ( n10305 , n10300 , n10304 );
and ( n10306 , n9408 , n9412 );
and ( n10307 , n9413 , n9416 );
or ( n10308 , n10306 , n10307 );
xor ( n10309 , n10305 , n10308 );
buf ( n10310 , n10309 );
buf ( n10311 , n10310 );
not ( n10312 , n10311 );
nor ( n10313 , n10312 , n8739 );
xor ( n10314 , n10043 , n10313 );
and ( n10315 , n9163 , n9421 );
and ( n10316 , n9422 , n9425 );
or ( n10317 , n10315 , n10316 );
xor ( n10318 , n10314 , n10317 );
buf ( n10319 , n10318 );
buf ( n10320 , n10319 );
not ( n10321 , n10320 );
buf ( n10322 , n537 );
not ( n10323 , n10322 );
nor ( n10324 , n10321 , n10323 );
xor ( n10325 , n9827 , n10324 );
xor ( n10326 , n9442 , n9824 );
nor ( n10327 , n9429 , n10323 );
and ( n10328 , n10326 , n10327 );
xor ( n10329 , n10326 , n10327 );
xor ( n10330 , n9451 , n9822 );
nor ( n10331 , n8949 , n10323 );
and ( n10332 , n10330 , n10331 );
xor ( n10333 , n10330 , n10331 );
xor ( n10334 , n9460 , n9820 );
nor ( n10335 , n9437 , n10323 );
and ( n10336 , n10334 , n10335 );
xor ( n10337 , n10334 , n10335 );
xor ( n10338 , n9469 , n9818 );
nor ( n10339 , n9446 , n10323 );
and ( n10340 , n10338 , n10339 );
xor ( n10341 , n10338 , n10339 );
xor ( n10342 , n9478 , n9816 );
nor ( n10343 , n9455 , n10323 );
and ( n10344 , n10342 , n10343 );
xor ( n10345 , n10342 , n10343 );
xor ( n10346 , n9487 , n9814 );
nor ( n10347 , n9464 , n10323 );
and ( n10348 , n10346 , n10347 );
xor ( n10349 , n10346 , n10347 );
xor ( n10350 , n9496 , n9812 );
nor ( n10351 , n9473 , n10323 );
and ( n10352 , n10350 , n10351 );
xor ( n10353 , n10350 , n10351 );
xor ( n10354 , n9505 , n9810 );
nor ( n10355 , n9482 , n10323 );
and ( n10356 , n10354 , n10355 );
xor ( n10357 , n10354 , n10355 );
xor ( n10358 , n9514 , n9808 );
nor ( n10359 , n9491 , n10323 );
and ( n10360 , n10358 , n10359 );
xor ( n10361 , n10358 , n10359 );
xor ( n10362 , n9523 , n9806 );
nor ( n10363 , n9500 , n10323 );
and ( n10364 , n10362 , n10363 );
xor ( n10365 , n10362 , n10363 );
xor ( n10366 , n9532 , n9804 );
nor ( n10367 , n9509 , n10323 );
and ( n10368 , n10366 , n10367 );
xor ( n10369 , n10366 , n10367 );
xor ( n10370 , n9541 , n9802 );
nor ( n10371 , n9518 , n10323 );
and ( n10372 , n10370 , n10371 );
xor ( n10373 , n10370 , n10371 );
xor ( n10374 , n9550 , n9800 );
nor ( n10375 , n9527 , n10323 );
and ( n10376 , n10374 , n10375 );
xor ( n10377 , n10374 , n10375 );
xor ( n10378 , n9559 , n9798 );
nor ( n10379 , n9536 , n10323 );
and ( n10380 , n10378 , n10379 );
xor ( n10381 , n10378 , n10379 );
xor ( n10382 , n9568 , n9796 );
nor ( n10383 , n9545 , n10323 );
and ( n10384 , n10382 , n10383 );
xor ( n10385 , n10382 , n10383 );
xor ( n10386 , n9577 , n9794 );
nor ( n10387 , n9554 , n10323 );
and ( n10388 , n10386 , n10387 );
xor ( n10389 , n10386 , n10387 );
xor ( n10390 , n9586 , n9792 );
nor ( n10391 , n9563 , n10323 );
and ( n10392 , n10390 , n10391 );
xor ( n10393 , n10390 , n10391 );
xor ( n10394 , n9595 , n9790 );
nor ( n10395 , n9572 , n10323 );
and ( n10396 , n10394 , n10395 );
xor ( n10397 , n10394 , n10395 );
xor ( n10398 , n9604 , n9788 );
nor ( n10399 , n9581 , n10323 );
and ( n10400 , n10398 , n10399 );
xor ( n10401 , n10398 , n10399 );
xor ( n10402 , n9613 , n9786 );
nor ( n10403 , n9590 , n10323 );
and ( n10404 , n10402 , n10403 );
xor ( n10405 , n10402 , n10403 );
xor ( n10406 , n9622 , n9784 );
nor ( n10407 , n9599 , n10323 );
and ( n10408 , n10406 , n10407 );
xor ( n10409 , n10406 , n10407 );
xor ( n10410 , n9631 , n9782 );
nor ( n10411 , n9608 , n10323 );
and ( n10412 , n10410 , n10411 );
xor ( n10413 , n10410 , n10411 );
xor ( n10414 , n9640 , n9780 );
nor ( n10415 , n9617 , n10323 );
and ( n10416 , n10414 , n10415 );
xor ( n10417 , n10414 , n10415 );
xor ( n10418 , n9649 , n9778 );
nor ( n10419 , n9626 , n10323 );
and ( n10420 , n10418 , n10419 );
xor ( n10421 , n10418 , n10419 );
xor ( n10422 , n9658 , n9776 );
nor ( n10423 , n9635 , n10323 );
and ( n10424 , n10422 , n10423 );
xor ( n10425 , n10422 , n10423 );
xor ( n10426 , n9667 , n9774 );
nor ( n10427 , n9644 , n10323 );
and ( n10428 , n10426 , n10427 );
xor ( n10429 , n10426 , n10427 );
xor ( n10430 , n9676 , n9772 );
nor ( n10431 , n9653 , n10323 );
and ( n10432 , n10430 , n10431 );
xor ( n10433 , n10430 , n10431 );
xor ( n10434 , n9685 , n9770 );
nor ( n10435 , n9662 , n10323 );
and ( n10436 , n10434 , n10435 );
xor ( n10437 , n10434 , n10435 );
xor ( n10438 , n9694 , n9768 );
nor ( n10439 , n9671 , n10323 );
and ( n10440 , n10438 , n10439 );
xor ( n10441 , n10438 , n10439 );
xor ( n10442 , n9703 , n9766 );
nor ( n10443 , n9680 , n10323 );
and ( n10444 , n10442 , n10443 );
xor ( n10445 , n10442 , n10443 );
xor ( n10446 , n9712 , n9764 );
nor ( n10447 , n9689 , n10323 );
and ( n10448 , n10446 , n10447 );
xor ( n10449 , n10446 , n10447 );
xor ( n10450 , n9721 , n9762 );
nor ( n10451 , n9698 , n10323 );
and ( n10452 , n10450 , n10451 );
xor ( n10453 , n10450 , n10451 );
xor ( n10454 , n9730 , n9760 );
nor ( n10455 , n9707 , n10323 );
and ( n10456 , n10454 , n10455 );
xor ( n10457 , n10454 , n10455 );
xor ( n10458 , n9739 , n9758 );
nor ( n10459 , n9716 , n10323 );
and ( n10460 , n10458 , n10459 );
xor ( n10461 , n10458 , n10459 );
xor ( n10462 , n9748 , n9756 );
nor ( n10463 , n9725 , n10323 );
and ( n10464 , n10462 , n10463 );
xor ( n10465 , n10462 , n10463 );
xor ( n10466 , n9754 , n9755 );
nor ( n10467 , n9734 , n10323 );
and ( n10468 , n10466 , n10467 );
xor ( n10469 , n10466 , n10467 );
nor ( n10470 , n9752 , n9431 );
nor ( n10471 , n9743 , n10323 );
and ( n10472 , n10470 , n10471 );
and ( n10473 , n10469 , n10472 );
or ( n10474 , n10468 , n10473 );
and ( n10475 , n10465 , n10474 );
or ( n10476 , n10464 , n10475 );
and ( n10477 , n10461 , n10476 );
or ( n10478 , n10460 , n10477 );
and ( n10479 , n10457 , n10478 );
or ( n10480 , n10456 , n10479 );
and ( n10481 , n10453 , n10480 );
or ( n10482 , n10452 , n10481 );
and ( n10483 , n10449 , n10482 );
or ( n10484 , n10448 , n10483 );
and ( n10485 , n10445 , n10484 );
or ( n10486 , n10444 , n10485 );
and ( n10487 , n10441 , n10486 );
or ( n10488 , n10440 , n10487 );
and ( n10489 , n10437 , n10488 );
or ( n10490 , n10436 , n10489 );
and ( n10491 , n10433 , n10490 );
or ( n10492 , n10432 , n10491 );
and ( n10493 , n10429 , n10492 );
or ( n10494 , n10428 , n10493 );
and ( n10495 , n10425 , n10494 );
or ( n10496 , n10424 , n10495 );
and ( n10497 , n10421 , n10496 );
or ( n10498 , n10420 , n10497 );
and ( n10499 , n10417 , n10498 );
or ( n10500 , n10416 , n10499 );
and ( n10501 , n10413 , n10500 );
or ( n10502 , n10412 , n10501 );
and ( n10503 , n10409 , n10502 );
or ( n10504 , n10408 , n10503 );
and ( n10505 , n10405 , n10504 );
or ( n10506 , n10404 , n10505 );
and ( n10507 , n10401 , n10506 );
or ( n10508 , n10400 , n10507 );
and ( n10509 , n10397 , n10508 );
or ( n10510 , n10396 , n10509 );
and ( n10511 , n10393 , n10510 );
or ( n10512 , n10392 , n10511 );
and ( n10513 , n10389 , n10512 );
or ( n10514 , n10388 , n10513 );
and ( n10515 , n10385 , n10514 );
or ( n10516 , n10384 , n10515 );
and ( n10517 , n10381 , n10516 );
or ( n10518 , n10380 , n10517 );
and ( n10519 , n10377 , n10518 );
or ( n10520 , n10376 , n10519 );
and ( n10521 , n10373 , n10520 );
or ( n10522 , n10372 , n10521 );
and ( n10523 , n10369 , n10522 );
or ( n10524 , n10368 , n10523 );
and ( n10525 , n10365 , n10524 );
or ( n10526 , n10364 , n10525 );
and ( n10527 , n10361 , n10526 );
or ( n10528 , n10360 , n10527 );
and ( n10529 , n10357 , n10528 );
or ( n10530 , n10356 , n10529 );
and ( n10531 , n10353 , n10530 );
or ( n10532 , n10352 , n10531 );
and ( n10533 , n10349 , n10532 );
or ( n10534 , n10348 , n10533 );
and ( n10535 , n10345 , n10534 );
or ( n10536 , n10344 , n10535 );
and ( n10537 , n10341 , n10536 );
or ( n10538 , n10340 , n10537 );
and ( n10539 , n10337 , n10538 );
or ( n10540 , n10336 , n10539 );
and ( n10541 , n10333 , n10540 );
or ( n10542 , n10332 , n10541 );
and ( n10543 , n10329 , n10542 );
or ( n10544 , n10328 , n10543 );
xor ( n10545 , n10325 , n10544 );
buf ( n10546 , n495 );
not ( n10547 , n10546 );
nor ( n10548 , n601 , n10547 );
buf ( n10549 , n10548 );
nor ( n10550 , n622 , n8955 );
xor ( n10551 , n10549 , n10550 );
buf ( n10552 , n10551 );
nor ( n10553 , n646 , n603 );
xor ( n10554 , n10552 , n10553 );
and ( n10555 , n9831 , n9832 );
buf ( n10556 , n10555 );
xor ( n10557 , n10554 , n10556 );
nor ( n10558 , n684 , n652 );
xor ( n10559 , n10557 , n10558 );
and ( n10560 , n9834 , n9835 );
and ( n10561 , n9836 , n9838 );
or ( n10562 , n10560 , n10561 );
xor ( n10563 , n10559 , n10562 );
nor ( n10564 , n733 , n624 );
xor ( n10565 , n10563 , n10564 );
and ( n10566 , n9839 , n9840 );
and ( n10567 , n9841 , n9844 );
or ( n10568 , n10566 , n10567 );
xor ( n10569 , n10565 , n10568 );
nor ( n10570 , n796 , n648 );
xor ( n10571 , n10569 , n10570 );
and ( n10572 , n9845 , n9846 );
and ( n10573 , n9847 , n9850 );
or ( n10574 , n10572 , n10573 );
xor ( n10575 , n10571 , n10574 );
nor ( n10576 , n868 , n686 );
xor ( n10577 , n10575 , n10576 );
and ( n10578 , n9851 , n9852 );
and ( n10579 , n9853 , n9856 );
or ( n10580 , n10578 , n10579 );
xor ( n10581 , n10577 , n10580 );
nor ( n10582 , n958 , n735 );
xor ( n10583 , n10581 , n10582 );
and ( n10584 , n9857 , n9858 );
and ( n10585 , n9859 , n9862 );
or ( n10586 , n10584 , n10585 );
xor ( n10587 , n10583 , n10586 );
nor ( n10588 , n1062 , n798 );
xor ( n10589 , n10587 , n10588 );
and ( n10590 , n9863 , n9864 );
and ( n10591 , n9865 , n9868 );
or ( n10592 , n10590 , n10591 );
xor ( n10593 , n10589 , n10592 );
nor ( n10594 , n1176 , n870 );
xor ( n10595 , n10593 , n10594 );
and ( n10596 , n9869 , n9870 );
and ( n10597 , n9871 , n9874 );
or ( n10598 , n10596 , n10597 );
xor ( n10599 , n10595 , n10598 );
nor ( n10600 , n1303 , n960 );
xor ( n10601 , n10599 , n10600 );
and ( n10602 , n9875 , n9876 );
and ( n10603 , n9877 , n9880 );
or ( n10604 , n10602 , n10603 );
xor ( n10605 , n10601 , n10604 );
nor ( n10606 , n1445 , n1064 );
xor ( n10607 , n10605 , n10606 );
and ( n10608 , n9881 , n9882 );
and ( n10609 , n9883 , n9886 );
or ( n10610 , n10608 , n10609 );
xor ( n10611 , n10607 , n10610 );
nor ( n10612 , n1598 , n1178 );
xor ( n10613 , n10611 , n10612 );
and ( n10614 , n9887 , n9888 );
and ( n10615 , n9889 , n9892 );
or ( n10616 , n10614 , n10615 );
xor ( n10617 , n10613 , n10616 );
nor ( n10618 , n1766 , n1305 );
xor ( n10619 , n10617 , n10618 );
and ( n10620 , n9893 , n9894 );
and ( n10621 , n9895 , n9898 );
or ( n10622 , n10620 , n10621 );
xor ( n10623 , n10619 , n10622 );
nor ( n10624 , n1945 , n1447 );
xor ( n10625 , n10623 , n10624 );
and ( n10626 , n9899 , n9900 );
and ( n10627 , n9901 , n9904 );
or ( n10628 , n10626 , n10627 );
xor ( n10629 , n10625 , n10628 );
nor ( n10630 , n2137 , n1600 );
xor ( n10631 , n10629 , n10630 );
and ( n10632 , n9905 , n9906 );
and ( n10633 , n9907 , n9910 );
or ( n10634 , n10632 , n10633 );
xor ( n10635 , n10631 , n10634 );
nor ( n10636 , n2343 , n1768 );
xor ( n10637 , n10635 , n10636 );
and ( n10638 , n9911 , n9912 );
and ( n10639 , n9913 , n9916 );
or ( n10640 , n10638 , n10639 );
xor ( n10641 , n10637 , n10640 );
nor ( n10642 , n2566 , n1947 );
xor ( n10643 , n10641 , n10642 );
and ( n10644 , n9917 , n9918 );
and ( n10645 , n9919 , n9922 );
or ( n10646 , n10644 , n10645 );
xor ( n10647 , n10643 , n10646 );
nor ( n10648 , n2797 , n2139 );
xor ( n10649 , n10647 , n10648 );
and ( n10650 , n9923 , n9924 );
and ( n10651 , n9925 , n9928 );
or ( n10652 , n10650 , n10651 );
xor ( n10653 , n10649 , n10652 );
nor ( n10654 , n3043 , n2345 );
xor ( n10655 , n10653 , n10654 );
and ( n10656 , n9929 , n9930 );
and ( n10657 , n9931 , n9934 );
or ( n10658 , n10656 , n10657 );
xor ( n10659 , n10655 , n10658 );
nor ( n10660 , n3300 , n2568 );
xor ( n10661 , n10659 , n10660 );
and ( n10662 , n9935 , n9936 );
and ( n10663 , n9937 , n9940 );
or ( n10664 , n10662 , n10663 );
xor ( n10665 , n10661 , n10664 );
nor ( n10666 , n3570 , n2799 );
xor ( n10667 , n10665 , n10666 );
and ( n10668 , n9941 , n9942 );
and ( n10669 , n9943 , n9946 );
or ( n10670 , n10668 , n10669 );
xor ( n10671 , n10667 , n10670 );
nor ( n10672 , n3853 , n3045 );
xor ( n10673 , n10671 , n10672 );
and ( n10674 , n9947 , n9948 );
and ( n10675 , n9949 , n9952 );
or ( n10676 , n10674 , n10675 );
xor ( n10677 , n10673 , n10676 );
nor ( n10678 , n4151 , n3302 );
xor ( n10679 , n10677 , n10678 );
and ( n10680 , n9953 , n9954 );
and ( n10681 , n9955 , n9958 );
or ( n10682 , n10680 , n10681 );
xor ( n10683 , n10679 , n10682 );
nor ( n10684 , n4458 , n3572 );
xor ( n10685 , n10683 , n10684 );
and ( n10686 , n9959 , n9960 );
and ( n10687 , n9961 , n9964 );
or ( n10688 , n10686 , n10687 );
xor ( n10689 , n10685 , n10688 );
nor ( n10690 , n4786 , n3855 );
xor ( n10691 , n10689 , n10690 );
and ( n10692 , n9965 , n9966 );
and ( n10693 , n9967 , n9970 );
or ( n10694 , n10692 , n10693 );
xor ( n10695 , n10691 , n10694 );
nor ( n10696 , n5126 , n4153 );
xor ( n10697 , n10695 , n10696 );
and ( n10698 , n9971 , n9972 );
and ( n10699 , n9973 , n9976 );
or ( n10700 , n10698 , n10699 );
xor ( n10701 , n10697 , n10700 );
nor ( n10702 , n5477 , n4460 );
xor ( n10703 , n10701 , n10702 );
and ( n10704 , n9977 , n9978 );
and ( n10705 , n9979 , n9982 );
or ( n10706 , n10704 , n10705 );
xor ( n10707 , n10703 , n10706 );
nor ( n10708 , n5838 , n4788 );
xor ( n10709 , n10707 , n10708 );
and ( n10710 , n9983 , n9984 );
and ( n10711 , n9985 , n9988 );
or ( n10712 , n10710 , n10711 );
xor ( n10713 , n10709 , n10712 );
nor ( n10714 , n6212 , n5128 );
xor ( n10715 , n10713 , n10714 );
and ( n10716 , n9989 , n9990 );
and ( n10717 , n9991 , n9994 );
or ( n10718 , n10716 , n10717 );
xor ( n10719 , n10715 , n10718 );
nor ( n10720 , n6596 , n5479 );
xor ( n10721 , n10719 , n10720 );
and ( n10722 , n9995 , n9996 );
and ( n10723 , n9997 , n10000 );
or ( n10724 , n10722 , n10723 );
xor ( n10725 , n10721 , n10724 );
nor ( n10726 , n6997 , n5840 );
xor ( n10727 , n10725 , n10726 );
and ( n10728 , n10001 , n10002 );
and ( n10729 , n10003 , n10006 );
or ( n10730 , n10728 , n10729 );
xor ( n10731 , n10727 , n10730 );
nor ( n10732 , n7413 , n6214 );
xor ( n10733 , n10731 , n10732 );
and ( n10734 , n10007 , n10008 );
and ( n10735 , n10009 , n10012 );
or ( n10736 , n10734 , n10735 );
xor ( n10737 , n10733 , n10736 );
nor ( n10738 , n7841 , n6598 );
xor ( n10739 , n10737 , n10738 );
and ( n10740 , n10013 , n10014 );
and ( n10741 , n10015 , n10018 );
or ( n10742 , n10740 , n10741 );
xor ( n10743 , n10739 , n10742 );
nor ( n10744 , n8281 , n6999 );
xor ( n10745 , n10743 , n10744 );
and ( n10746 , n10019 , n10020 );
and ( n10747 , n10021 , n10024 );
or ( n10748 , n10746 , n10747 );
xor ( n10749 , n10745 , n10748 );
nor ( n10750 , n8737 , n7415 );
xor ( n10751 , n10749 , n10750 );
and ( n10752 , n10025 , n10026 );
and ( n10753 , n10027 , n10030 );
or ( n10754 , n10752 , n10753 );
xor ( n10755 , n10751 , n10754 );
nor ( n10756 , n9420 , n7843 );
xor ( n10757 , n10755 , n10756 );
and ( n10758 , n10031 , n10032 );
and ( n10759 , n10033 , n10036 );
or ( n10760 , n10758 , n10759 );
xor ( n10761 , n10757 , n10760 );
nor ( n10762 , n10312 , n8283 );
xor ( n10763 , n10761 , n10762 );
and ( n10764 , n10037 , n10038 );
and ( n10765 , n10039 , n10042 );
or ( n10766 , n10764 , n10765 );
xor ( n10767 , n10763 , n10766 );
and ( n10768 , n10270 , n10271 );
and ( n10769 , n10271 , n10297 );
and ( n10770 , n10270 , n10297 );
or ( n10771 , n10768 , n10769 , n10770 );
and ( n10772 , n10056 , n10265 );
and ( n10773 , n10265 , n10298 );
and ( n10774 , n10056 , n10298 );
or ( n10775 , n10772 , n10773 , n10774 );
xor ( n10776 , n10771 , n10775 );
and ( n10777 , n10060 , n10138 );
and ( n10778 , n10138 , n10264 );
and ( n10779 , n10060 , n10264 );
or ( n10780 , n10777 , n10778 , n10779 );
and ( n10781 , n10143 , n10192 );
and ( n10782 , n10192 , n10263 );
and ( n10783 , n10143 , n10263 );
or ( n10784 , n10781 , n10782 , n10783 );
and ( n10785 , n10073 , n10110 );
and ( n10786 , n10110 , n10136 );
and ( n10787 , n10073 , n10136 );
or ( n10788 , n10785 , n10786 , n10787 );
and ( n10789 , n10147 , n10151 );
and ( n10790 , n10151 , n10191 );
and ( n10791 , n10147 , n10191 );
or ( n10792 , n10789 , n10790 , n10791 );
xor ( n10793 , n10788 , n10792 );
and ( n10794 , n10115 , n10119 );
and ( n10795 , n10119 , n10135 );
and ( n10796 , n10115 , n10135 );
or ( n10797 , n10794 , n10795 , n10796 );
and ( n10798 , n10097 , n10102 );
and ( n10799 , n10102 , n10108 );
and ( n10800 , n10097 , n10108 );
or ( n10801 , n10798 , n10799 , n10800 );
and ( n10802 , n10087 , n10088 );
and ( n10803 , n10088 , n10090 );
and ( n10804 , n10087 , n10090 );
or ( n10805 , n10802 , n10803 , n10804 );
and ( n10806 , n10098 , n10099 );
and ( n10807 , n10099 , n10101 );
and ( n10808 , n10098 , n10101 );
or ( n10809 , n10806 , n10807 , n10808 );
xor ( n10810 , n10805 , n10809 );
and ( n10811 , n7385 , n771 );
and ( n10812 , n7808 , n719 );
xor ( n10813 , n10811 , n10812 );
and ( n10814 , n8079 , n663 );
xor ( n10815 , n10813 , n10814 );
xor ( n10816 , n10810 , n10815 );
xor ( n10817 , n10801 , n10816 );
and ( n10818 , n10104 , n10105 );
and ( n10819 , n10105 , n10107 );
and ( n10820 , n10104 , n10107 );
or ( n10821 , n10818 , n10819 , n10820 );
and ( n10822 , n6187 , n1034 );
and ( n10823 , n6569 , n940 );
xor ( n10824 , n10822 , n10823 );
and ( n10825 , n6816 , n840 );
xor ( n10826 , n10824 , n10825 );
xor ( n10827 , n10821 , n10826 );
and ( n10828 , n4959 , n1424 );
and ( n10829 , n5459 , n1254 );
xor ( n10830 , n10828 , n10829 );
and ( n10831 , n5819 , n1134 );
xor ( n10832 , n10830 , n10831 );
xor ( n10833 , n10827 , n10832 );
xor ( n10834 , n10817 , n10833 );
xor ( n10835 , n10797 , n10834 );
and ( n10836 , n10124 , n10128 );
and ( n10837 , n10128 , n10134 );
and ( n10838 , n10124 , n10134 );
or ( n10839 , n10836 , n10837 , n10838 );
and ( n10840 , n10178 , n10183 );
and ( n10841 , n10183 , n10189 );
and ( n10842 , n10178 , n10189 );
or ( n10843 , n10840 , n10841 , n10842 );
xor ( n10844 , n10839 , n10843 );
and ( n10845 , n10130 , n10131 );
and ( n10846 , n10131 , n10133 );
and ( n10847 , n10130 , n10133 );
or ( n10848 , n10845 , n10846 , n10847 );
and ( n10849 , n10179 , n10180 );
and ( n10850 , n10180 , n10182 );
and ( n10851 , n10179 , n10182 );
or ( n10852 , n10849 , n10850 , n10851 );
xor ( n10853 , n10848 , n10852 );
and ( n10854 , n4132 , n1882 );
and ( n10855 , n4438 , n1738 );
xor ( n10856 , n10854 , n10855 );
and ( n10857 , n4766 , n1551 );
xor ( n10858 , n10856 , n10857 );
xor ( n10859 , n10853 , n10858 );
xor ( n10860 , n10844 , n10859 );
xor ( n10861 , n10835 , n10860 );
xor ( n10862 , n10793 , n10861 );
xor ( n10863 , n10784 , n10862 );
and ( n10864 , n10197 , n10223 );
and ( n10865 , n10223 , n10262 );
and ( n10866 , n10197 , n10262 );
or ( n10867 , n10864 , n10865 , n10866 );
and ( n10868 , n10156 , n10171 );
and ( n10869 , n10171 , n10190 );
and ( n10870 , n10156 , n10190 );
or ( n10871 , n10868 , n10869 , n10870 );
and ( n10872 , n10201 , n10205 );
and ( n10873 , n10205 , n10222 );
and ( n10874 , n10201 , n10222 );
or ( n10875 , n10872 , n10873 , n10874 );
xor ( n10876 , n10871 , n10875 );
and ( n10877 , n10160 , n10164 );
and ( n10878 , n10164 , n10170 );
and ( n10879 , n10160 , n10170 );
or ( n10880 , n10877 , n10878 , n10879 );
and ( n10881 , n10185 , n10186 );
and ( n10882 , n10186 , n10188 );
and ( n10883 , n10185 , n10188 );
or ( n10884 , n10881 , n10882 , n10883 );
and ( n10885 , n3182 , n2544 );
and ( n10886 , n3545 , n2298 );
xor ( n10887 , n10885 , n10886 );
and ( n10888 , n3801 , n2100 );
xor ( n10889 , n10887 , n10888 );
xor ( n10890 , n10884 , n10889 );
and ( n10891 , n2462 , n3271 );
and ( n10892 , n2779 , n2981 );
xor ( n10893 , n10891 , n10892 );
and ( n10894 , n3024 , n2739 );
xor ( n10895 , n10893 , n10894 );
xor ( n10896 , n10890 , n10895 );
xor ( n10897 , n10880 , n10896 );
and ( n10898 , n10166 , n10167 );
and ( n10899 , n10167 , n10169 );
and ( n10900 , n10166 , n10169 );
or ( n10901 , n10898 , n10899 , n10900 );
and ( n10902 , n10211 , n10212 );
and ( n10903 , n10212 , n10214 );
and ( n10904 , n10211 , n10214 );
or ( n10905 , n10902 , n10903 , n10904 );
xor ( n10906 , n10901 , n10905 );
and ( n10907 , n1933 , n4102 );
and ( n10908 , n2120 , n3749 );
xor ( n10909 , n10907 , n10908 );
and ( n10910 , n2324 , n3495 );
xor ( n10911 , n10909 , n10910 );
xor ( n10912 , n10906 , n10911 );
xor ( n10913 , n10897 , n10912 );
xor ( n10914 , n10876 , n10913 );
xor ( n10915 , n10867 , n10914 );
and ( n10916 , n10228 , n10245 );
and ( n10917 , n10245 , n10261 );
and ( n10918 , n10228 , n10261 );
or ( n10919 , n10916 , n10917 , n10918 );
and ( n10920 , n10250 , n10254 );
and ( n10921 , n10254 , n10260 );
and ( n10922 , n10250 , n10260 );
or ( n10923 , n10920 , n10921 , n10922 );
and ( n10924 , n10210 , n10215 );
and ( n10925 , n10215 , n10221 );
and ( n10926 , n10210 , n10221 );
or ( n10927 , n10924 , n10925 , n10926 );
xor ( n10928 , n10923 , n10927 );
and ( n10929 , n10217 , n10218 );
and ( n10930 , n10218 , n10220 );
and ( n10931 , n10217 , n10220 );
or ( n10932 , n10929 , n10930 , n10931 );
and ( n10933 , n1383 , n5103 );
and ( n10934 , n1580 , n4730 );
xor ( n10935 , n10933 , n10934 );
and ( n10936 , n1694 , n4403 );
xor ( n10937 , n10935 , n10936 );
xor ( n10938 , n10932 , n10937 );
and ( n10939 , n1047 , n6132 );
and ( n10940 , n1164 , n5765 );
xor ( n10941 , n10939 , n10940 );
and ( n10942 , n1287 , n5408 );
xor ( n10943 , n10941 , n10942 );
xor ( n10944 , n10938 , n10943 );
xor ( n10945 , n10928 , n10944 );
xor ( n10946 , n10919 , n10945 );
and ( n10947 , n10232 , n10237 );
and ( n10948 , n10237 , n10244 );
and ( n10949 , n10232 , n10244 );
or ( n10950 , n10947 , n10948 , n10949 );
and ( n10951 , n10256 , n10257 );
and ( n10952 , n10257 , n10259 );
and ( n10953 , n10256 , n10259 );
or ( n10954 , n10951 , n10952 , n10953 );
and ( n10955 , n10233 , n10234 );
and ( n10956 , n10234 , n10236 );
and ( n10957 , n10233 , n10236 );
or ( n10958 , n10955 , n10956 , n10957 );
xor ( n10959 , n10954 , n10958 );
and ( n10960 , n783 , n7310 );
and ( n10961 , n856 , n6971 );
xor ( n10962 , n10960 , n10961 );
and ( n10963 , n925 , n6504 );
xor ( n10964 , n10962 , n10963 );
xor ( n10965 , n10959 , n10964 );
xor ( n10966 , n10950 , n10965 );
and ( n10967 , n10240 , n10241 );
and ( n10968 , n10241 , n10243 );
and ( n10969 , n10240 , n10243 );
or ( n10970 , n10967 , n10968 , n10969 );
and ( n10971 , n632 , n8669 );
and ( n10972 , n671 , n8243 );
xor ( n10973 , n10971 , n10972 );
and ( n10974 , n715 , n7662 );
xor ( n10975 , n10973 , n10974 );
xor ( n10976 , n10970 , n10975 );
buf ( n10977 , n431 );
and ( n10978 , n599 , n10977 );
and ( n10979 , n608 , n10239 );
xor ( n10980 , n10978 , n10979 );
and ( n10981 , n611 , n9348 );
xor ( n10982 , n10980 , n10981 );
xor ( n10983 , n10976 , n10982 );
xor ( n10984 , n10966 , n10983 );
xor ( n10985 , n10946 , n10984 );
xor ( n10986 , n10915 , n10985 );
xor ( n10987 , n10863 , n10986 );
xor ( n10988 , n10780 , n10987 );
and ( n10989 , n10064 , n10068 );
and ( n10990 , n10068 , n10137 );
and ( n10991 , n10064 , n10137 );
or ( n10992 , n10989 , n10990 , n10991 );
and ( n10993 , n10276 , n10296 );
xor ( n10994 , n10992 , n10993 );
and ( n10995 , n10280 , n10281 );
and ( n10996 , n10281 , n10295 );
and ( n10997 , n10280 , n10295 );
or ( n10998 , n10995 , n10996 , n10997 );
and ( n10999 , n10077 , n10092 );
and ( n11000 , n10092 , n10109 );
and ( n11001 , n10077 , n10109 );
or ( n11002 , n10999 , n11000 , n11001 );
and ( n11003 , n10286 , n10294 );
xor ( n11004 , n11002 , n11003 );
and ( n11005 , n10081 , n10085 );
and ( n11006 , n10085 , n10091 );
and ( n11007 , n10081 , n10091 );
or ( n11008 , n11005 , n11006 , n11007 );
and ( n11009 , n10287 , n10293 );
xor ( n11010 , n11008 , n11009 );
and ( n11011 , n10288 , n10289 );
and ( n11012 , n10289 , n10292 );
and ( n11013 , n10288 , n10292 );
or ( n11014 , n11011 , n11012 , n11013 );
buf ( n11015 , n431 );
and ( n11016 , n11015 , n612 );
xor ( n11017 , n11014 , n11016 );
and ( n11018 , n8718 , n635 );
and ( n11019 , n9400 , n606 );
xor ( n11020 , n11018 , n11019 );
and ( n11021 , n10291 , n615 );
xor ( n11022 , n11020 , n11021 );
xor ( n11023 , n11017 , n11022 );
xor ( n11024 , n11010 , n11023 );
xor ( n11025 , n11004 , n11024 );
xor ( n11026 , n10998 , n11025 );
xor ( n11027 , n10994 , n11026 );
xor ( n11028 , n10988 , n11027 );
xor ( n11029 , n10776 , n11028 );
and ( n11030 , n10047 , n10051 );
and ( n11031 , n10051 , n10299 );
and ( n11032 , n10047 , n10299 );
or ( n11033 , n11030 , n11031 , n11032 );
xor ( n11034 , n11029 , n11033 );
and ( n11035 , n10300 , n10304 );
and ( n11036 , n10305 , n10308 );
or ( n11037 , n11035 , n11036 );
xor ( n11038 , n11034 , n11037 );
buf ( n11039 , n11038 );
buf ( n11040 , n11039 );
not ( n11041 , n11040 );
nor ( n11042 , n11041 , n8739 );
xor ( n11043 , n10767 , n11042 );
and ( n11044 , n10043 , n10313 );
and ( n11045 , n10314 , n10317 );
or ( n11046 , n11044 , n11045 );
xor ( n11047 , n11043 , n11046 );
buf ( n11048 , n11047 );
buf ( n11049 , n11048 );
not ( n11050 , n11049 );
buf ( n11051 , n538 );
not ( n11052 , n11051 );
nor ( n11053 , n11050 , n11052 );
xor ( n11054 , n10545 , n11053 );
xor ( n11055 , n10329 , n10542 );
nor ( n11056 , n10321 , n11052 );
and ( n11057 , n11055 , n11056 );
xor ( n11058 , n11055 , n11056 );
xor ( n11059 , n10333 , n10540 );
nor ( n11060 , n9429 , n11052 );
and ( n11061 , n11059 , n11060 );
xor ( n11062 , n11059 , n11060 );
xor ( n11063 , n10337 , n10538 );
nor ( n11064 , n8949 , n11052 );
and ( n11065 , n11063 , n11064 );
xor ( n11066 , n11063 , n11064 );
xor ( n11067 , n10341 , n10536 );
nor ( n11068 , n9437 , n11052 );
and ( n11069 , n11067 , n11068 );
xor ( n11070 , n11067 , n11068 );
xor ( n11071 , n10345 , n10534 );
nor ( n11072 , n9446 , n11052 );
and ( n11073 , n11071 , n11072 );
xor ( n11074 , n11071 , n11072 );
xor ( n11075 , n10349 , n10532 );
nor ( n11076 , n9455 , n11052 );
and ( n11077 , n11075 , n11076 );
xor ( n11078 , n11075 , n11076 );
xor ( n11079 , n10353 , n10530 );
nor ( n11080 , n9464 , n11052 );
and ( n11081 , n11079 , n11080 );
xor ( n11082 , n11079 , n11080 );
xor ( n11083 , n10357 , n10528 );
nor ( n11084 , n9473 , n11052 );
and ( n11085 , n11083 , n11084 );
xor ( n11086 , n11083 , n11084 );
xor ( n11087 , n10361 , n10526 );
nor ( n11088 , n9482 , n11052 );
and ( n11089 , n11087 , n11088 );
xor ( n11090 , n11087 , n11088 );
xor ( n11091 , n10365 , n10524 );
nor ( n11092 , n9491 , n11052 );
and ( n11093 , n11091 , n11092 );
xor ( n11094 , n11091 , n11092 );
xor ( n11095 , n10369 , n10522 );
nor ( n11096 , n9500 , n11052 );
and ( n11097 , n11095 , n11096 );
xor ( n11098 , n11095 , n11096 );
xor ( n11099 , n10373 , n10520 );
nor ( n11100 , n9509 , n11052 );
and ( n11101 , n11099 , n11100 );
xor ( n11102 , n11099 , n11100 );
xor ( n11103 , n10377 , n10518 );
nor ( n11104 , n9518 , n11052 );
and ( n11105 , n11103 , n11104 );
xor ( n11106 , n11103 , n11104 );
xor ( n11107 , n10381 , n10516 );
nor ( n11108 , n9527 , n11052 );
and ( n11109 , n11107 , n11108 );
xor ( n11110 , n11107 , n11108 );
xor ( n11111 , n10385 , n10514 );
nor ( n11112 , n9536 , n11052 );
and ( n11113 , n11111 , n11112 );
xor ( n11114 , n11111 , n11112 );
xor ( n11115 , n10389 , n10512 );
nor ( n11116 , n9545 , n11052 );
and ( n11117 , n11115 , n11116 );
xor ( n11118 , n11115 , n11116 );
xor ( n11119 , n10393 , n10510 );
nor ( n11120 , n9554 , n11052 );
and ( n11121 , n11119 , n11120 );
xor ( n11122 , n11119 , n11120 );
xor ( n11123 , n10397 , n10508 );
nor ( n11124 , n9563 , n11052 );
and ( n11125 , n11123 , n11124 );
xor ( n11126 , n11123 , n11124 );
xor ( n11127 , n10401 , n10506 );
nor ( n11128 , n9572 , n11052 );
and ( n11129 , n11127 , n11128 );
xor ( n11130 , n11127 , n11128 );
xor ( n11131 , n10405 , n10504 );
nor ( n11132 , n9581 , n11052 );
and ( n11133 , n11131 , n11132 );
xor ( n11134 , n11131 , n11132 );
xor ( n11135 , n10409 , n10502 );
nor ( n11136 , n9590 , n11052 );
and ( n11137 , n11135 , n11136 );
xor ( n11138 , n11135 , n11136 );
xor ( n11139 , n10413 , n10500 );
nor ( n11140 , n9599 , n11052 );
and ( n11141 , n11139 , n11140 );
xor ( n11142 , n11139 , n11140 );
xor ( n11143 , n10417 , n10498 );
nor ( n11144 , n9608 , n11052 );
and ( n11145 , n11143 , n11144 );
xor ( n11146 , n11143 , n11144 );
xor ( n11147 , n10421 , n10496 );
nor ( n11148 , n9617 , n11052 );
and ( n11149 , n11147 , n11148 );
xor ( n11150 , n11147 , n11148 );
xor ( n11151 , n10425 , n10494 );
nor ( n11152 , n9626 , n11052 );
and ( n11153 , n11151 , n11152 );
xor ( n11154 , n11151 , n11152 );
xor ( n11155 , n10429 , n10492 );
nor ( n11156 , n9635 , n11052 );
and ( n11157 , n11155 , n11156 );
xor ( n11158 , n11155 , n11156 );
xor ( n11159 , n10433 , n10490 );
nor ( n11160 , n9644 , n11052 );
and ( n11161 , n11159 , n11160 );
xor ( n11162 , n11159 , n11160 );
xor ( n11163 , n10437 , n10488 );
nor ( n11164 , n9653 , n11052 );
and ( n11165 , n11163 , n11164 );
xor ( n11166 , n11163 , n11164 );
xor ( n11167 , n10441 , n10486 );
nor ( n11168 , n9662 , n11052 );
and ( n11169 , n11167 , n11168 );
xor ( n11170 , n11167 , n11168 );
xor ( n11171 , n10445 , n10484 );
nor ( n11172 , n9671 , n11052 );
and ( n11173 , n11171 , n11172 );
xor ( n11174 , n11171 , n11172 );
xor ( n11175 , n10449 , n10482 );
nor ( n11176 , n9680 , n11052 );
and ( n11177 , n11175 , n11176 );
xor ( n11178 , n11175 , n11176 );
xor ( n11179 , n10453 , n10480 );
nor ( n11180 , n9689 , n11052 );
and ( n11181 , n11179 , n11180 );
xor ( n11182 , n11179 , n11180 );
xor ( n11183 , n10457 , n10478 );
nor ( n11184 , n9698 , n11052 );
and ( n11185 , n11183 , n11184 );
xor ( n11186 , n11183 , n11184 );
xor ( n11187 , n10461 , n10476 );
nor ( n11188 , n9707 , n11052 );
and ( n11189 , n11187 , n11188 );
xor ( n11190 , n11187 , n11188 );
xor ( n11191 , n10465 , n10474 );
nor ( n11192 , n9716 , n11052 );
and ( n11193 , n11191 , n11192 );
xor ( n11194 , n11191 , n11192 );
xor ( n11195 , n10469 , n10472 );
nor ( n11196 , n9725 , n11052 );
and ( n11197 , n11195 , n11196 );
xor ( n11198 , n11195 , n11196 );
xor ( n11199 , n10470 , n10471 );
nor ( n11200 , n9734 , n11052 );
and ( n11201 , n11199 , n11200 );
xor ( n11202 , n11199 , n11200 );
nor ( n11203 , n9752 , n10323 );
nor ( n11204 , n9743 , n11052 );
and ( n11205 , n11203 , n11204 );
and ( n11206 , n11202 , n11205 );
or ( n11207 , n11201 , n11206 );
and ( n11208 , n11198 , n11207 );
or ( n11209 , n11197 , n11208 );
and ( n11210 , n11194 , n11209 );
or ( n11211 , n11193 , n11210 );
and ( n11212 , n11190 , n11211 );
or ( n11213 , n11189 , n11212 );
and ( n11214 , n11186 , n11213 );
or ( n11215 , n11185 , n11214 );
and ( n11216 , n11182 , n11215 );
or ( n11217 , n11181 , n11216 );
and ( n11218 , n11178 , n11217 );
or ( n11219 , n11177 , n11218 );
and ( n11220 , n11174 , n11219 );
or ( n11221 , n11173 , n11220 );
and ( n11222 , n11170 , n11221 );
or ( n11223 , n11169 , n11222 );
and ( n11224 , n11166 , n11223 );
or ( n11225 , n11165 , n11224 );
and ( n11226 , n11162 , n11225 );
or ( n11227 , n11161 , n11226 );
and ( n11228 , n11158 , n11227 );
or ( n11229 , n11157 , n11228 );
and ( n11230 , n11154 , n11229 );
or ( n11231 , n11153 , n11230 );
and ( n11232 , n11150 , n11231 );
or ( n11233 , n11149 , n11232 );
and ( n11234 , n11146 , n11233 );
or ( n11235 , n11145 , n11234 );
and ( n11236 , n11142 , n11235 );
or ( n11237 , n11141 , n11236 );
and ( n11238 , n11138 , n11237 );
or ( n11239 , n11137 , n11238 );
and ( n11240 , n11134 , n11239 );
or ( n11241 , n11133 , n11240 );
and ( n11242 , n11130 , n11241 );
or ( n11243 , n11129 , n11242 );
and ( n11244 , n11126 , n11243 );
or ( n11245 , n11125 , n11244 );
and ( n11246 , n11122 , n11245 );
or ( n11247 , n11121 , n11246 );
and ( n11248 , n11118 , n11247 );
or ( n11249 , n11117 , n11248 );
and ( n11250 , n11114 , n11249 );
or ( n11251 , n11113 , n11250 );
and ( n11252 , n11110 , n11251 );
or ( n11253 , n11109 , n11252 );
and ( n11254 , n11106 , n11253 );
or ( n11255 , n11105 , n11254 );
and ( n11256 , n11102 , n11255 );
or ( n11257 , n11101 , n11256 );
and ( n11258 , n11098 , n11257 );
or ( n11259 , n11097 , n11258 );
and ( n11260 , n11094 , n11259 );
or ( n11261 , n11093 , n11260 );
and ( n11262 , n11090 , n11261 );
or ( n11263 , n11089 , n11262 );
and ( n11264 , n11086 , n11263 );
or ( n11265 , n11085 , n11264 );
and ( n11266 , n11082 , n11265 );
or ( n11267 , n11081 , n11266 );
and ( n11268 , n11078 , n11267 );
or ( n11269 , n11077 , n11268 );
and ( n11270 , n11074 , n11269 );
or ( n11271 , n11073 , n11270 );
and ( n11272 , n11070 , n11271 );
or ( n11273 , n11069 , n11272 );
and ( n11274 , n11066 , n11273 );
or ( n11275 , n11065 , n11274 );
and ( n11276 , n11062 , n11275 );
or ( n11277 , n11061 , n11276 );
and ( n11278 , n11058 , n11277 );
or ( n11279 , n11057 , n11278 );
xor ( n11280 , n11054 , n11279 );
buf ( n11281 , n494 );
not ( n11282 , n11281 );
nor ( n11283 , n601 , n11282 );
buf ( n11284 , n11283 );
nor ( n11285 , n622 , n9829 );
xor ( n11286 , n11284 , n11285 );
buf ( n11287 , n11286 );
nor ( n11288 , n646 , n8955 );
xor ( n11289 , n11287 , n11288 );
and ( n11290 , n10549 , n10550 );
buf ( n11291 , n11290 );
xor ( n11292 , n11289 , n11291 );
nor ( n11293 , n684 , n603 );
xor ( n11294 , n11292 , n11293 );
and ( n11295 , n10552 , n10553 );
and ( n11296 , n10554 , n10556 );
or ( n11297 , n11295 , n11296 );
xor ( n11298 , n11294 , n11297 );
nor ( n11299 , n733 , n652 );
xor ( n11300 , n11298 , n11299 );
and ( n11301 , n10557 , n10558 );
and ( n11302 , n10559 , n10562 );
or ( n11303 , n11301 , n11302 );
xor ( n11304 , n11300 , n11303 );
nor ( n11305 , n796 , n624 );
xor ( n11306 , n11304 , n11305 );
and ( n11307 , n10563 , n10564 );
and ( n11308 , n10565 , n10568 );
or ( n11309 , n11307 , n11308 );
xor ( n11310 , n11306 , n11309 );
nor ( n11311 , n868 , n648 );
xor ( n11312 , n11310 , n11311 );
and ( n11313 , n10569 , n10570 );
and ( n11314 , n10571 , n10574 );
or ( n11315 , n11313 , n11314 );
xor ( n11316 , n11312 , n11315 );
nor ( n11317 , n958 , n686 );
xor ( n11318 , n11316 , n11317 );
and ( n11319 , n10575 , n10576 );
and ( n11320 , n10577 , n10580 );
or ( n11321 , n11319 , n11320 );
xor ( n11322 , n11318 , n11321 );
nor ( n11323 , n1062 , n735 );
xor ( n11324 , n11322 , n11323 );
and ( n11325 , n10581 , n10582 );
and ( n11326 , n10583 , n10586 );
or ( n11327 , n11325 , n11326 );
xor ( n11328 , n11324 , n11327 );
nor ( n11329 , n1176 , n798 );
xor ( n11330 , n11328 , n11329 );
and ( n11331 , n10587 , n10588 );
and ( n11332 , n10589 , n10592 );
or ( n11333 , n11331 , n11332 );
xor ( n11334 , n11330 , n11333 );
nor ( n11335 , n1303 , n870 );
xor ( n11336 , n11334 , n11335 );
and ( n11337 , n10593 , n10594 );
and ( n11338 , n10595 , n10598 );
or ( n11339 , n11337 , n11338 );
xor ( n11340 , n11336 , n11339 );
nor ( n11341 , n1445 , n960 );
xor ( n11342 , n11340 , n11341 );
and ( n11343 , n10599 , n10600 );
and ( n11344 , n10601 , n10604 );
or ( n11345 , n11343 , n11344 );
xor ( n11346 , n11342 , n11345 );
nor ( n11347 , n1598 , n1064 );
xor ( n11348 , n11346 , n11347 );
and ( n11349 , n10605 , n10606 );
and ( n11350 , n10607 , n10610 );
or ( n11351 , n11349 , n11350 );
xor ( n11352 , n11348 , n11351 );
nor ( n11353 , n1766 , n1178 );
xor ( n11354 , n11352 , n11353 );
and ( n11355 , n10611 , n10612 );
and ( n11356 , n10613 , n10616 );
or ( n11357 , n11355 , n11356 );
xor ( n11358 , n11354 , n11357 );
nor ( n11359 , n1945 , n1305 );
xor ( n11360 , n11358 , n11359 );
and ( n11361 , n10617 , n10618 );
and ( n11362 , n10619 , n10622 );
or ( n11363 , n11361 , n11362 );
xor ( n11364 , n11360 , n11363 );
nor ( n11365 , n2137 , n1447 );
xor ( n11366 , n11364 , n11365 );
and ( n11367 , n10623 , n10624 );
and ( n11368 , n10625 , n10628 );
or ( n11369 , n11367 , n11368 );
xor ( n11370 , n11366 , n11369 );
nor ( n11371 , n2343 , n1600 );
xor ( n11372 , n11370 , n11371 );
and ( n11373 , n10629 , n10630 );
and ( n11374 , n10631 , n10634 );
or ( n11375 , n11373 , n11374 );
xor ( n11376 , n11372 , n11375 );
nor ( n11377 , n2566 , n1768 );
xor ( n11378 , n11376 , n11377 );
and ( n11379 , n10635 , n10636 );
and ( n11380 , n10637 , n10640 );
or ( n11381 , n11379 , n11380 );
xor ( n11382 , n11378 , n11381 );
nor ( n11383 , n2797 , n1947 );
xor ( n11384 , n11382 , n11383 );
and ( n11385 , n10641 , n10642 );
and ( n11386 , n10643 , n10646 );
or ( n11387 , n11385 , n11386 );
xor ( n11388 , n11384 , n11387 );
nor ( n11389 , n3043 , n2139 );
xor ( n11390 , n11388 , n11389 );
and ( n11391 , n10647 , n10648 );
and ( n11392 , n10649 , n10652 );
or ( n11393 , n11391 , n11392 );
xor ( n11394 , n11390 , n11393 );
nor ( n11395 , n3300 , n2345 );
xor ( n11396 , n11394 , n11395 );
and ( n11397 , n10653 , n10654 );
and ( n11398 , n10655 , n10658 );
or ( n11399 , n11397 , n11398 );
xor ( n11400 , n11396 , n11399 );
nor ( n11401 , n3570 , n2568 );
xor ( n11402 , n11400 , n11401 );
and ( n11403 , n10659 , n10660 );
and ( n11404 , n10661 , n10664 );
or ( n11405 , n11403 , n11404 );
xor ( n11406 , n11402 , n11405 );
nor ( n11407 , n3853 , n2799 );
xor ( n11408 , n11406 , n11407 );
and ( n11409 , n10665 , n10666 );
and ( n11410 , n10667 , n10670 );
or ( n11411 , n11409 , n11410 );
xor ( n11412 , n11408 , n11411 );
nor ( n11413 , n4151 , n3045 );
xor ( n11414 , n11412 , n11413 );
and ( n11415 , n10671 , n10672 );
and ( n11416 , n10673 , n10676 );
or ( n11417 , n11415 , n11416 );
xor ( n11418 , n11414 , n11417 );
nor ( n11419 , n4458 , n3302 );
xor ( n11420 , n11418 , n11419 );
and ( n11421 , n10677 , n10678 );
and ( n11422 , n10679 , n10682 );
or ( n11423 , n11421 , n11422 );
xor ( n11424 , n11420 , n11423 );
nor ( n11425 , n4786 , n3572 );
xor ( n11426 , n11424 , n11425 );
and ( n11427 , n10683 , n10684 );
and ( n11428 , n10685 , n10688 );
or ( n11429 , n11427 , n11428 );
xor ( n11430 , n11426 , n11429 );
nor ( n11431 , n5126 , n3855 );
xor ( n11432 , n11430 , n11431 );
and ( n11433 , n10689 , n10690 );
and ( n11434 , n10691 , n10694 );
or ( n11435 , n11433 , n11434 );
xor ( n11436 , n11432 , n11435 );
nor ( n11437 , n5477 , n4153 );
xor ( n11438 , n11436 , n11437 );
and ( n11439 , n10695 , n10696 );
and ( n11440 , n10697 , n10700 );
or ( n11441 , n11439 , n11440 );
xor ( n11442 , n11438 , n11441 );
nor ( n11443 , n5838 , n4460 );
xor ( n11444 , n11442 , n11443 );
and ( n11445 , n10701 , n10702 );
and ( n11446 , n10703 , n10706 );
or ( n11447 , n11445 , n11446 );
xor ( n11448 , n11444 , n11447 );
nor ( n11449 , n6212 , n4788 );
xor ( n11450 , n11448 , n11449 );
and ( n11451 , n10707 , n10708 );
and ( n11452 , n10709 , n10712 );
or ( n11453 , n11451 , n11452 );
xor ( n11454 , n11450 , n11453 );
nor ( n11455 , n6596 , n5128 );
xor ( n11456 , n11454 , n11455 );
and ( n11457 , n10713 , n10714 );
and ( n11458 , n10715 , n10718 );
or ( n11459 , n11457 , n11458 );
xor ( n11460 , n11456 , n11459 );
nor ( n11461 , n6997 , n5479 );
xor ( n11462 , n11460 , n11461 );
and ( n11463 , n10719 , n10720 );
and ( n11464 , n10721 , n10724 );
or ( n11465 , n11463 , n11464 );
xor ( n11466 , n11462 , n11465 );
nor ( n11467 , n7413 , n5840 );
xor ( n11468 , n11466 , n11467 );
and ( n11469 , n10725 , n10726 );
and ( n11470 , n10727 , n10730 );
or ( n11471 , n11469 , n11470 );
xor ( n11472 , n11468 , n11471 );
nor ( n11473 , n7841 , n6214 );
xor ( n11474 , n11472 , n11473 );
and ( n11475 , n10731 , n10732 );
and ( n11476 , n10733 , n10736 );
or ( n11477 , n11475 , n11476 );
xor ( n11478 , n11474 , n11477 );
nor ( n11479 , n8281 , n6598 );
xor ( n11480 , n11478 , n11479 );
and ( n11481 , n10737 , n10738 );
and ( n11482 , n10739 , n10742 );
or ( n11483 , n11481 , n11482 );
xor ( n11484 , n11480 , n11483 );
nor ( n11485 , n8737 , n6999 );
xor ( n11486 , n11484 , n11485 );
and ( n11487 , n10743 , n10744 );
and ( n11488 , n10745 , n10748 );
or ( n11489 , n11487 , n11488 );
xor ( n11490 , n11486 , n11489 );
nor ( n11491 , n9420 , n7415 );
xor ( n11492 , n11490 , n11491 );
and ( n11493 , n10749 , n10750 );
and ( n11494 , n10751 , n10754 );
or ( n11495 , n11493 , n11494 );
xor ( n11496 , n11492 , n11495 );
nor ( n11497 , n10312 , n7843 );
xor ( n11498 , n11496 , n11497 );
and ( n11499 , n10755 , n10756 );
and ( n11500 , n10757 , n10760 );
or ( n11501 , n11499 , n11500 );
xor ( n11502 , n11498 , n11501 );
nor ( n11503 , n11041 , n8283 );
xor ( n11504 , n11502 , n11503 );
and ( n11505 , n10761 , n10762 );
and ( n11506 , n10763 , n10766 );
or ( n11507 , n11505 , n11506 );
xor ( n11508 , n11504 , n11507 );
and ( n11509 , n10992 , n10993 );
and ( n11510 , n10993 , n11026 );
and ( n11511 , n10992 , n11026 );
or ( n11512 , n11509 , n11510 , n11511 );
and ( n11513 , n10780 , n10987 );
and ( n11514 , n10987 , n11027 );
and ( n11515 , n10780 , n11027 );
or ( n11516 , n11513 , n11514 , n11515 );
xor ( n11517 , n11512 , n11516 );
and ( n11518 , n10784 , n10862 );
and ( n11519 , n10862 , n10986 );
and ( n11520 , n10784 , n10986 );
or ( n11521 , n11518 , n11519 , n11520 );
and ( n11522 , n10867 , n10914 );
and ( n11523 , n10914 , n10985 );
and ( n11524 , n10867 , n10985 );
or ( n11525 , n11522 , n11523 , n11524 );
and ( n11526 , n10797 , n10834 );
and ( n11527 , n10834 , n10860 );
and ( n11528 , n10797 , n10860 );
or ( n11529 , n11526 , n11527 , n11528 );
and ( n11530 , n10871 , n10875 );
and ( n11531 , n10875 , n10913 );
and ( n11532 , n10871 , n10913 );
or ( n11533 , n11530 , n11531 , n11532 );
xor ( n11534 , n11529 , n11533 );
and ( n11535 , n10839 , n10843 );
and ( n11536 , n10843 , n10859 );
and ( n11537 , n10839 , n10859 );
or ( n11538 , n11535 , n11536 , n11537 );
and ( n11539 , n10821 , n10826 );
and ( n11540 , n10826 , n10832 );
and ( n11541 , n10821 , n10832 );
or ( n11542 , n11539 , n11540 , n11541 );
and ( n11543 , n10811 , n10812 );
and ( n11544 , n10812 , n10814 );
and ( n11545 , n10811 , n10814 );
or ( n11546 , n11543 , n11544 , n11545 );
and ( n11547 , n10822 , n10823 );
and ( n11548 , n10823 , n10825 );
and ( n11549 , n10822 , n10825 );
or ( n11550 , n11547 , n11548 , n11549 );
xor ( n11551 , n11546 , n11550 );
and ( n11552 , n7385 , n840 );
and ( n11553 , n7808 , n771 );
xor ( n11554 , n11552 , n11553 );
and ( n11555 , n8079 , n719 );
xor ( n11556 , n11554 , n11555 );
xor ( n11557 , n11551 , n11556 );
xor ( n11558 , n11542 , n11557 );
and ( n11559 , n10828 , n10829 );
and ( n11560 , n10829 , n10831 );
and ( n11561 , n10828 , n10831 );
or ( n11562 , n11559 , n11560 , n11561 );
and ( n11563 , n6187 , n1134 );
and ( n11564 , n6569 , n1034 );
xor ( n11565 , n11563 , n11564 );
and ( n11566 , n6816 , n940 );
xor ( n11567 , n11565 , n11566 );
xor ( n11568 , n11562 , n11567 );
and ( n11569 , n4959 , n1551 );
and ( n11570 , n5459 , n1424 );
xor ( n11571 , n11569 , n11570 );
and ( n11572 , n5819 , n1254 );
xor ( n11573 , n11571 , n11572 );
xor ( n11574 , n11568 , n11573 );
xor ( n11575 , n11558 , n11574 );
xor ( n11576 , n11538 , n11575 );
and ( n11577 , n10848 , n10852 );
and ( n11578 , n10852 , n10858 );
and ( n11579 , n10848 , n10858 );
or ( n11580 , n11577 , n11578 , n11579 );
and ( n11581 , n10884 , n10889 );
and ( n11582 , n10889 , n10895 );
and ( n11583 , n10884 , n10895 );
or ( n11584 , n11581 , n11582 , n11583 );
xor ( n11585 , n11580 , n11584 );
and ( n11586 , n10854 , n10855 );
and ( n11587 , n10855 , n10857 );
and ( n11588 , n10854 , n10857 );
or ( n11589 , n11586 , n11587 , n11588 );
and ( n11590 , n10885 , n10886 );
and ( n11591 , n10886 , n10888 );
and ( n11592 , n10885 , n10888 );
or ( n11593 , n11590 , n11591 , n11592 );
xor ( n11594 , n11589 , n11593 );
and ( n11595 , n4132 , n2100 );
and ( n11596 , n4438 , n1882 );
xor ( n11597 , n11595 , n11596 );
and ( n11598 , n4766 , n1738 );
xor ( n11599 , n11597 , n11598 );
xor ( n11600 , n11594 , n11599 );
xor ( n11601 , n11585 , n11600 );
xor ( n11602 , n11576 , n11601 );
xor ( n11603 , n11534 , n11602 );
xor ( n11604 , n11525 , n11603 );
and ( n11605 , n10919 , n10945 );
and ( n11606 , n10945 , n10984 );
and ( n11607 , n10919 , n10984 );
or ( n11608 , n11605 , n11606 , n11607 );
and ( n11609 , n10880 , n10896 );
and ( n11610 , n10896 , n10912 );
and ( n11611 , n10880 , n10912 );
or ( n11612 , n11609 , n11610 , n11611 );
and ( n11613 , n10923 , n10927 );
and ( n11614 , n10927 , n10944 );
and ( n11615 , n10923 , n10944 );
or ( n11616 , n11613 , n11614 , n11615 );
xor ( n11617 , n11612 , n11616 );
and ( n11618 , n10901 , n10905 );
and ( n11619 , n10905 , n10911 );
and ( n11620 , n10901 , n10911 );
or ( n11621 , n11618 , n11619 , n11620 );
and ( n11622 , n10891 , n10892 );
and ( n11623 , n10892 , n10894 );
and ( n11624 , n10891 , n10894 );
or ( n11625 , n11622 , n11623 , n11624 );
and ( n11626 , n3182 , n2739 );
and ( n11627 , n3545 , n2544 );
xor ( n11628 , n11626 , n11627 );
and ( n11629 , n3801 , n2298 );
xor ( n11630 , n11628 , n11629 );
xor ( n11631 , n11625 , n11630 );
and ( n11632 , n2462 , n3495 );
and ( n11633 , n2779 , n3271 );
xor ( n11634 , n11632 , n11633 );
buf ( n11635 , n3024 );
xor ( n11636 , n11634 , n11635 );
xor ( n11637 , n11631 , n11636 );
xor ( n11638 , n11621 , n11637 );
and ( n11639 , n10907 , n10908 );
and ( n11640 , n10908 , n10910 );
and ( n11641 , n10907 , n10910 );
or ( n11642 , n11639 , n11640 , n11641 );
and ( n11643 , n10933 , n10934 );
and ( n11644 , n10934 , n10936 );
and ( n11645 , n10933 , n10936 );
or ( n11646 , n11643 , n11644 , n11645 );
xor ( n11647 , n11642 , n11646 );
and ( n11648 , n1933 , n4403 );
and ( n11649 , n2120 , n4102 );
xor ( n11650 , n11648 , n11649 );
and ( n11651 , n2324 , n3749 );
xor ( n11652 , n11650 , n11651 );
xor ( n11653 , n11647 , n11652 );
xor ( n11654 , n11638 , n11653 );
xor ( n11655 , n11617 , n11654 );
xor ( n11656 , n11608 , n11655 );
and ( n11657 , n10950 , n10965 );
and ( n11658 , n10965 , n10983 );
and ( n11659 , n10950 , n10983 );
or ( n11660 , n11657 , n11658 , n11659 );
and ( n11661 , n10932 , n10937 );
and ( n11662 , n10937 , n10943 );
and ( n11663 , n10932 , n10943 );
or ( n11664 , n11661 , n11662 , n11663 );
and ( n11665 , n10954 , n10958 );
and ( n11666 , n10958 , n10964 );
and ( n11667 , n10954 , n10964 );
or ( n11668 , n11665 , n11666 , n11667 );
xor ( n11669 , n11664 , n11668 );
and ( n11670 , n10939 , n10940 );
and ( n11671 , n10940 , n10942 );
and ( n11672 , n10939 , n10942 );
or ( n11673 , n11670 , n11671 , n11672 );
and ( n11674 , n1383 , n5408 );
and ( n11675 , n1580 , n5103 );
xor ( n11676 , n11674 , n11675 );
and ( n11677 , n1694 , n4730 );
xor ( n11678 , n11676 , n11677 );
xor ( n11679 , n11673 , n11678 );
and ( n11680 , n1047 , n6504 );
and ( n11681 , n1164 , n6132 );
xor ( n11682 , n11680 , n11681 );
and ( n11683 , n1287 , n5765 );
xor ( n11684 , n11682 , n11683 );
xor ( n11685 , n11679 , n11684 );
xor ( n11686 , n11669 , n11685 );
xor ( n11687 , n11660 , n11686 );
and ( n11688 , n10970 , n10975 );
and ( n11689 , n10975 , n10982 );
and ( n11690 , n10970 , n10982 );
or ( n11691 , n11688 , n11689 , n11690 );
and ( n11692 , n10960 , n10961 );
and ( n11693 , n10961 , n10963 );
and ( n11694 , n10960 , n10963 );
or ( n11695 , n11692 , n11693 , n11694 );
and ( n11696 , n10971 , n10972 );
and ( n11697 , n10972 , n10974 );
and ( n11698 , n10971 , n10974 );
or ( n11699 , n11696 , n11697 , n11698 );
xor ( n11700 , n11695 , n11699 );
and ( n11701 , n783 , n7662 );
and ( n11702 , n856 , n7310 );
xor ( n11703 , n11701 , n11702 );
and ( n11704 , n925 , n6971 );
xor ( n11705 , n11703 , n11704 );
xor ( n11706 , n11700 , n11705 );
xor ( n11707 , n11691 , n11706 );
and ( n11708 , n10978 , n10979 );
and ( n11709 , n10979 , n10981 );
and ( n11710 , n10978 , n10981 );
or ( n11711 , n11708 , n11709 , n11710 );
and ( n11712 , n632 , n9348 );
and ( n11713 , n671 , n8669 );
xor ( n11714 , n11712 , n11713 );
and ( n11715 , n715 , n8243 );
xor ( n11716 , n11714 , n11715 );
xor ( n11717 , n11711 , n11716 );
buf ( n11718 , n430 );
and ( n11719 , n599 , n11718 );
and ( n11720 , n608 , n10977 );
xor ( n11721 , n11719 , n11720 );
and ( n11722 , n611 , n10239 );
xor ( n11723 , n11721 , n11722 );
xor ( n11724 , n11717 , n11723 );
xor ( n11725 , n11707 , n11724 );
xor ( n11726 , n11687 , n11725 );
xor ( n11727 , n11656 , n11726 );
xor ( n11728 , n11604 , n11727 );
xor ( n11729 , n11521 , n11728 );
and ( n11730 , n10788 , n10792 );
and ( n11731 , n10792 , n10861 );
and ( n11732 , n10788 , n10861 );
or ( n11733 , n11730 , n11731 , n11732 );
and ( n11734 , n10998 , n11025 );
xor ( n11735 , n11733 , n11734 );
and ( n11736 , n11002 , n11003 );
and ( n11737 , n11003 , n11024 );
and ( n11738 , n11002 , n11024 );
or ( n11739 , n11736 , n11737 , n11738 );
and ( n11740 , n11008 , n11009 );
and ( n11741 , n11009 , n11023 );
and ( n11742 , n11008 , n11023 );
or ( n11743 , n11740 , n11741 , n11742 );
and ( n11744 , n10801 , n10816 );
and ( n11745 , n10816 , n10833 );
and ( n11746 , n10801 , n10833 );
or ( n11747 , n11744 , n11745 , n11746 );
xor ( n11748 , n11743 , n11747 );
and ( n11749 , n11014 , n11016 );
and ( n11750 , n11016 , n11022 );
and ( n11751 , n11014 , n11022 );
or ( n11752 , n11749 , n11750 , n11751 );
and ( n11753 , n10805 , n10809 );
and ( n11754 , n10809 , n10815 );
and ( n11755 , n10805 , n10815 );
or ( n11756 , n11753 , n11754 , n11755 );
xor ( n11757 , n11752 , n11756 );
and ( n11758 , n11018 , n11019 );
and ( n11759 , n11019 , n11021 );
and ( n11760 , n11018 , n11021 );
or ( n11761 , n11758 , n11759 , n11760 );
and ( n11762 , n8718 , n663 );
and ( n11763 , n9400 , n635 );
xor ( n11764 , n11762 , n11763 );
and ( n11765 , n10291 , n606 );
xor ( n11766 , n11764 , n11765 );
xor ( n11767 , n11761 , n11766 );
and ( n11768 , n11015 , n615 );
buf ( n11769 , n430 );
and ( n11770 , n11769 , n612 );
xor ( n11771 , n11768 , n11770 );
xor ( n11772 , n11767 , n11771 );
xor ( n11773 , n11757 , n11772 );
xor ( n11774 , n11748 , n11773 );
xor ( n11775 , n11739 , n11774 );
xor ( n11776 , n11735 , n11775 );
xor ( n11777 , n11729 , n11776 );
xor ( n11778 , n11517 , n11777 );
and ( n11779 , n10771 , n10775 );
and ( n11780 , n10775 , n11028 );
and ( n11781 , n10771 , n11028 );
or ( n11782 , n11779 , n11780 , n11781 );
xor ( n11783 , n11778 , n11782 );
and ( n11784 , n11029 , n11033 );
and ( n11785 , n11034 , n11037 );
or ( n11786 , n11784 , n11785 );
xor ( n11787 , n11783 , n11786 );
buf ( n11788 , n11787 );
buf ( n11789 , n11788 );
not ( n11790 , n11789 );
nor ( n11791 , n11790 , n8739 );
xor ( n11792 , n11508 , n11791 );
and ( n11793 , n10767 , n11042 );
and ( n11794 , n11043 , n11046 );
or ( n11795 , n11793 , n11794 );
xor ( n11796 , n11792 , n11795 );
buf ( n11797 , n11796 );
buf ( n11798 , n11797 );
not ( n11799 , n11798 );
buf ( n11800 , n539 );
not ( n11801 , n11800 );
nor ( n11802 , n11799 , n11801 );
xor ( n11803 , n11280 , n11802 );
xor ( n11804 , n11058 , n11277 );
nor ( n11805 , n11050 , n11801 );
and ( n11806 , n11804 , n11805 );
xor ( n11807 , n11804 , n11805 );
xor ( n11808 , n11062 , n11275 );
nor ( n11809 , n10321 , n11801 );
and ( n11810 , n11808 , n11809 );
xor ( n11811 , n11808 , n11809 );
xor ( n11812 , n11066 , n11273 );
nor ( n11813 , n9429 , n11801 );
and ( n11814 , n11812 , n11813 );
xor ( n11815 , n11812 , n11813 );
xor ( n11816 , n11070 , n11271 );
nor ( n11817 , n8949 , n11801 );
and ( n11818 , n11816 , n11817 );
xor ( n11819 , n11816 , n11817 );
xor ( n11820 , n11074 , n11269 );
nor ( n11821 , n9437 , n11801 );
and ( n11822 , n11820 , n11821 );
xor ( n11823 , n11820 , n11821 );
xor ( n11824 , n11078 , n11267 );
nor ( n11825 , n9446 , n11801 );
and ( n11826 , n11824 , n11825 );
xor ( n11827 , n11824 , n11825 );
xor ( n11828 , n11082 , n11265 );
nor ( n11829 , n9455 , n11801 );
and ( n11830 , n11828 , n11829 );
xor ( n11831 , n11828 , n11829 );
xor ( n11832 , n11086 , n11263 );
nor ( n11833 , n9464 , n11801 );
and ( n11834 , n11832 , n11833 );
xor ( n11835 , n11832 , n11833 );
xor ( n11836 , n11090 , n11261 );
nor ( n11837 , n9473 , n11801 );
and ( n11838 , n11836 , n11837 );
xor ( n11839 , n11836 , n11837 );
xor ( n11840 , n11094 , n11259 );
nor ( n11841 , n9482 , n11801 );
and ( n11842 , n11840 , n11841 );
xor ( n11843 , n11840 , n11841 );
xor ( n11844 , n11098 , n11257 );
nor ( n11845 , n9491 , n11801 );
and ( n11846 , n11844 , n11845 );
xor ( n11847 , n11844 , n11845 );
xor ( n11848 , n11102 , n11255 );
nor ( n11849 , n9500 , n11801 );
and ( n11850 , n11848 , n11849 );
xor ( n11851 , n11848 , n11849 );
xor ( n11852 , n11106 , n11253 );
nor ( n11853 , n9509 , n11801 );
and ( n11854 , n11852 , n11853 );
xor ( n11855 , n11852 , n11853 );
xor ( n11856 , n11110 , n11251 );
nor ( n11857 , n9518 , n11801 );
and ( n11858 , n11856 , n11857 );
xor ( n11859 , n11856 , n11857 );
xor ( n11860 , n11114 , n11249 );
nor ( n11861 , n9527 , n11801 );
and ( n11862 , n11860 , n11861 );
xor ( n11863 , n11860 , n11861 );
xor ( n11864 , n11118 , n11247 );
nor ( n11865 , n9536 , n11801 );
and ( n11866 , n11864 , n11865 );
xor ( n11867 , n11864 , n11865 );
xor ( n11868 , n11122 , n11245 );
nor ( n11869 , n9545 , n11801 );
and ( n11870 , n11868 , n11869 );
xor ( n11871 , n11868 , n11869 );
xor ( n11872 , n11126 , n11243 );
nor ( n11873 , n9554 , n11801 );
and ( n11874 , n11872 , n11873 );
xor ( n11875 , n11872 , n11873 );
xor ( n11876 , n11130 , n11241 );
nor ( n11877 , n9563 , n11801 );
and ( n11878 , n11876 , n11877 );
xor ( n11879 , n11876 , n11877 );
xor ( n11880 , n11134 , n11239 );
nor ( n11881 , n9572 , n11801 );
and ( n11882 , n11880 , n11881 );
xor ( n11883 , n11880 , n11881 );
xor ( n11884 , n11138 , n11237 );
nor ( n11885 , n9581 , n11801 );
and ( n11886 , n11884 , n11885 );
xor ( n11887 , n11884 , n11885 );
xor ( n11888 , n11142 , n11235 );
nor ( n11889 , n9590 , n11801 );
and ( n11890 , n11888 , n11889 );
xor ( n11891 , n11888 , n11889 );
xor ( n11892 , n11146 , n11233 );
nor ( n11893 , n9599 , n11801 );
and ( n11894 , n11892 , n11893 );
xor ( n11895 , n11892 , n11893 );
xor ( n11896 , n11150 , n11231 );
nor ( n11897 , n9608 , n11801 );
and ( n11898 , n11896 , n11897 );
xor ( n11899 , n11896 , n11897 );
xor ( n11900 , n11154 , n11229 );
nor ( n11901 , n9617 , n11801 );
and ( n11902 , n11900 , n11901 );
xor ( n11903 , n11900 , n11901 );
xor ( n11904 , n11158 , n11227 );
nor ( n11905 , n9626 , n11801 );
and ( n11906 , n11904 , n11905 );
xor ( n11907 , n11904 , n11905 );
xor ( n11908 , n11162 , n11225 );
nor ( n11909 , n9635 , n11801 );
and ( n11910 , n11908 , n11909 );
xor ( n11911 , n11908 , n11909 );
xor ( n11912 , n11166 , n11223 );
nor ( n11913 , n9644 , n11801 );
and ( n11914 , n11912 , n11913 );
xor ( n11915 , n11912 , n11913 );
xor ( n11916 , n11170 , n11221 );
nor ( n11917 , n9653 , n11801 );
and ( n11918 , n11916 , n11917 );
xor ( n11919 , n11916 , n11917 );
xor ( n11920 , n11174 , n11219 );
nor ( n11921 , n9662 , n11801 );
and ( n11922 , n11920 , n11921 );
xor ( n11923 , n11920 , n11921 );
xor ( n11924 , n11178 , n11217 );
nor ( n11925 , n9671 , n11801 );
and ( n11926 , n11924 , n11925 );
xor ( n11927 , n11924 , n11925 );
xor ( n11928 , n11182 , n11215 );
nor ( n11929 , n9680 , n11801 );
and ( n11930 , n11928 , n11929 );
xor ( n11931 , n11928 , n11929 );
xor ( n11932 , n11186 , n11213 );
nor ( n11933 , n9689 , n11801 );
and ( n11934 , n11932 , n11933 );
xor ( n11935 , n11932 , n11933 );
xor ( n11936 , n11190 , n11211 );
nor ( n11937 , n9698 , n11801 );
and ( n11938 , n11936 , n11937 );
xor ( n11939 , n11936 , n11937 );
xor ( n11940 , n11194 , n11209 );
nor ( n11941 , n9707 , n11801 );
and ( n11942 , n11940 , n11941 );
xor ( n11943 , n11940 , n11941 );
xor ( n11944 , n11198 , n11207 );
nor ( n11945 , n9716 , n11801 );
and ( n11946 , n11944 , n11945 );
xor ( n11947 , n11944 , n11945 );
xor ( n11948 , n11202 , n11205 );
nor ( n11949 , n9725 , n11801 );
and ( n11950 , n11948 , n11949 );
xor ( n11951 , n11948 , n11949 );
xor ( n11952 , n11203 , n11204 );
nor ( n11953 , n9734 , n11801 );
and ( n11954 , n11952 , n11953 );
xor ( n11955 , n11952 , n11953 );
nor ( n11956 , n9752 , n11052 );
nor ( n11957 , n9743 , n11801 );
and ( n11958 , n11956 , n11957 );
and ( n11959 , n11955 , n11958 );
or ( n11960 , n11954 , n11959 );
and ( n11961 , n11951 , n11960 );
or ( n11962 , n11950 , n11961 );
and ( n11963 , n11947 , n11962 );
or ( n11964 , n11946 , n11963 );
and ( n11965 , n11943 , n11964 );
or ( n11966 , n11942 , n11965 );
and ( n11967 , n11939 , n11966 );
or ( n11968 , n11938 , n11967 );
and ( n11969 , n11935 , n11968 );
or ( n11970 , n11934 , n11969 );
and ( n11971 , n11931 , n11970 );
or ( n11972 , n11930 , n11971 );
and ( n11973 , n11927 , n11972 );
or ( n11974 , n11926 , n11973 );
and ( n11975 , n11923 , n11974 );
or ( n11976 , n11922 , n11975 );
and ( n11977 , n11919 , n11976 );
or ( n11978 , n11918 , n11977 );
and ( n11979 , n11915 , n11978 );
or ( n11980 , n11914 , n11979 );
and ( n11981 , n11911 , n11980 );
or ( n11982 , n11910 , n11981 );
and ( n11983 , n11907 , n11982 );
or ( n11984 , n11906 , n11983 );
and ( n11985 , n11903 , n11984 );
or ( n11986 , n11902 , n11985 );
and ( n11987 , n11899 , n11986 );
or ( n11988 , n11898 , n11987 );
and ( n11989 , n11895 , n11988 );
or ( n11990 , n11894 , n11989 );
and ( n11991 , n11891 , n11990 );
or ( n11992 , n11890 , n11991 );
and ( n11993 , n11887 , n11992 );
or ( n11994 , n11886 , n11993 );
and ( n11995 , n11883 , n11994 );
or ( n11996 , n11882 , n11995 );
and ( n11997 , n11879 , n11996 );
or ( n11998 , n11878 , n11997 );
and ( n11999 , n11875 , n11998 );
or ( n12000 , n11874 , n11999 );
and ( n12001 , n11871 , n12000 );
or ( n12002 , n11870 , n12001 );
and ( n12003 , n11867 , n12002 );
or ( n12004 , n11866 , n12003 );
and ( n12005 , n11863 , n12004 );
or ( n12006 , n11862 , n12005 );
and ( n12007 , n11859 , n12006 );
or ( n12008 , n11858 , n12007 );
and ( n12009 , n11855 , n12008 );
or ( n12010 , n11854 , n12009 );
and ( n12011 , n11851 , n12010 );
or ( n12012 , n11850 , n12011 );
and ( n12013 , n11847 , n12012 );
or ( n12014 , n11846 , n12013 );
and ( n12015 , n11843 , n12014 );
or ( n12016 , n11842 , n12015 );
and ( n12017 , n11839 , n12016 );
or ( n12018 , n11838 , n12017 );
and ( n12019 , n11835 , n12018 );
or ( n12020 , n11834 , n12019 );
and ( n12021 , n11831 , n12020 );
or ( n12022 , n11830 , n12021 );
and ( n12023 , n11827 , n12022 );
or ( n12024 , n11826 , n12023 );
and ( n12025 , n11823 , n12024 );
or ( n12026 , n11822 , n12025 );
and ( n12027 , n11819 , n12026 );
or ( n12028 , n11818 , n12027 );
and ( n12029 , n11815 , n12028 );
or ( n12030 , n11814 , n12029 );
and ( n12031 , n11811 , n12030 );
or ( n12032 , n11810 , n12031 );
and ( n12033 , n11807 , n12032 );
or ( n12034 , n11806 , n12033 );
xor ( n12035 , n11803 , n12034 );
buf ( n12036 , n493 );
not ( n12037 , n12036 );
nor ( n12038 , n601 , n12037 );
buf ( n12039 , n12038 );
nor ( n12040 , n622 , n10547 );
xor ( n12041 , n12039 , n12040 );
buf ( n12042 , n12041 );
nor ( n12043 , n646 , n9829 );
xor ( n12044 , n12042 , n12043 );
and ( n12045 , n11284 , n11285 );
buf ( n12046 , n12045 );
xor ( n12047 , n12044 , n12046 );
nor ( n12048 , n684 , n8955 );
xor ( n12049 , n12047 , n12048 );
and ( n12050 , n11287 , n11288 );
and ( n12051 , n11289 , n11291 );
or ( n12052 , n12050 , n12051 );
xor ( n12053 , n12049 , n12052 );
nor ( n12054 , n733 , n603 );
xor ( n12055 , n12053 , n12054 );
and ( n12056 , n11292 , n11293 );
and ( n12057 , n11294 , n11297 );
or ( n12058 , n12056 , n12057 );
xor ( n12059 , n12055 , n12058 );
nor ( n12060 , n796 , n652 );
xor ( n12061 , n12059 , n12060 );
and ( n12062 , n11298 , n11299 );
and ( n12063 , n11300 , n11303 );
or ( n12064 , n12062 , n12063 );
xor ( n12065 , n12061 , n12064 );
nor ( n12066 , n868 , n624 );
xor ( n12067 , n12065 , n12066 );
and ( n12068 , n11304 , n11305 );
and ( n12069 , n11306 , n11309 );
or ( n12070 , n12068 , n12069 );
xor ( n12071 , n12067 , n12070 );
nor ( n12072 , n958 , n648 );
xor ( n12073 , n12071 , n12072 );
and ( n12074 , n11310 , n11311 );
and ( n12075 , n11312 , n11315 );
or ( n12076 , n12074 , n12075 );
xor ( n12077 , n12073 , n12076 );
nor ( n12078 , n1062 , n686 );
xor ( n12079 , n12077 , n12078 );
and ( n12080 , n11316 , n11317 );
and ( n12081 , n11318 , n11321 );
or ( n12082 , n12080 , n12081 );
xor ( n12083 , n12079 , n12082 );
nor ( n12084 , n1176 , n735 );
xor ( n12085 , n12083 , n12084 );
and ( n12086 , n11322 , n11323 );
and ( n12087 , n11324 , n11327 );
or ( n12088 , n12086 , n12087 );
xor ( n12089 , n12085 , n12088 );
nor ( n12090 , n1303 , n798 );
xor ( n12091 , n12089 , n12090 );
and ( n12092 , n11328 , n11329 );
and ( n12093 , n11330 , n11333 );
or ( n12094 , n12092 , n12093 );
xor ( n12095 , n12091 , n12094 );
nor ( n12096 , n1445 , n870 );
xor ( n12097 , n12095 , n12096 );
and ( n12098 , n11334 , n11335 );
and ( n12099 , n11336 , n11339 );
or ( n12100 , n12098 , n12099 );
xor ( n12101 , n12097 , n12100 );
nor ( n12102 , n1598 , n960 );
xor ( n12103 , n12101 , n12102 );
and ( n12104 , n11340 , n11341 );
and ( n12105 , n11342 , n11345 );
or ( n12106 , n12104 , n12105 );
xor ( n12107 , n12103 , n12106 );
nor ( n12108 , n1766 , n1064 );
xor ( n12109 , n12107 , n12108 );
and ( n12110 , n11346 , n11347 );
and ( n12111 , n11348 , n11351 );
or ( n12112 , n12110 , n12111 );
xor ( n12113 , n12109 , n12112 );
nor ( n12114 , n1945 , n1178 );
xor ( n12115 , n12113 , n12114 );
and ( n12116 , n11352 , n11353 );
and ( n12117 , n11354 , n11357 );
or ( n12118 , n12116 , n12117 );
xor ( n12119 , n12115 , n12118 );
nor ( n12120 , n2137 , n1305 );
xor ( n12121 , n12119 , n12120 );
and ( n12122 , n11358 , n11359 );
and ( n12123 , n11360 , n11363 );
or ( n12124 , n12122 , n12123 );
xor ( n12125 , n12121 , n12124 );
nor ( n12126 , n2343 , n1447 );
xor ( n12127 , n12125 , n12126 );
and ( n12128 , n11364 , n11365 );
and ( n12129 , n11366 , n11369 );
or ( n12130 , n12128 , n12129 );
xor ( n12131 , n12127 , n12130 );
nor ( n12132 , n2566 , n1600 );
xor ( n12133 , n12131 , n12132 );
and ( n12134 , n11370 , n11371 );
and ( n12135 , n11372 , n11375 );
or ( n12136 , n12134 , n12135 );
xor ( n12137 , n12133 , n12136 );
nor ( n12138 , n2797 , n1768 );
xor ( n12139 , n12137 , n12138 );
and ( n12140 , n11376 , n11377 );
and ( n12141 , n11378 , n11381 );
or ( n12142 , n12140 , n12141 );
xor ( n12143 , n12139 , n12142 );
nor ( n12144 , n3043 , n1947 );
xor ( n12145 , n12143 , n12144 );
and ( n12146 , n11382 , n11383 );
and ( n12147 , n11384 , n11387 );
or ( n12148 , n12146 , n12147 );
xor ( n12149 , n12145 , n12148 );
nor ( n12150 , n3300 , n2139 );
xor ( n12151 , n12149 , n12150 );
and ( n12152 , n11388 , n11389 );
and ( n12153 , n11390 , n11393 );
or ( n12154 , n12152 , n12153 );
xor ( n12155 , n12151 , n12154 );
nor ( n12156 , n3570 , n2345 );
xor ( n12157 , n12155 , n12156 );
and ( n12158 , n11394 , n11395 );
and ( n12159 , n11396 , n11399 );
or ( n12160 , n12158 , n12159 );
xor ( n12161 , n12157 , n12160 );
nor ( n12162 , n3853 , n2568 );
xor ( n12163 , n12161 , n12162 );
and ( n12164 , n11400 , n11401 );
and ( n12165 , n11402 , n11405 );
or ( n12166 , n12164 , n12165 );
xor ( n12167 , n12163 , n12166 );
nor ( n12168 , n4151 , n2799 );
xor ( n12169 , n12167 , n12168 );
and ( n12170 , n11406 , n11407 );
and ( n12171 , n11408 , n11411 );
or ( n12172 , n12170 , n12171 );
xor ( n12173 , n12169 , n12172 );
nor ( n12174 , n4458 , n3045 );
xor ( n12175 , n12173 , n12174 );
and ( n12176 , n11412 , n11413 );
and ( n12177 , n11414 , n11417 );
or ( n12178 , n12176 , n12177 );
xor ( n12179 , n12175 , n12178 );
nor ( n12180 , n4786 , n3302 );
xor ( n12181 , n12179 , n12180 );
and ( n12182 , n11418 , n11419 );
and ( n12183 , n11420 , n11423 );
or ( n12184 , n12182 , n12183 );
xor ( n12185 , n12181 , n12184 );
nor ( n12186 , n5126 , n3572 );
xor ( n12187 , n12185 , n12186 );
and ( n12188 , n11424 , n11425 );
and ( n12189 , n11426 , n11429 );
or ( n12190 , n12188 , n12189 );
xor ( n12191 , n12187 , n12190 );
nor ( n12192 , n5477 , n3855 );
xor ( n12193 , n12191 , n12192 );
and ( n12194 , n11430 , n11431 );
and ( n12195 , n11432 , n11435 );
or ( n12196 , n12194 , n12195 );
xor ( n12197 , n12193 , n12196 );
nor ( n12198 , n5838 , n4153 );
xor ( n12199 , n12197 , n12198 );
and ( n12200 , n11436 , n11437 );
and ( n12201 , n11438 , n11441 );
or ( n12202 , n12200 , n12201 );
xor ( n12203 , n12199 , n12202 );
nor ( n12204 , n6212 , n4460 );
xor ( n12205 , n12203 , n12204 );
and ( n12206 , n11442 , n11443 );
and ( n12207 , n11444 , n11447 );
or ( n12208 , n12206 , n12207 );
xor ( n12209 , n12205 , n12208 );
nor ( n12210 , n6596 , n4788 );
xor ( n12211 , n12209 , n12210 );
and ( n12212 , n11448 , n11449 );
and ( n12213 , n11450 , n11453 );
or ( n12214 , n12212 , n12213 );
xor ( n12215 , n12211 , n12214 );
nor ( n12216 , n6997 , n5128 );
xor ( n12217 , n12215 , n12216 );
and ( n12218 , n11454 , n11455 );
and ( n12219 , n11456 , n11459 );
or ( n12220 , n12218 , n12219 );
xor ( n12221 , n12217 , n12220 );
nor ( n12222 , n7413 , n5479 );
xor ( n12223 , n12221 , n12222 );
and ( n12224 , n11460 , n11461 );
and ( n12225 , n11462 , n11465 );
or ( n12226 , n12224 , n12225 );
xor ( n12227 , n12223 , n12226 );
nor ( n12228 , n7841 , n5840 );
xor ( n12229 , n12227 , n12228 );
and ( n12230 , n11466 , n11467 );
and ( n12231 , n11468 , n11471 );
or ( n12232 , n12230 , n12231 );
xor ( n12233 , n12229 , n12232 );
nor ( n12234 , n8281 , n6214 );
xor ( n12235 , n12233 , n12234 );
and ( n12236 , n11472 , n11473 );
and ( n12237 , n11474 , n11477 );
or ( n12238 , n12236 , n12237 );
xor ( n12239 , n12235 , n12238 );
nor ( n12240 , n8737 , n6598 );
xor ( n12241 , n12239 , n12240 );
and ( n12242 , n11478 , n11479 );
and ( n12243 , n11480 , n11483 );
or ( n12244 , n12242 , n12243 );
xor ( n12245 , n12241 , n12244 );
nor ( n12246 , n9420 , n6999 );
xor ( n12247 , n12245 , n12246 );
and ( n12248 , n11484 , n11485 );
and ( n12249 , n11486 , n11489 );
or ( n12250 , n12248 , n12249 );
xor ( n12251 , n12247 , n12250 );
nor ( n12252 , n10312 , n7415 );
xor ( n12253 , n12251 , n12252 );
and ( n12254 , n11490 , n11491 );
and ( n12255 , n11492 , n11495 );
or ( n12256 , n12254 , n12255 );
xor ( n12257 , n12253 , n12256 );
nor ( n12258 , n11041 , n7843 );
xor ( n12259 , n12257 , n12258 );
and ( n12260 , n11496 , n11497 );
and ( n12261 , n11498 , n11501 );
or ( n12262 , n12260 , n12261 );
xor ( n12263 , n12259 , n12262 );
nor ( n12264 , n11790 , n8283 );
xor ( n12265 , n12263 , n12264 );
and ( n12266 , n11502 , n11503 );
and ( n12267 , n11504 , n11507 );
or ( n12268 , n12266 , n12267 );
xor ( n12269 , n12265 , n12268 );
and ( n12270 , n11733 , n11734 );
and ( n12271 , n11734 , n11775 );
and ( n12272 , n11733 , n11775 );
or ( n12273 , n12270 , n12271 , n12272 );
and ( n12274 , n11521 , n11728 );
and ( n12275 , n11728 , n11776 );
and ( n12276 , n11521 , n11776 );
or ( n12277 , n12274 , n12275 , n12276 );
xor ( n12278 , n12273 , n12277 );
and ( n12279 , n11525 , n11603 );
and ( n12280 , n11603 , n11727 );
and ( n12281 , n11525 , n11727 );
or ( n12282 , n12279 , n12280 , n12281 );
and ( n12283 , n11529 , n11533 );
and ( n12284 , n11533 , n11602 );
and ( n12285 , n11529 , n11602 );
or ( n12286 , n12283 , n12284 , n12285 );
and ( n12287 , n11739 , n11774 );
xor ( n12288 , n12286 , n12287 );
and ( n12289 , n11768 , n11770 );
and ( n12290 , n11743 , n11747 );
and ( n12291 , n11747 , n11773 );
and ( n12292 , n11743 , n11773 );
or ( n12293 , n12290 , n12291 , n12292 );
xor ( n12294 , n12289 , n12293 );
and ( n12295 , n11542 , n11557 );
and ( n12296 , n11557 , n11574 );
and ( n12297 , n11542 , n11574 );
or ( n12298 , n12295 , n12296 , n12297 );
and ( n12299 , n11752 , n11756 );
and ( n12300 , n11756 , n11772 );
and ( n12301 , n11752 , n11772 );
or ( n12302 , n12299 , n12300 , n12301 );
xor ( n12303 , n12298 , n12302 );
and ( n12304 , n11546 , n11550 );
and ( n12305 , n11550 , n11556 );
and ( n12306 , n11546 , n11556 );
or ( n12307 , n12304 , n12305 , n12306 );
and ( n12308 , n11761 , n11766 );
and ( n12309 , n11766 , n11771 );
and ( n12310 , n11761 , n11771 );
or ( n12311 , n12308 , n12309 , n12310 );
xor ( n12312 , n12307 , n12311 );
and ( n12313 , n11762 , n11763 );
and ( n12314 , n11763 , n11765 );
and ( n12315 , n11762 , n11765 );
or ( n12316 , n12313 , n12314 , n12315 );
and ( n12317 , n11015 , n606 );
and ( n12318 , n11769 , n615 );
xor ( n12319 , n12317 , n12318 );
buf ( n12320 , n429 );
and ( n12321 , n12320 , n612 );
xor ( n12322 , n12319 , n12321 );
xor ( n12323 , n12316 , n12322 );
and ( n12324 , n8718 , n719 );
and ( n12325 , n9400 , n663 );
xor ( n12326 , n12324 , n12325 );
and ( n12327 , n10291 , n635 );
xor ( n12328 , n12326 , n12327 );
xor ( n12329 , n12323 , n12328 );
xor ( n12330 , n12312 , n12329 );
xor ( n12331 , n12303 , n12330 );
xor ( n12332 , n12294 , n12331 );
xor ( n12333 , n12288 , n12332 );
xor ( n12334 , n12282 , n12333 );
and ( n12335 , n11608 , n11655 );
and ( n12336 , n11655 , n11726 );
and ( n12337 , n11608 , n11726 );
or ( n12338 , n12335 , n12336 , n12337 );
and ( n12339 , n11538 , n11575 );
and ( n12340 , n11575 , n11601 );
and ( n12341 , n11538 , n11601 );
or ( n12342 , n12339 , n12340 , n12341 );
and ( n12343 , n11612 , n11616 );
and ( n12344 , n11616 , n11654 );
and ( n12345 , n11612 , n11654 );
or ( n12346 , n12343 , n12344 , n12345 );
xor ( n12347 , n12342 , n12346 );
and ( n12348 , n11580 , n11584 );
and ( n12349 , n11584 , n11600 );
and ( n12350 , n11580 , n11600 );
or ( n12351 , n12348 , n12349 , n12350 );
and ( n12352 , n11562 , n11567 );
and ( n12353 , n11567 , n11573 );
and ( n12354 , n11562 , n11573 );
or ( n12355 , n12352 , n12353 , n12354 );
and ( n12356 , n11552 , n11553 );
and ( n12357 , n11553 , n11555 );
and ( n12358 , n11552 , n11555 );
or ( n12359 , n12356 , n12357 , n12358 );
and ( n12360 , n11563 , n11564 );
and ( n12361 , n11564 , n11566 );
and ( n12362 , n11563 , n11566 );
or ( n12363 , n12360 , n12361 , n12362 );
xor ( n12364 , n12359 , n12363 );
and ( n12365 , n7385 , n940 );
and ( n12366 , n7808 , n840 );
xor ( n12367 , n12365 , n12366 );
and ( n12368 , n8079 , n771 );
xor ( n12369 , n12367 , n12368 );
xor ( n12370 , n12364 , n12369 );
xor ( n12371 , n12355 , n12370 );
and ( n12372 , n11569 , n11570 );
and ( n12373 , n11570 , n11572 );
and ( n12374 , n11569 , n11572 );
or ( n12375 , n12372 , n12373 , n12374 );
and ( n12376 , n6187 , n1254 );
and ( n12377 , n6569 , n1134 );
xor ( n12378 , n12376 , n12377 );
and ( n12379 , n6816 , n1034 );
xor ( n12380 , n12378 , n12379 );
xor ( n12381 , n12375 , n12380 );
and ( n12382 , n4959 , n1738 );
and ( n12383 , n5459 , n1551 );
xor ( n12384 , n12382 , n12383 );
and ( n12385 , n5819 , n1424 );
xor ( n12386 , n12384 , n12385 );
xor ( n12387 , n12381 , n12386 );
xor ( n12388 , n12371 , n12387 );
xor ( n12389 , n12351 , n12388 );
and ( n12390 , n11589 , n11593 );
and ( n12391 , n11593 , n11599 );
and ( n12392 , n11589 , n11599 );
or ( n12393 , n12390 , n12391 , n12392 );
and ( n12394 , n11625 , n11630 );
and ( n12395 , n11630 , n11636 );
and ( n12396 , n11625 , n11636 );
or ( n12397 , n12394 , n12395 , n12396 );
xor ( n12398 , n12393 , n12397 );
and ( n12399 , n11595 , n11596 );
and ( n12400 , n11596 , n11598 );
and ( n12401 , n11595 , n11598 );
or ( n12402 , n12399 , n12400 , n12401 );
and ( n12403 , n11626 , n11627 );
and ( n12404 , n11627 , n11629 );
and ( n12405 , n11626 , n11629 );
or ( n12406 , n12403 , n12404 , n12405 );
xor ( n12407 , n12402 , n12406 );
and ( n12408 , n4132 , n2298 );
and ( n12409 , n4438 , n2100 );
xor ( n12410 , n12408 , n12409 );
and ( n12411 , n4766 , n1882 );
xor ( n12412 , n12410 , n12411 );
xor ( n12413 , n12407 , n12412 );
xor ( n12414 , n12398 , n12413 );
xor ( n12415 , n12389 , n12414 );
xor ( n12416 , n12347 , n12415 );
xor ( n12417 , n12338 , n12416 );
and ( n12418 , n11660 , n11686 );
and ( n12419 , n11686 , n11725 );
and ( n12420 , n11660 , n11725 );
or ( n12421 , n12418 , n12419 , n12420 );
and ( n12422 , n11621 , n11637 );
and ( n12423 , n11637 , n11653 );
and ( n12424 , n11621 , n11653 );
or ( n12425 , n12422 , n12423 , n12424 );
and ( n12426 , n11664 , n11668 );
and ( n12427 , n11668 , n11685 );
and ( n12428 , n11664 , n11685 );
or ( n12429 , n12426 , n12427 , n12428 );
xor ( n12430 , n12425 , n12429 );
and ( n12431 , n11642 , n11646 );
and ( n12432 , n11646 , n11652 );
and ( n12433 , n11642 , n11652 );
or ( n12434 , n12431 , n12432 , n12433 );
and ( n12435 , n11632 , n11633 );
and ( n12436 , n11633 , n11635 );
and ( n12437 , n11632 , n11635 );
or ( n12438 , n12435 , n12436 , n12437 );
and ( n12439 , n3182 , n2981 );
and ( n12440 , n3545 , n2739 );
xor ( n12441 , n12439 , n12440 );
and ( n12442 , n3801 , n2544 );
xor ( n12443 , n12441 , n12442 );
xor ( n12444 , n12438 , n12443 );
and ( n12445 , n2462 , n3749 );
and ( n12446 , n2779 , n3495 );
xor ( n12447 , n12445 , n12446 );
and ( n12448 , n3024 , n3271 );
xor ( n12449 , n12447 , n12448 );
xor ( n12450 , n12444 , n12449 );
xor ( n12451 , n12434 , n12450 );
and ( n12452 , n11648 , n11649 );
and ( n12453 , n11649 , n11651 );
and ( n12454 , n11648 , n11651 );
or ( n12455 , n12452 , n12453 , n12454 );
and ( n12456 , n11674 , n11675 );
and ( n12457 , n11675 , n11677 );
and ( n12458 , n11674 , n11677 );
or ( n12459 , n12456 , n12457 , n12458 );
xor ( n12460 , n12455 , n12459 );
and ( n12461 , n1933 , n4730 );
and ( n12462 , n2120 , n4403 );
xor ( n12463 , n12461 , n12462 );
and ( n12464 , n2324 , n4102 );
xor ( n12465 , n12463 , n12464 );
xor ( n12466 , n12460 , n12465 );
xor ( n12467 , n12451 , n12466 );
xor ( n12468 , n12430 , n12467 );
xor ( n12469 , n12421 , n12468 );
and ( n12470 , n11691 , n11706 );
and ( n12471 , n11706 , n11724 );
and ( n12472 , n11691 , n11724 );
or ( n12473 , n12470 , n12471 , n12472 );
and ( n12474 , n11673 , n11678 );
and ( n12475 , n11678 , n11684 );
and ( n12476 , n11673 , n11684 );
or ( n12477 , n12474 , n12475 , n12476 );
and ( n12478 , n11695 , n11699 );
and ( n12479 , n11699 , n11705 );
and ( n12480 , n11695 , n11705 );
or ( n12481 , n12478 , n12479 , n12480 );
xor ( n12482 , n12477 , n12481 );
and ( n12483 , n11680 , n11681 );
and ( n12484 , n11681 , n11683 );
and ( n12485 , n11680 , n11683 );
or ( n12486 , n12483 , n12484 , n12485 );
and ( n12487 , n1383 , n5765 );
and ( n12488 , n1580 , n5408 );
xor ( n12489 , n12487 , n12488 );
and ( n12490 , n1694 , n5103 );
xor ( n12491 , n12489 , n12490 );
xor ( n12492 , n12486 , n12491 );
and ( n12493 , n1047 , n6971 );
and ( n12494 , n1164 , n6504 );
xor ( n12495 , n12493 , n12494 );
and ( n12496 , n1287 , n6132 );
xor ( n12497 , n12495 , n12496 );
xor ( n12498 , n12492 , n12497 );
xor ( n12499 , n12482 , n12498 );
xor ( n12500 , n12473 , n12499 );
and ( n12501 , n11711 , n11716 );
and ( n12502 , n11716 , n11723 );
and ( n12503 , n11711 , n11723 );
or ( n12504 , n12501 , n12502 , n12503 );
and ( n12505 , n11701 , n11702 );
and ( n12506 , n11702 , n11704 );
and ( n12507 , n11701 , n11704 );
or ( n12508 , n12505 , n12506 , n12507 );
and ( n12509 , n11712 , n11713 );
and ( n12510 , n11713 , n11715 );
and ( n12511 , n11712 , n11715 );
or ( n12512 , n12509 , n12510 , n12511 );
xor ( n12513 , n12508 , n12512 );
and ( n12514 , n783 , n8243 );
and ( n12515 , n856 , n7662 );
xor ( n12516 , n12514 , n12515 );
and ( n12517 , n925 , n7310 );
xor ( n12518 , n12516 , n12517 );
xor ( n12519 , n12513 , n12518 );
xor ( n12520 , n12504 , n12519 );
and ( n12521 , n11719 , n11720 );
and ( n12522 , n11720 , n11722 );
and ( n12523 , n11719 , n11722 );
or ( n12524 , n12521 , n12522 , n12523 );
and ( n12525 , n632 , n10239 );
and ( n12526 , n671 , n9348 );
xor ( n12527 , n12525 , n12526 );
and ( n12528 , n715 , n8669 );
xor ( n12529 , n12527 , n12528 );
xor ( n12530 , n12524 , n12529 );
buf ( n12531 , n429 );
and ( n12532 , n599 , n12531 );
and ( n12533 , n608 , n11718 );
xor ( n12534 , n12532 , n12533 );
and ( n12535 , n611 , n10977 );
xor ( n12536 , n12534 , n12535 );
xor ( n12537 , n12530 , n12536 );
xor ( n12538 , n12520 , n12537 );
xor ( n12539 , n12500 , n12538 );
xor ( n12540 , n12469 , n12539 );
xor ( n12541 , n12417 , n12540 );
xor ( n12542 , n12334 , n12541 );
xor ( n12543 , n12278 , n12542 );
and ( n12544 , n11512 , n11516 );
and ( n12545 , n11516 , n11777 );
and ( n12546 , n11512 , n11777 );
or ( n12547 , n12544 , n12545 , n12546 );
xor ( n12548 , n12543 , n12547 );
and ( n12549 , n11778 , n11782 );
and ( n12550 , n11783 , n11786 );
or ( n12551 , n12549 , n12550 );
xor ( n12552 , n12548 , n12551 );
buf ( n12553 , n12552 );
buf ( n12554 , n12553 );
not ( n12555 , n12554 );
nor ( n12556 , n12555 , n8739 );
xor ( n12557 , n12269 , n12556 );
and ( n12558 , n11508 , n11791 );
and ( n12559 , n11792 , n11795 );
or ( n12560 , n12558 , n12559 );
xor ( n12561 , n12557 , n12560 );
buf ( n12562 , n12561 );
buf ( n12563 , n12562 );
not ( n12564 , n12563 );
buf ( n12565 , n540 );
not ( n12566 , n12565 );
nor ( n12567 , n12564 , n12566 );
xor ( n12568 , n12035 , n12567 );
xor ( n12569 , n11807 , n12032 );
nor ( n12570 , n11799 , n12566 );
and ( n12571 , n12569 , n12570 );
xor ( n12572 , n12569 , n12570 );
xor ( n12573 , n11811 , n12030 );
nor ( n12574 , n11050 , n12566 );
and ( n12575 , n12573 , n12574 );
xor ( n12576 , n12573 , n12574 );
xor ( n12577 , n11815 , n12028 );
nor ( n12578 , n10321 , n12566 );
and ( n12579 , n12577 , n12578 );
xor ( n12580 , n12577 , n12578 );
xor ( n12581 , n11819 , n12026 );
nor ( n12582 , n9429 , n12566 );
and ( n12583 , n12581 , n12582 );
xor ( n12584 , n12581 , n12582 );
xor ( n12585 , n11823 , n12024 );
nor ( n12586 , n8949 , n12566 );
and ( n12587 , n12585 , n12586 );
xor ( n12588 , n12585 , n12586 );
xor ( n12589 , n11827 , n12022 );
nor ( n12590 , n9437 , n12566 );
and ( n12591 , n12589 , n12590 );
xor ( n12592 , n12589 , n12590 );
xor ( n12593 , n11831 , n12020 );
nor ( n12594 , n9446 , n12566 );
and ( n12595 , n12593 , n12594 );
xor ( n12596 , n12593 , n12594 );
xor ( n12597 , n11835 , n12018 );
nor ( n12598 , n9455 , n12566 );
and ( n12599 , n12597 , n12598 );
xor ( n12600 , n12597 , n12598 );
xor ( n12601 , n11839 , n12016 );
nor ( n12602 , n9464 , n12566 );
and ( n12603 , n12601 , n12602 );
xor ( n12604 , n12601 , n12602 );
xor ( n12605 , n11843 , n12014 );
nor ( n12606 , n9473 , n12566 );
and ( n12607 , n12605 , n12606 );
xor ( n12608 , n12605 , n12606 );
xor ( n12609 , n11847 , n12012 );
nor ( n12610 , n9482 , n12566 );
and ( n12611 , n12609 , n12610 );
xor ( n12612 , n12609 , n12610 );
xor ( n12613 , n11851 , n12010 );
nor ( n12614 , n9491 , n12566 );
and ( n12615 , n12613 , n12614 );
xor ( n12616 , n12613 , n12614 );
xor ( n12617 , n11855 , n12008 );
nor ( n12618 , n9500 , n12566 );
and ( n12619 , n12617 , n12618 );
xor ( n12620 , n12617 , n12618 );
xor ( n12621 , n11859 , n12006 );
nor ( n12622 , n9509 , n12566 );
and ( n12623 , n12621 , n12622 );
xor ( n12624 , n12621 , n12622 );
xor ( n12625 , n11863 , n12004 );
nor ( n12626 , n9518 , n12566 );
and ( n12627 , n12625 , n12626 );
xor ( n12628 , n12625 , n12626 );
xor ( n12629 , n11867 , n12002 );
nor ( n12630 , n9527 , n12566 );
and ( n12631 , n12629 , n12630 );
xor ( n12632 , n12629 , n12630 );
xor ( n12633 , n11871 , n12000 );
nor ( n12634 , n9536 , n12566 );
and ( n12635 , n12633 , n12634 );
xor ( n12636 , n12633 , n12634 );
xor ( n12637 , n11875 , n11998 );
nor ( n12638 , n9545 , n12566 );
and ( n12639 , n12637 , n12638 );
xor ( n12640 , n12637 , n12638 );
xor ( n12641 , n11879 , n11996 );
nor ( n12642 , n9554 , n12566 );
and ( n12643 , n12641 , n12642 );
xor ( n12644 , n12641 , n12642 );
xor ( n12645 , n11883 , n11994 );
nor ( n12646 , n9563 , n12566 );
and ( n12647 , n12645 , n12646 );
xor ( n12648 , n12645 , n12646 );
xor ( n12649 , n11887 , n11992 );
nor ( n12650 , n9572 , n12566 );
and ( n12651 , n12649 , n12650 );
xor ( n12652 , n12649 , n12650 );
xor ( n12653 , n11891 , n11990 );
nor ( n12654 , n9581 , n12566 );
and ( n12655 , n12653 , n12654 );
xor ( n12656 , n12653 , n12654 );
xor ( n12657 , n11895 , n11988 );
nor ( n12658 , n9590 , n12566 );
and ( n12659 , n12657 , n12658 );
xor ( n12660 , n12657 , n12658 );
xor ( n12661 , n11899 , n11986 );
nor ( n12662 , n9599 , n12566 );
and ( n12663 , n12661 , n12662 );
xor ( n12664 , n12661 , n12662 );
xor ( n12665 , n11903 , n11984 );
nor ( n12666 , n9608 , n12566 );
and ( n12667 , n12665 , n12666 );
xor ( n12668 , n12665 , n12666 );
xor ( n12669 , n11907 , n11982 );
nor ( n12670 , n9617 , n12566 );
and ( n12671 , n12669 , n12670 );
xor ( n12672 , n12669 , n12670 );
xor ( n12673 , n11911 , n11980 );
nor ( n12674 , n9626 , n12566 );
and ( n12675 , n12673 , n12674 );
xor ( n12676 , n12673 , n12674 );
xor ( n12677 , n11915 , n11978 );
nor ( n12678 , n9635 , n12566 );
and ( n12679 , n12677 , n12678 );
xor ( n12680 , n12677 , n12678 );
xor ( n12681 , n11919 , n11976 );
nor ( n12682 , n9644 , n12566 );
and ( n12683 , n12681 , n12682 );
xor ( n12684 , n12681 , n12682 );
xor ( n12685 , n11923 , n11974 );
nor ( n12686 , n9653 , n12566 );
and ( n12687 , n12685 , n12686 );
xor ( n12688 , n12685 , n12686 );
xor ( n12689 , n11927 , n11972 );
nor ( n12690 , n9662 , n12566 );
and ( n12691 , n12689 , n12690 );
xor ( n12692 , n12689 , n12690 );
xor ( n12693 , n11931 , n11970 );
nor ( n12694 , n9671 , n12566 );
and ( n12695 , n12693 , n12694 );
xor ( n12696 , n12693 , n12694 );
xor ( n12697 , n11935 , n11968 );
nor ( n12698 , n9680 , n12566 );
and ( n12699 , n12697 , n12698 );
xor ( n12700 , n12697 , n12698 );
xor ( n12701 , n11939 , n11966 );
nor ( n12702 , n9689 , n12566 );
and ( n12703 , n12701 , n12702 );
xor ( n12704 , n12701 , n12702 );
xor ( n12705 , n11943 , n11964 );
nor ( n12706 , n9698 , n12566 );
and ( n12707 , n12705 , n12706 );
xor ( n12708 , n12705 , n12706 );
xor ( n12709 , n11947 , n11962 );
nor ( n12710 , n9707 , n12566 );
and ( n12711 , n12709 , n12710 );
xor ( n12712 , n12709 , n12710 );
xor ( n12713 , n11951 , n11960 );
nor ( n12714 , n9716 , n12566 );
and ( n12715 , n12713 , n12714 );
xor ( n12716 , n12713 , n12714 );
xor ( n12717 , n11955 , n11958 );
nor ( n12718 , n9725 , n12566 );
and ( n12719 , n12717 , n12718 );
xor ( n12720 , n12717 , n12718 );
xor ( n12721 , n11956 , n11957 );
nor ( n12722 , n9734 , n12566 );
and ( n12723 , n12721 , n12722 );
xor ( n12724 , n12721 , n12722 );
nor ( n12725 , n9752 , n11801 );
nor ( n12726 , n9743 , n12566 );
and ( n12727 , n12725 , n12726 );
and ( n12728 , n12724 , n12727 );
or ( n12729 , n12723 , n12728 );
and ( n12730 , n12720 , n12729 );
or ( n12731 , n12719 , n12730 );
and ( n12732 , n12716 , n12731 );
or ( n12733 , n12715 , n12732 );
and ( n12734 , n12712 , n12733 );
or ( n12735 , n12711 , n12734 );
and ( n12736 , n12708 , n12735 );
or ( n12737 , n12707 , n12736 );
and ( n12738 , n12704 , n12737 );
or ( n12739 , n12703 , n12738 );
and ( n12740 , n12700 , n12739 );
or ( n12741 , n12699 , n12740 );
and ( n12742 , n12696 , n12741 );
or ( n12743 , n12695 , n12742 );
and ( n12744 , n12692 , n12743 );
or ( n12745 , n12691 , n12744 );
and ( n12746 , n12688 , n12745 );
or ( n12747 , n12687 , n12746 );
and ( n12748 , n12684 , n12747 );
or ( n12749 , n12683 , n12748 );
and ( n12750 , n12680 , n12749 );
or ( n12751 , n12679 , n12750 );
and ( n12752 , n12676 , n12751 );
or ( n12753 , n12675 , n12752 );
and ( n12754 , n12672 , n12753 );
or ( n12755 , n12671 , n12754 );
and ( n12756 , n12668 , n12755 );
or ( n12757 , n12667 , n12756 );
and ( n12758 , n12664 , n12757 );
or ( n12759 , n12663 , n12758 );
and ( n12760 , n12660 , n12759 );
or ( n12761 , n12659 , n12760 );
and ( n12762 , n12656 , n12761 );
or ( n12763 , n12655 , n12762 );
and ( n12764 , n12652 , n12763 );
or ( n12765 , n12651 , n12764 );
and ( n12766 , n12648 , n12765 );
or ( n12767 , n12647 , n12766 );
and ( n12768 , n12644 , n12767 );
or ( n12769 , n12643 , n12768 );
and ( n12770 , n12640 , n12769 );
or ( n12771 , n12639 , n12770 );
and ( n12772 , n12636 , n12771 );
or ( n12773 , n12635 , n12772 );
and ( n12774 , n12632 , n12773 );
or ( n12775 , n12631 , n12774 );
and ( n12776 , n12628 , n12775 );
or ( n12777 , n12627 , n12776 );
and ( n12778 , n12624 , n12777 );
or ( n12779 , n12623 , n12778 );
and ( n12780 , n12620 , n12779 );
or ( n12781 , n12619 , n12780 );
and ( n12782 , n12616 , n12781 );
or ( n12783 , n12615 , n12782 );
and ( n12784 , n12612 , n12783 );
or ( n12785 , n12611 , n12784 );
and ( n12786 , n12608 , n12785 );
or ( n12787 , n12607 , n12786 );
and ( n12788 , n12604 , n12787 );
or ( n12789 , n12603 , n12788 );
and ( n12790 , n12600 , n12789 );
or ( n12791 , n12599 , n12790 );
and ( n12792 , n12596 , n12791 );
or ( n12793 , n12595 , n12792 );
and ( n12794 , n12592 , n12793 );
or ( n12795 , n12591 , n12794 );
and ( n12796 , n12588 , n12795 );
or ( n12797 , n12587 , n12796 );
and ( n12798 , n12584 , n12797 );
or ( n12799 , n12583 , n12798 );
and ( n12800 , n12580 , n12799 );
or ( n12801 , n12579 , n12800 );
and ( n12802 , n12576 , n12801 );
or ( n12803 , n12575 , n12802 );
and ( n12804 , n12572 , n12803 );
or ( n12805 , n12571 , n12804 );
xor ( n12806 , n12568 , n12805 );
buf ( n12807 , n492 );
not ( n12808 , n12807 );
nor ( n12809 , n601 , n12808 );
buf ( n12810 , n12809 );
nor ( n12811 , n622 , n11282 );
xor ( n12812 , n12810 , n12811 );
buf ( n12813 , n12812 );
nor ( n12814 , n646 , n10547 );
xor ( n12815 , n12813 , n12814 );
and ( n12816 , n12039 , n12040 );
buf ( n12817 , n12816 );
xor ( n12818 , n12815 , n12817 );
nor ( n12819 , n684 , n9829 );
xor ( n12820 , n12818 , n12819 );
and ( n12821 , n12042 , n12043 );
and ( n12822 , n12044 , n12046 );
or ( n12823 , n12821 , n12822 );
xor ( n12824 , n12820 , n12823 );
nor ( n12825 , n733 , n8955 );
xor ( n12826 , n12824 , n12825 );
and ( n12827 , n12047 , n12048 );
and ( n12828 , n12049 , n12052 );
or ( n12829 , n12827 , n12828 );
xor ( n12830 , n12826 , n12829 );
nor ( n12831 , n796 , n603 );
xor ( n12832 , n12830 , n12831 );
and ( n12833 , n12053 , n12054 );
and ( n12834 , n12055 , n12058 );
or ( n12835 , n12833 , n12834 );
xor ( n12836 , n12832 , n12835 );
nor ( n12837 , n868 , n652 );
xor ( n12838 , n12836 , n12837 );
and ( n12839 , n12059 , n12060 );
and ( n12840 , n12061 , n12064 );
or ( n12841 , n12839 , n12840 );
xor ( n12842 , n12838 , n12841 );
nor ( n12843 , n958 , n624 );
xor ( n12844 , n12842 , n12843 );
and ( n12845 , n12065 , n12066 );
and ( n12846 , n12067 , n12070 );
or ( n12847 , n12845 , n12846 );
xor ( n12848 , n12844 , n12847 );
nor ( n12849 , n1062 , n648 );
xor ( n12850 , n12848 , n12849 );
and ( n12851 , n12071 , n12072 );
and ( n12852 , n12073 , n12076 );
or ( n12853 , n12851 , n12852 );
xor ( n12854 , n12850 , n12853 );
nor ( n12855 , n1176 , n686 );
xor ( n12856 , n12854 , n12855 );
and ( n12857 , n12077 , n12078 );
and ( n12858 , n12079 , n12082 );
or ( n12859 , n12857 , n12858 );
xor ( n12860 , n12856 , n12859 );
nor ( n12861 , n1303 , n735 );
xor ( n12862 , n12860 , n12861 );
and ( n12863 , n12083 , n12084 );
and ( n12864 , n12085 , n12088 );
or ( n12865 , n12863 , n12864 );
xor ( n12866 , n12862 , n12865 );
nor ( n12867 , n1445 , n798 );
xor ( n12868 , n12866 , n12867 );
and ( n12869 , n12089 , n12090 );
and ( n12870 , n12091 , n12094 );
or ( n12871 , n12869 , n12870 );
xor ( n12872 , n12868 , n12871 );
nor ( n12873 , n1598 , n870 );
xor ( n12874 , n12872 , n12873 );
and ( n12875 , n12095 , n12096 );
and ( n12876 , n12097 , n12100 );
or ( n12877 , n12875 , n12876 );
xor ( n12878 , n12874 , n12877 );
nor ( n12879 , n1766 , n960 );
xor ( n12880 , n12878 , n12879 );
and ( n12881 , n12101 , n12102 );
and ( n12882 , n12103 , n12106 );
or ( n12883 , n12881 , n12882 );
xor ( n12884 , n12880 , n12883 );
nor ( n12885 , n1945 , n1064 );
xor ( n12886 , n12884 , n12885 );
and ( n12887 , n12107 , n12108 );
and ( n12888 , n12109 , n12112 );
or ( n12889 , n12887 , n12888 );
xor ( n12890 , n12886 , n12889 );
nor ( n12891 , n2137 , n1178 );
xor ( n12892 , n12890 , n12891 );
and ( n12893 , n12113 , n12114 );
and ( n12894 , n12115 , n12118 );
or ( n12895 , n12893 , n12894 );
xor ( n12896 , n12892 , n12895 );
nor ( n12897 , n2343 , n1305 );
xor ( n12898 , n12896 , n12897 );
and ( n12899 , n12119 , n12120 );
and ( n12900 , n12121 , n12124 );
or ( n12901 , n12899 , n12900 );
xor ( n12902 , n12898 , n12901 );
nor ( n12903 , n2566 , n1447 );
xor ( n12904 , n12902 , n12903 );
and ( n12905 , n12125 , n12126 );
and ( n12906 , n12127 , n12130 );
or ( n12907 , n12905 , n12906 );
xor ( n12908 , n12904 , n12907 );
nor ( n12909 , n2797 , n1600 );
xor ( n12910 , n12908 , n12909 );
and ( n12911 , n12131 , n12132 );
and ( n12912 , n12133 , n12136 );
or ( n12913 , n12911 , n12912 );
xor ( n12914 , n12910 , n12913 );
nor ( n12915 , n3043 , n1768 );
xor ( n12916 , n12914 , n12915 );
and ( n12917 , n12137 , n12138 );
and ( n12918 , n12139 , n12142 );
or ( n12919 , n12917 , n12918 );
xor ( n12920 , n12916 , n12919 );
nor ( n12921 , n3300 , n1947 );
xor ( n12922 , n12920 , n12921 );
and ( n12923 , n12143 , n12144 );
and ( n12924 , n12145 , n12148 );
or ( n12925 , n12923 , n12924 );
xor ( n12926 , n12922 , n12925 );
nor ( n12927 , n3570 , n2139 );
xor ( n12928 , n12926 , n12927 );
and ( n12929 , n12149 , n12150 );
and ( n12930 , n12151 , n12154 );
or ( n12931 , n12929 , n12930 );
xor ( n12932 , n12928 , n12931 );
nor ( n12933 , n3853 , n2345 );
xor ( n12934 , n12932 , n12933 );
and ( n12935 , n12155 , n12156 );
and ( n12936 , n12157 , n12160 );
or ( n12937 , n12935 , n12936 );
xor ( n12938 , n12934 , n12937 );
nor ( n12939 , n4151 , n2568 );
xor ( n12940 , n12938 , n12939 );
and ( n12941 , n12161 , n12162 );
and ( n12942 , n12163 , n12166 );
or ( n12943 , n12941 , n12942 );
xor ( n12944 , n12940 , n12943 );
nor ( n12945 , n4458 , n2799 );
xor ( n12946 , n12944 , n12945 );
and ( n12947 , n12167 , n12168 );
and ( n12948 , n12169 , n12172 );
or ( n12949 , n12947 , n12948 );
xor ( n12950 , n12946 , n12949 );
nor ( n12951 , n4786 , n3045 );
xor ( n12952 , n12950 , n12951 );
and ( n12953 , n12173 , n12174 );
and ( n12954 , n12175 , n12178 );
or ( n12955 , n12953 , n12954 );
xor ( n12956 , n12952 , n12955 );
nor ( n12957 , n5126 , n3302 );
xor ( n12958 , n12956 , n12957 );
and ( n12959 , n12179 , n12180 );
and ( n12960 , n12181 , n12184 );
or ( n12961 , n12959 , n12960 );
xor ( n12962 , n12958 , n12961 );
nor ( n12963 , n5477 , n3572 );
xor ( n12964 , n12962 , n12963 );
and ( n12965 , n12185 , n12186 );
and ( n12966 , n12187 , n12190 );
or ( n12967 , n12965 , n12966 );
xor ( n12968 , n12964 , n12967 );
nor ( n12969 , n5838 , n3855 );
xor ( n12970 , n12968 , n12969 );
and ( n12971 , n12191 , n12192 );
and ( n12972 , n12193 , n12196 );
or ( n12973 , n12971 , n12972 );
xor ( n12974 , n12970 , n12973 );
nor ( n12975 , n6212 , n4153 );
xor ( n12976 , n12974 , n12975 );
and ( n12977 , n12197 , n12198 );
and ( n12978 , n12199 , n12202 );
or ( n12979 , n12977 , n12978 );
xor ( n12980 , n12976 , n12979 );
nor ( n12981 , n6596 , n4460 );
xor ( n12982 , n12980 , n12981 );
and ( n12983 , n12203 , n12204 );
and ( n12984 , n12205 , n12208 );
or ( n12985 , n12983 , n12984 );
xor ( n12986 , n12982 , n12985 );
nor ( n12987 , n6997 , n4788 );
xor ( n12988 , n12986 , n12987 );
and ( n12989 , n12209 , n12210 );
and ( n12990 , n12211 , n12214 );
or ( n12991 , n12989 , n12990 );
xor ( n12992 , n12988 , n12991 );
nor ( n12993 , n7413 , n5128 );
xor ( n12994 , n12992 , n12993 );
and ( n12995 , n12215 , n12216 );
and ( n12996 , n12217 , n12220 );
or ( n12997 , n12995 , n12996 );
xor ( n12998 , n12994 , n12997 );
nor ( n12999 , n7841 , n5479 );
xor ( n13000 , n12998 , n12999 );
and ( n13001 , n12221 , n12222 );
and ( n13002 , n12223 , n12226 );
or ( n13003 , n13001 , n13002 );
xor ( n13004 , n13000 , n13003 );
nor ( n13005 , n8281 , n5840 );
xor ( n13006 , n13004 , n13005 );
and ( n13007 , n12227 , n12228 );
and ( n13008 , n12229 , n12232 );
or ( n13009 , n13007 , n13008 );
xor ( n13010 , n13006 , n13009 );
nor ( n13011 , n8737 , n6214 );
xor ( n13012 , n13010 , n13011 );
and ( n13013 , n12233 , n12234 );
and ( n13014 , n12235 , n12238 );
or ( n13015 , n13013 , n13014 );
xor ( n13016 , n13012 , n13015 );
nor ( n13017 , n9420 , n6598 );
xor ( n13018 , n13016 , n13017 );
and ( n13019 , n12239 , n12240 );
and ( n13020 , n12241 , n12244 );
or ( n13021 , n13019 , n13020 );
xor ( n13022 , n13018 , n13021 );
nor ( n13023 , n10312 , n6999 );
xor ( n13024 , n13022 , n13023 );
and ( n13025 , n12245 , n12246 );
and ( n13026 , n12247 , n12250 );
or ( n13027 , n13025 , n13026 );
xor ( n13028 , n13024 , n13027 );
nor ( n13029 , n11041 , n7415 );
xor ( n13030 , n13028 , n13029 );
and ( n13031 , n12251 , n12252 );
and ( n13032 , n12253 , n12256 );
or ( n13033 , n13031 , n13032 );
xor ( n13034 , n13030 , n13033 );
nor ( n13035 , n11790 , n7843 );
xor ( n13036 , n13034 , n13035 );
and ( n13037 , n12257 , n12258 );
and ( n13038 , n12259 , n12262 );
or ( n13039 , n13037 , n13038 );
xor ( n13040 , n13036 , n13039 );
nor ( n13041 , n12555 , n8283 );
xor ( n13042 , n13040 , n13041 );
and ( n13043 , n12263 , n12264 );
and ( n13044 , n12265 , n12268 );
or ( n13045 , n13043 , n13044 );
xor ( n13046 , n13042 , n13045 );
and ( n13047 , n12286 , n12287 );
and ( n13048 , n12287 , n12332 );
and ( n13049 , n12286 , n12332 );
or ( n13050 , n13047 , n13048 , n13049 );
and ( n13051 , n12282 , n12333 );
and ( n13052 , n12333 , n12541 );
and ( n13053 , n12282 , n12541 );
or ( n13054 , n13051 , n13052 , n13053 );
xor ( n13055 , n13050 , n13054 );
and ( n13056 , n12338 , n12416 );
and ( n13057 , n12416 , n12540 );
and ( n13058 , n12338 , n12540 );
or ( n13059 , n13056 , n13057 , n13058 );
and ( n13060 , n12421 , n12468 );
and ( n13061 , n12468 , n12539 );
and ( n13062 , n12421 , n12539 );
or ( n13063 , n13060 , n13061 , n13062 );
and ( n13064 , n12351 , n12388 );
and ( n13065 , n12388 , n12414 );
and ( n13066 , n12351 , n12414 );
or ( n13067 , n13064 , n13065 , n13066 );
and ( n13068 , n12425 , n12429 );
and ( n13069 , n12429 , n12467 );
and ( n13070 , n12425 , n12467 );
or ( n13071 , n13068 , n13069 , n13070 );
xor ( n13072 , n13067 , n13071 );
and ( n13073 , n12393 , n12397 );
and ( n13074 , n12397 , n12413 );
and ( n13075 , n12393 , n12413 );
or ( n13076 , n13073 , n13074 , n13075 );
and ( n13077 , n12375 , n12380 );
and ( n13078 , n12380 , n12386 );
and ( n13079 , n12375 , n12386 );
or ( n13080 , n13077 , n13078 , n13079 );
and ( n13081 , n12365 , n12366 );
and ( n13082 , n12366 , n12368 );
and ( n13083 , n12365 , n12368 );
or ( n13084 , n13081 , n13082 , n13083 );
and ( n13085 , n12376 , n12377 );
and ( n13086 , n12377 , n12379 );
and ( n13087 , n12376 , n12379 );
or ( n13088 , n13085 , n13086 , n13087 );
xor ( n13089 , n13084 , n13088 );
and ( n13090 , n7385 , n1034 );
and ( n13091 , n7808 , n940 );
xor ( n13092 , n13090 , n13091 );
and ( n13093 , n8079 , n840 );
xor ( n13094 , n13092 , n13093 );
xor ( n13095 , n13089 , n13094 );
xor ( n13096 , n13080 , n13095 );
and ( n13097 , n12382 , n12383 );
and ( n13098 , n12383 , n12385 );
and ( n13099 , n12382 , n12385 );
or ( n13100 , n13097 , n13098 , n13099 );
and ( n13101 , n6187 , n1424 );
and ( n13102 , n6569 , n1254 );
xor ( n13103 , n13101 , n13102 );
and ( n13104 , n6816 , n1134 );
xor ( n13105 , n13103 , n13104 );
xor ( n13106 , n13100 , n13105 );
and ( n13107 , n4959 , n1882 );
and ( n13108 , n5459 , n1738 );
xor ( n13109 , n13107 , n13108 );
and ( n13110 , n5819 , n1551 );
xor ( n13111 , n13109 , n13110 );
xor ( n13112 , n13106 , n13111 );
xor ( n13113 , n13096 , n13112 );
xor ( n13114 , n13076 , n13113 );
and ( n13115 , n12402 , n12406 );
and ( n13116 , n12406 , n12412 );
and ( n13117 , n12402 , n12412 );
or ( n13118 , n13115 , n13116 , n13117 );
and ( n13119 , n12438 , n12443 );
and ( n13120 , n12443 , n12449 );
and ( n13121 , n12438 , n12449 );
or ( n13122 , n13119 , n13120 , n13121 );
xor ( n13123 , n13118 , n13122 );
and ( n13124 , n12408 , n12409 );
and ( n13125 , n12409 , n12411 );
and ( n13126 , n12408 , n12411 );
or ( n13127 , n13124 , n13125 , n13126 );
and ( n13128 , n12439 , n12440 );
and ( n13129 , n12440 , n12442 );
and ( n13130 , n12439 , n12442 );
or ( n13131 , n13128 , n13129 , n13130 );
xor ( n13132 , n13127 , n13131 );
and ( n13133 , n4132 , n2544 );
and ( n13134 , n4438 , n2298 );
xor ( n13135 , n13133 , n13134 );
and ( n13136 , n4766 , n2100 );
xor ( n13137 , n13135 , n13136 );
xor ( n13138 , n13132 , n13137 );
xor ( n13139 , n13123 , n13138 );
xor ( n13140 , n13114 , n13139 );
xor ( n13141 , n13072 , n13140 );
xor ( n13142 , n13063 , n13141 );
and ( n13143 , n12473 , n12499 );
and ( n13144 , n12499 , n12538 );
and ( n13145 , n12473 , n12538 );
or ( n13146 , n13143 , n13144 , n13145 );
and ( n13147 , n12434 , n12450 );
and ( n13148 , n12450 , n12466 );
and ( n13149 , n12434 , n12466 );
or ( n13150 , n13147 , n13148 , n13149 );
and ( n13151 , n12477 , n12481 );
and ( n13152 , n12481 , n12498 );
and ( n13153 , n12477 , n12498 );
or ( n13154 , n13151 , n13152 , n13153 );
xor ( n13155 , n13150 , n13154 );
and ( n13156 , n12455 , n12459 );
and ( n13157 , n12459 , n12465 );
and ( n13158 , n12455 , n12465 );
or ( n13159 , n13156 , n13157 , n13158 );
and ( n13160 , n12445 , n12446 );
and ( n13161 , n12446 , n12448 );
and ( n13162 , n12445 , n12448 );
or ( n13163 , n13160 , n13161 , n13162 );
buf ( n13164 , n3182 );
and ( n13165 , n3545 , n2981 );
xor ( n13166 , n13164 , n13165 );
and ( n13167 , n3801 , n2739 );
xor ( n13168 , n13166 , n13167 );
xor ( n13169 , n13163 , n13168 );
and ( n13170 , n2462 , n4102 );
and ( n13171 , n2779 , n3749 );
xor ( n13172 , n13170 , n13171 );
and ( n13173 , n3024 , n3495 );
xor ( n13174 , n13172 , n13173 );
xor ( n13175 , n13169 , n13174 );
xor ( n13176 , n13159 , n13175 );
and ( n13177 , n12461 , n12462 );
and ( n13178 , n12462 , n12464 );
and ( n13179 , n12461 , n12464 );
or ( n13180 , n13177 , n13178 , n13179 );
and ( n13181 , n12487 , n12488 );
and ( n13182 , n12488 , n12490 );
and ( n13183 , n12487 , n12490 );
or ( n13184 , n13181 , n13182 , n13183 );
xor ( n13185 , n13180 , n13184 );
and ( n13186 , n1933 , n5103 );
and ( n13187 , n2120 , n4730 );
xor ( n13188 , n13186 , n13187 );
and ( n13189 , n2324 , n4403 );
xor ( n13190 , n13188 , n13189 );
xor ( n13191 , n13185 , n13190 );
xor ( n13192 , n13176 , n13191 );
xor ( n13193 , n13155 , n13192 );
xor ( n13194 , n13146 , n13193 );
and ( n13195 , n12504 , n12519 );
and ( n13196 , n12519 , n12537 );
and ( n13197 , n12504 , n12537 );
or ( n13198 , n13195 , n13196 , n13197 );
and ( n13199 , n12486 , n12491 );
and ( n13200 , n12491 , n12497 );
and ( n13201 , n12486 , n12497 );
or ( n13202 , n13199 , n13200 , n13201 );
and ( n13203 , n12508 , n12512 );
and ( n13204 , n12512 , n12518 );
and ( n13205 , n12508 , n12518 );
or ( n13206 , n13203 , n13204 , n13205 );
xor ( n13207 , n13202 , n13206 );
and ( n13208 , n12493 , n12494 );
and ( n13209 , n12494 , n12496 );
and ( n13210 , n12493 , n12496 );
or ( n13211 , n13208 , n13209 , n13210 );
and ( n13212 , n1383 , n6132 );
and ( n13213 , n1580 , n5765 );
xor ( n13214 , n13212 , n13213 );
and ( n13215 , n1694 , n5408 );
xor ( n13216 , n13214 , n13215 );
xor ( n13217 , n13211 , n13216 );
and ( n13218 , n1047 , n7310 );
and ( n13219 , n1164 , n6971 );
xor ( n13220 , n13218 , n13219 );
and ( n13221 , n1287 , n6504 );
xor ( n13222 , n13220 , n13221 );
xor ( n13223 , n13217 , n13222 );
xor ( n13224 , n13207 , n13223 );
xor ( n13225 , n13198 , n13224 );
and ( n13226 , n12524 , n12529 );
and ( n13227 , n12529 , n12536 );
and ( n13228 , n12524 , n12536 );
or ( n13229 , n13226 , n13227 , n13228 );
and ( n13230 , n12514 , n12515 );
and ( n13231 , n12515 , n12517 );
and ( n13232 , n12514 , n12517 );
or ( n13233 , n13230 , n13231 , n13232 );
and ( n13234 , n12525 , n12526 );
and ( n13235 , n12526 , n12528 );
and ( n13236 , n12525 , n12528 );
or ( n13237 , n13234 , n13235 , n13236 );
xor ( n13238 , n13233 , n13237 );
and ( n13239 , n783 , n8669 );
and ( n13240 , n856 , n8243 );
xor ( n13241 , n13239 , n13240 );
and ( n13242 , n925 , n7662 );
xor ( n13243 , n13241 , n13242 );
xor ( n13244 , n13238 , n13243 );
xor ( n13245 , n13229 , n13244 );
and ( n13246 , n12532 , n12533 );
and ( n13247 , n12533 , n12535 );
and ( n13248 , n12532 , n12535 );
or ( n13249 , n13246 , n13247 , n13248 );
and ( n13250 , n632 , n10977 );
and ( n13251 , n671 , n10239 );
xor ( n13252 , n13250 , n13251 );
and ( n13253 , n715 , n9348 );
xor ( n13254 , n13252 , n13253 );
xor ( n13255 , n13249 , n13254 );
buf ( n13256 , n428 );
and ( n13257 , n599 , n13256 );
and ( n13258 , n608 , n12531 );
xor ( n13259 , n13257 , n13258 );
and ( n13260 , n611 , n11718 );
xor ( n13261 , n13259 , n13260 );
xor ( n13262 , n13255 , n13261 );
xor ( n13263 , n13245 , n13262 );
xor ( n13264 , n13225 , n13263 );
xor ( n13265 , n13194 , n13264 );
xor ( n13266 , n13142 , n13265 );
xor ( n13267 , n13059 , n13266 );
and ( n13268 , n12289 , n12293 );
and ( n13269 , n12293 , n12331 );
and ( n13270 , n12289 , n12331 );
or ( n13271 , n13268 , n13269 , n13270 );
and ( n13272 , n12342 , n12346 );
and ( n13273 , n12346 , n12415 );
and ( n13274 , n12342 , n12415 );
or ( n13275 , n13272 , n13273 , n13274 );
xor ( n13276 , n13271 , n13275 );
and ( n13277 , n12298 , n12302 );
and ( n13278 , n12302 , n12330 );
and ( n13279 , n12298 , n12330 );
or ( n13280 , n13277 , n13278 , n13279 );
and ( n13281 , n12307 , n12311 );
and ( n13282 , n12311 , n12329 );
and ( n13283 , n12307 , n12329 );
or ( n13284 , n13281 , n13282 , n13283 );
and ( n13285 , n12355 , n12370 );
and ( n13286 , n12370 , n12387 );
and ( n13287 , n12355 , n12387 );
or ( n13288 , n13285 , n13286 , n13287 );
xor ( n13289 , n13284 , n13288 );
and ( n13290 , n12316 , n12322 );
and ( n13291 , n12322 , n12328 );
and ( n13292 , n12316 , n12328 );
or ( n13293 , n13290 , n13291 , n13292 );
and ( n13294 , n12359 , n12363 );
and ( n13295 , n12363 , n12369 );
and ( n13296 , n12359 , n12369 );
or ( n13297 , n13294 , n13295 , n13296 );
xor ( n13298 , n13293 , n13297 );
and ( n13299 , n12324 , n12325 );
and ( n13300 , n12325 , n12327 );
and ( n13301 , n12324 , n12327 );
or ( n13302 , n13299 , n13300 , n13301 );
and ( n13303 , n11015 , n635 );
and ( n13304 , n11769 , n606 );
xor ( n13305 , n13303 , n13304 );
and ( n13306 , n12320 , n615 );
xor ( n13307 , n13305 , n13306 );
xor ( n13308 , n13302 , n13307 );
and ( n13309 , n8718 , n771 );
and ( n13310 , n9400 , n719 );
xor ( n13311 , n13309 , n13310 );
and ( n13312 , n10291 , n663 );
xor ( n13313 , n13311 , n13312 );
xor ( n13314 , n13308 , n13313 );
xor ( n13315 , n13298 , n13314 );
xor ( n13316 , n13289 , n13315 );
xor ( n13317 , n13280 , n13316 );
and ( n13318 , n12317 , n12318 );
and ( n13319 , n12318 , n12321 );
and ( n13320 , n12317 , n12321 );
or ( n13321 , n13318 , n13319 , n13320 );
buf ( n13322 , n428 );
and ( n13323 , n13322 , n612 );
xor ( n13324 , n13321 , n13323 );
xor ( n13325 , n13317 , n13324 );
xor ( n13326 , n13276 , n13325 );
xor ( n13327 , n13267 , n13326 );
xor ( n13328 , n13055 , n13327 );
and ( n13329 , n12273 , n12277 );
and ( n13330 , n12277 , n12542 );
and ( n13331 , n12273 , n12542 );
or ( n13332 , n13329 , n13330 , n13331 );
xor ( n13333 , n13328 , n13332 );
and ( n13334 , n12543 , n12547 );
and ( n13335 , n12548 , n12551 );
or ( n13336 , n13334 , n13335 );
xor ( n13337 , n13333 , n13336 );
buf ( n13338 , n13337 );
buf ( n13339 , n13338 );
not ( n13340 , n13339 );
nor ( n13341 , n13340 , n8739 );
xor ( n13342 , n13046 , n13341 );
and ( n13343 , n12269 , n12556 );
and ( n13344 , n12557 , n12560 );
or ( n13345 , n13343 , n13344 );
xor ( n13346 , n13342 , n13345 );
buf ( n13347 , n13346 );
buf ( n13348 , n13347 );
not ( n13349 , n13348 );
buf ( n13350 , n541 );
not ( n13351 , n13350 );
nor ( n13352 , n13349 , n13351 );
xor ( n13353 , n12806 , n13352 );
xor ( n13354 , n12572 , n12803 );
nor ( n13355 , n12564 , n13351 );
and ( n13356 , n13354 , n13355 );
xor ( n13357 , n13354 , n13355 );
xor ( n13358 , n12576 , n12801 );
nor ( n13359 , n11799 , n13351 );
and ( n13360 , n13358 , n13359 );
xor ( n13361 , n13358 , n13359 );
xor ( n13362 , n12580 , n12799 );
nor ( n13363 , n11050 , n13351 );
and ( n13364 , n13362 , n13363 );
xor ( n13365 , n13362 , n13363 );
xor ( n13366 , n12584 , n12797 );
nor ( n13367 , n10321 , n13351 );
and ( n13368 , n13366 , n13367 );
xor ( n13369 , n13366 , n13367 );
xor ( n13370 , n12588 , n12795 );
nor ( n13371 , n9429 , n13351 );
and ( n13372 , n13370 , n13371 );
xor ( n13373 , n13370 , n13371 );
xor ( n13374 , n12592 , n12793 );
nor ( n13375 , n8949 , n13351 );
and ( n13376 , n13374 , n13375 );
xor ( n13377 , n13374 , n13375 );
xor ( n13378 , n12596 , n12791 );
nor ( n13379 , n9437 , n13351 );
and ( n13380 , n13378 , n13379 );
xor ( n13381 , n13378 , n13379 );
xor ( n13382 , n12600 , n12789 );
nor ( n13383 , n9446 , n13351 );
and ( n13384 , n13382 , n13383 );
xor ( n13385 , n13382 , n13383 );
xor ( n13386 , n12604 , n12787 );
nor ( n13387 , n9455 , n13351 );
and ( n13388 , n13386 , n13387 );
xor ( n13389 , n13386 , n13387 );
xor ( n13390 , n12608 , n12785 );
nor ( n13391 , n9464 , n13351 );
and ( n13392 , n13390 , n13391 );
xor ( n13393 , n13390 , n13391 );
xor ( n13394 , n12612 , n12783 );
nor ( n13395 , n9473 , n13351 );
and ( n13396 , n13394 , n13395 );
xor ( n13397 , n13394 , n13395 );
xor ( n13398 , n12616 , n12781 );
nor ( n13399 , n9482 , n13351 );
and ( n13400 , n13398 , n13399 );
xor ( n13401 , n13398 , n13399 );
xor ( n13402 , n12620 , n12779 );
nor ( n13403 , n9491 , n13351 );
and ( n13404 , n13402 , n13403 );
xor ( n13405 , n13402 , n13403 );
xor ( n13406 , n12624 , n12777 );
nor ( n13407 , n9500 , n13351 );
and ( n13408 , n13406 , n13407 );
xor ( n13409 , n13406 , n13407 );
xor ( n13410 , n12628 , n12775 );
nor ( n13411 , n9509 , n13351 );
and ( n13412 , n13410 , n13411 );
xor ( n13413 , n13410 , n13411 );
xor ( n13414 , n12632 , n12773 );
nor ( n13415 , n9518 , n13351 );
and ( n13416 , n13414 , n13415 );
xor ( n13417 , n13414 , n13415 );
xor ( n13418 , n12636 , n12771 );
nor ( n13419 , n9527 , n13351 );
and ( n13420 , n13418 , n13419 );
xor ( n13421 , n13418 , n13419 );
xor ( n13422 , n12640 , n12769 );
nor ( n13423 , n9536 , n13351 );
and ( n13424 , n13422 , n13423 );
xor ( n13425 , n13422 , n13423 );
xor ( n13426 , n12644 , n12767 );
nor ( n13427 , n9545 , n13351 );
and ( n13428 , n13426 , n13427 );
xor ( n13429 , n13426 , n13427 );
xor ( n13430 , n12648 , n12765 );
nor ( n13431 , n9554 , n13351 );
and ( n13432 , n13430 , n13431 );
xor ( n13433 , n13430 , n13431 );
xor ( n13434 , n12652 , n12763 );
nor ( n13435 , n9563 , n13351 );
and ( n13436 , n13434 , n13435 );
xor ( n13437 , n13434 , n13435 );
xor ( n13438 , n12656 , n12761 );
nor ( n13439 , n9572 , n13351 );
and ( n13440 , n13438 , n13439 );
xor ( n13441 , n13438 , n13439 );
xor ( n13442 , n12660 , n12759 );
nor ( n13443 , n9581 , n13351 );
and ( n13444 , n13442 , n13443 );
xor ( n13445 , n13442 , n13443 );
xor ( n13446 , n12664 , n12757 );
nor ( n13447 , n9590 , n13351 );
and ( n13448 , n13446 , n13447 );
xor ( n13449 , n13446 , n13447 );
xor ( n13450 , n12668 , n12755 );
nor ( n13451 , n9599 , n13351 );
and ( n13452 , n13450 , n13451 );
xor ( n13453 , n13450 , n13451 );
xor ( n13454 , n12672 , n12753 );
nor ( n13455 , n9608 , n13351 );
and ( n13456 , n13454 , n13455 );
xor ( n13457 , n13454 , n13455 );
xor ( n13458 , n12676 , n12751 );
nor ( n13459 , n9617 , n13351 );
and ( n13460 , n13458 , n13459 );
xor ( n13461 , n13458 , n13459 );
xor ( n13462 , n12680 , n12749 );
nor ( n13463 , n9626 , n13351 );
and ( n13464 , n13462 , n13463 );
xor ( n13465 , n13462 , n13463 );
xor ( n13466 , n12684 , n12747 );
nor ( n13467 , n9635 , n13351 );
and ( n13468 , n13466 , n13467 );
xor ( n13469 , n13466 , n13467 );
xor ( n13470 , n12688 , n12745 );
nor ( n13471 , n9644 , n13351 );
and ( n13472 , n13470 , n13471 );
xor ( n13473 , n13470 , n13471 );
xor ( n13474 , n12692 , n12743 );
nor ( n13475 , n9653 , n13351 );
and ( n13476 , n13474 , n13475 );
xor ( n13477 , n13474 , n13475 );
xor ( n13478 , n12696 , n12741 );
nor ( n13479 , n9662 , n13351 );
and ( n13480 , n13478 , n13479 );
xor ( n13481 , n13478 , n13479 );
xor ( n13482 , n12700 , n12739 );
nor ( n13483 , n9671 , n13351 );
and ( n13484 , n13482 , n13483 );
xor ( n13485 , n13482 , n13483 );
xor ( n13486 , n12704 , n12737 );
nor ( n13487 , n9680 , n13351 );
and ( n13488 , n13486 , n13487 );
xor ( n13489 , n13486 , n13487 );
xor ( n13490 , n12708 , n12735 );
nor ( n13491 , n9689 , n13351 );
and ( n13492 , n13490 , n13491 );
xor ( n13493 , n13490 , n13491 );
xor ( n13494 , n12712 , n12733 );
nor ( n13495 , n9698 , n13351 );
and ( n13496 , n13494 , n13495 );
xor ( n13497 , n13494 , n13495 );
xor ( n13498 , n12716 , n12731 );
nor ( n13499 , n9707 , n13351 );
and ( n13500 , n13498 , n13499 );
xor ( n13501 , n13498 , n13499 );
xor ( n13502 , n12720 , n12729 );
nor ( n13503 , n9716 , n13351 );
and ( n13504 , n13502 , n13503 );
xor ( n13505 , n13502 , n13503 );
xor ( n13506 , n12724 , n12727 );
nor ( n13507 , n9725 , n13351 );
and ( n13508 , n13506 , n13507 );
xor ( n13509 , n13506 , n13507 );
xor ( n13510 , n12725 , n12726 );
nor ( n13511 , n9734 , n13351 );
and ( n13512 , n13510 , n13511 );
xor ( n13513 , n13510 , n13511 );
nor ( n13514 , n9752 , n12566 );
nor ( n13515 , n9743 , n13351 );
and ( n13516 , n13514 , n13515 );
and ( n13517 , n13513 , n13516 );
or ( n13518 , n13512 , n13517 );
and ( n13519 , n13509 , n13518 );
or ( n13520 , n13508 , n13519 );
and ( n13521 , n13505 , n13520 );
or ( n13522 , n13504 , n13521 );
and ( n13523 , n13501 , n13522 );
or ( n13524 , n13500 , n13523 );
and ( n13525 , n13497 , n13524 );
or ( n13526 , n13496 , n13525 );
and ( n13527 , n13493 , n13526 );
or ( n13528 , n13492 , n13527 );
and ( n13529 , n13489 , n13528 );
or ( n13530 , n13488 , n13529 );
and ( n13531 , n13485 , n13530 );
or ( n13532 , n13484 , n13531 );
and ( n13533 , n13481 , n13532 );
or ( n13534 , n13480 , n13533 );
and ( n13535 , n13477 , n13534 );
or ( n13536 , n13476 , n13535 );
and ( n13537 , n13473 , n13536 );
or ( n13538 , n13472 , n13537 );
and ( n13539 , n13469 , n13538 );
or ( n13540 , n13468 , n13539 );
and ( n13541 , n13465 , n13540 );
or ( n13542 , n13464 , n13541 );
and ( n13543 , n13461 , n13542 );
or ( n13544 , n13460 , n13543 );
and ( n13545 , n13457 , n13544 );
or ( n13546 , n13456 , n13545 );
and ( n13547 , n13453 , n13546 );
or ( n13548 , n13452 , n13547 );
and ( n13549 , n13449 , n13548 );
or ( n13550 , n13448 , n13549 );
and ( n13551 , n13445 , n13550 );
or ( n13552 , n13444 , n13551 );
and ( n13553 , n13441 , n13552 );
or ( n13554 , n13440 , n13553 );
and ( n13555 , n13437 , n13554 );
or ( n13556 , n13436 , n13555 );
and ( n13557 , n13433 , n13556 );
or ( n13558 , n13432 , n13557 );
and ( n13559 , n13429 , n13558 );
or ( n13560 , n13428 , n13559 );
and ( n13561 , n13425 , n13560 );
or ( n13562 , n13424 , n13561 );
and ( n13563 , n13421 , n13562 );
or ( n13564 , n13420 , n13563 );
and ( n13565 , n13417 , n13564 );
or ( n13566 , n13416 , n13565 );
and ( n13567 , n13413 , n13566 );
or ( n13568 , n13412 , n13567 );
and ( n13569 , n13409 , n13568 );
or ( n13570 , n13408 , n13569 );
and ( n13571 , n13405 , n13570 );
or ( n13572 , n13404 , n13571 );
and ( n13573 , n13401 , n13572 );
or ( n13574 , n13400 , n13573 );
and ( n13575 , n13397 , n13574 );
or ( n13576 , n13396 , n13575 );
and ( n13577 , n13393 , n13576 );
or ( n13578 , n13392 , n13577 );
and ( n13579 , n13389 , n13578 );
or ( n13580 , n13388 , n13579 );
and ( n13581 , n13385 , n13580 );
or ( n13582 , n13384 , n13581 );
and ( n13583 , n13381 , n13582 );
or ( n13584 , n13380 , n13583 );
and ( n13585 , n13377 , n13584 );
or ( n13586 , n13376 , n13585 );
and ( n13587 , n13373 , n13586 );
or ( n13588 , n13372 , n13587 );
and ( n13589 , n13369 , n13588 );
or ( n13590 , n13368 , n13589 );
and ( n13591 , n13365 , n13590 );
or ( n13592 , n13364 , n13591 );
and ( n13593 , n13361 , n13592 );
or ( n13594 , n13360 , n13593 );
and ( n13595 , n13357 , n13594 );
or ( n13596 , n13356 , n13595 );
xor ( n13597 , n13353 , n13596 );
buf ( n13598 , n491 );
not ( n13599 , n13598 );
nor ( n13600 , n601 , n13599 );
buf ( n13601 , n13600 );
nor ( n13602 , n622 , n12037 );
xor ( n13603 , n13601 , n13602 );
buf ( n13604 , n13603 );
nor ( n13605 , n646 , n11282 );
xor ( n13606 , n13604 , n13605 );
and ( n13607 , n12810 , n12811 );
buf ( n13608 , n13607 );
xor ( n13609 , n13606 , n13608 );
nor ( n13610 , n684 , n10547 );
xor ( n13611 , n13609 , n13610 );
and ( n13612 , n12813 , n12814 );
and ( n13613 , n12815 , n12817 );
or ( n13614 , n13612 , n13613 );
xor ( n13615 , n13611 , n13614 );
nor ( n13616 , n733 , n9829 );
xor ( n13617 , n13615 , n13616 );
and ( n13618 , n12818 , n12819 );
and ( n13619 , n12820 , n12823 );
or ( n13620 , n13618 , n13619 );
xor ( n13621 , n13617 , n13620 );
nor ( n13622 , n796 , n8955 );
xor ( n13623 , n13621 , n13622 );
and ( n13624 , n12824 , n12825 );
and ( n13625 , n12826 , n12829 );
or ( n13626 , n13624 , n13625 );
xor ( n13627 , n13623 , n13626 );
nor ( n13628 , n868 , n603 );
xor ( n13629 , n13627 , n13628 );
and ( n13630 , n12830 , n12831 );
and ( n13631 , n12832 , n12835 );
or ( n13632 , n13630 , n13631 );
xor ( n13633 , n13629 , n13632 );
nor ( n13634 , n958 , n652 );
xor ( n13635 , n13633 , n13634 );
and ( n13636 , n12836 , n12837 );
and ( n13637 , n12838 , n12841 );
or ( n13638 , n13636 , n13637 );
xor ( n13639 , n13635 , n13638 );
nor ( n13640 , n1062 , n624 );
xor ( n13641 , n13639 , n13640 );
and ( n13642 , n12842 , n12843 );
and ( n13643 , n12844 , n12847 );
or ( n13644 , n13642 , n13643 );
xor ( n13645 , n13641 , n13644 );
nor ( n13646 , n1176 , n648 );
xor ( n13647 , n13645 , n13646 );
and ( n13648 , n12848 , n12849 );
and ( n13649 , n12850 , n12853 );
or ( n13650 , n13648 , n13649 );
xor ( n13651 , n13647 , n13650 );
nor ( n13652 , n1303 , n686 );
xor ( n13653 , n13651 , n13652 );
and ( n13654 , n12854 , n12855 );
and ( n13655 , n12856 , n12859 );
or ( n13656 , n13654 , n13655 );
xor ( n13657 , n13653 , n13656 );
nor ( n13658 , n1445 , n735 );
xor ( n13659 , n13657 , n13658 );
and ( n13660 , n12860 , n12861 );
and ( n13661 , n12862 , n12865 );
or ( n13662 , n13660 , n13661 );
xor ( n13663 , n13659 , n13662 );
nor ( n13664 , n1598 , n798 );
xor ( n13665 , n13663 , n13664 );
and ( n13666 , n12866 , n12867 );
and ( n13667 , n12868 , n12871 );
or ( n13668 , n13666 , n13667 );
xor ( n13669 , n13665 , n13668 );
nor ( n13670 , n1766 , n870 );
xor ( n13671 , n13669 , n13670 );
and ( n13672 , n12872 , n12873 );
and ( n13673 , n12874 , n12877 );
or ( n13674 , n13672 , n13673 );
xor ( n13675 , n13671 , n13674 );
nor ( n13676 , n1945 , n960 );
xor ( n13677 , n13675 , n13676 );
and ( n13678 , n12878 , n12879 );
and ( n13679 , n12880 , n12883 );
or ( n13680 , n13678 , n13679 );
xor ( n13681 , n13677 , n13680 );
nor ( n13682 , n2137 , n1064 );
xor ( n13683 , n13681 , n13682 );
and ( n13684 , n12884 , n12885 );
and ( n13685 , n12886 , n12889 );
or ( n13686 , n13684 , n13685 );
xor ( n13687 , n13683 , n13686 );
nor ( n13688 , n2343 , n1178 );
xor ( n13689 , n13687 , n13688 );
and ( n13690 , n12890 , n12891 );
and ( n13691 , n12892 , n12895 );
or ( n13692 , n13690 , n13691 );
xor ( n13693 , n13689 , n13692 );
nor ( n13694 , n2566 , n1305 );
xor ( n13695 , n13693 , n13694 );
and ( n13696 , n12896 , n12897 );
and ( n13697 , n12898 , n12901 );
or ( n13698 , n13696 , n13697 );
xor ( n13699 , n13695 , n13698 );
nor ( n13700 , n2797 , n1447 );
xor ( n13701 , n13699 , n13700 );
and ( n13702 , n12902 , n12903 );
and ( n13703 , n12904 , n12907 );
or ( n13704 , n13702 , n13703 );
xor ( n13705 , n13701 , n13704 );
nor ( n13706 , n3043 , n1600 );
xor ( n13707 , n13705 , n13706 );
and ( n13708 , n12908 , n12909 );
and ( n13709 , n12910 , n12913 );
or ( n13710 , n13708 , n13709 );
xor ( n13711 , n13707 , n13710 );
nor ( n13712 , n3300 , n1768 );
xor ( n13713 , n13711 , n13712 );
and ( n13714 , n12914 , n12915 );
and ( n13715 , n12916 , n12919 );
or ( n13716 , n13714 , n13715 );
xor ( n13717 , n13713 , n13716 );
nor ( n13718 , n3570 , n1947 );
xor ( n13719 , n13717 , n13718 );
and ( n13720 , n12920 , n12921 );
and ( n13721 , n12922 , n12925 );
or ( n13722 , n13720 , n13721 );
xor ( n13723 , n13719 , n13722 );
nor ( n13724 , n3853 , n2139 );
xor ( n13725 , n13723 , n13724 );
and ( n13726 , n12926 , n12927 );
and ( n13727 , n12928 , n12931 );
or ( n13728 , n13726 , n13727 );
xor ( n13729 , n13725 , n13728 );
nor ( n13730 , n4151 , n2345 );
xor ( n13731 , n13729 , n13730 );
and ( n13732 , n12932 , n12933 );
and ( n13733 , n12934 , n12937 );
or ( n13734 , n13732 , n13733 );
xor ( n13735 , n13731 , n13734 );
nor ( n13736 , n4458 , n2568 );
xor ( n13737 , n13735 , n13736 );
and ( n13738 , n12938 , n12939 );
and ( n13739 , n12940 , n12943 );
or ( n13740 , n13738 , n13739 );
xor ( n13741 , n13737 , n13740 );
nor ( n13742 , n4786 , n2799 );
xor ( n13743 , n13741 , n13742 );
and ( n13744 , n12944 , n12945 );
and ( n13745 , n12946 , n12949 );
or ( n13746 , n13744 , n13745 );
xor ( n13747 , n13743 , n13746 );
nor ( n13748 , n5126 , n3045 );
xor ( n13749 , n13747 , n13748 );
and ( n13750 , n12950 , n12951 );
and ( n13751 , n12952 , n12955 );
or ( n13752 , n13750 , n13751 );
xor ( n13753 , n13749 , n13752 );
nor ( n13754 , n5477 , n3302 );
xor ( n13755 , n13753 , n13754 );
and ( n13756 , n12956 , n12957 );
and ( n13757 , n12958 , n12961 );
or ( n13758 , n13756 , n13757 );
xor ( n13759 , n13755 , n13758 );
nor ( n13760 , n5838 , n3572 );
xor ( n13761 , n13759 , n13760 );
and ( n13762 , n12962 , n12963 );
and ( n13763 , n12964 , n12967 );
or ( n13764 , n13762 , n13763 );
xor ( n13765 , n13761 , n13764 );
nor ( n13766 , n6212 , n3855 );
xor ( n13767 , n13765 , n13766 );
and ( n13768 , n12968 , n12969 );
and ( n13769 , n12970 , n12973 );
or ( n13770 , n13768 , n13769 );
xor ( n13771 , n13767 , n13770 );
nor ( n13772 , n6596 , n4153 );
xor ( n13773 , n13771 , n13772 );
and ( n13774 , n12974 , n12975 );
and ( n13775 , n12976 , n12979 );
or ( n13776 , n13774 , n13775 );
xor ( n13777 , n13773 , n13776 );
nor ( n13778 , n6997 , n4460 );
xor ( n13779 , n13777 , n13778 );
and ( n13780 , n12980 , n12981 );
and ( n13781 , n12982 , n12985 );
or ( n13782 , n13780 , n13781 );
xor ( n13783 , n13779 , n13782 );
nor ( n13784 , n7413 , n4788 );
xor ( n13785 , n13783 , n13784 );
and ( n13786 , n12986 , n12987 );
and ( n13787 , n12988 , n12991 );
or ( n13788 , n13786 , n13787 );
xor ( n13789 , n13785 , n13788 );
nor ( n13790 , n7841 , n5128 );
xor ( n13791 , n13789 , n13790 );
and ( n13792 , n12992 , n12993 );
and ( n13793 , n12994 , n12997 );
or ( n13794 , n13792 , n13793 );
xor ( n13795 , n13791 , n13794 );
nor ( n13796 , n8281 , n5479 );
xor ( n13797 , n13795 , n13796 );
and ( n13798 , n12998 , n12999 );
and ( n13799 , n13000 , n13003 );
or ( n13800 , n13798 , n13799 );
xor ( n13801 , n13797 , n13800 );
nor ( n13802 , n8737 , n5840 );
xor ( n13803 , n13801 , n13802 );
and ( n13804 , n13004 , n13005 );
and ( n13805 , n13006 , n13009 );
or ( n13806 , n13804 , n13805 );
xor ( n13807 , n13803 , n13806 );
nor ( n13808 , n9420 , n6214 );
xor ( n13809 , n13807 , n13808 );
and ( n13810 , n13010 , n13011 );
and ( n13811 , n13012 , n13015 );
or ( n13812 , n13810 , n13811 );
xor ( n13813 , n13809 , n13812 );
nor ( n13814 , n10312 , n6598 );
xor ( n13815 , n13813 , n13814 );
and ( n13816 , n13016 , n13017 );
and ( n13817 , n13018 , n13021 );
or ( n13818 , n13816 , n13817 );
xor ( n13819 , n13815 , n13818 );
nor ( n13820 , n11041 , n6999 );
xor ( n13821 , n13819 , n13820 );
and ( n13822 , n13022 , n13023 );
and ( n13823 , n13024 , n13027 );
or ( n13824 , n13822 , n13823 );
xor ( n13825 , n13821 , n13824 );
nor ( n13826 , n11790 , n7415 );
xor ( n13827 , n13825 , n13826 );
and ( n13828 , n13028 , n13029 );
and ( n13829 , n13030 , n13033 );
or ( n13830 , n13828 , n13829 );
xor ( n13831 , n13827 , n13830 );
nor ( n13832 , n12555 , n7843 );
xor ( n13833 , n13831 , n13832 );
and ( n13834 , n13034 , n13035 );
and ( n13835 , n13036 , n13039 );
or ( n13836 , n13834 , n13835 );
xor ( n13837 , n13833 , n13836 );
nor ( n13838 , n13340 , n8283 );
xor ( n13839 , n13837 , n13838 );
and ( n13840 , n13040 , n13041 );
and ( n13841 , n13042 , n13045 );
or ( n13842 , n13840 , n13841 );
xor ( n13843 , n13839 , n13842 );
and ( n13844 , n13271 , n13275 );
and ( n13845 , n13275 , n13325 );
and ( n13846 , n13271 , n13325 );
or ( n13847 , n13844 , n13845 , n13846 );
and ( n13848 , n13059 , n13266 );
and ( n13849 , n13266 , n13326 );
and ( n13850 , n13059 , n13326 );
or ( n13851 , n13848 , n13849 , n13850 );
xor ( n13852 , n13847 , n13851 );
and ( n13853 , n13063 , n13141 );
and ( n13854 , n13141 , n13265 );
and ( n13855 , n13063 , n13265 );
or ( n13856 , n13853 , n13854 , n13855 );
and ( n13857 , n13146 , n13193 );
and ( n13858 , n13193 , n13264 );
and ( n13859 , n13146 , n13264 );
or ( n13860 , n13857 , n13858 , n13859 );
and ( n13861 , n13076 , n13113 );
and ( n13862 , n13113 , n13139 );
and ( n13863 , n13076 , n13139 );
or ( n13864 , n13861 , n13862 , n13863 );
and ( n13865 , n13150 , n13154 );
and ( n13866 , n13154 , n13192 );
and ( n13867 , n13150 , n13192 );
or ( n13868 , n13865 , n13866 , n13867 );
xor ( n13869 , n13864 , n13868 );
and ( n13870 , n13118 , n13122 );
and ( n13871 , n13122 , n13138 );
and ( n13872 , n13118 , n13138 );
or ( n13873 , n13870 , n13871 , n13872 );
and ( n13874 , n13100 , n13105 );
and ( n13875 , n13105 , n13111 );
and ( n13876 , n13100 , n13111 );
or ( n13877 , n13874 , n13875 , n13876 );
and ( n13878 , n13090 , n13091 );
and ( n13879 , n13091 , n13093 );
and ( n13880 , n13090 , n13093 );
or ( n13881 , n13878 , n13879 , n13880 );
and ( n13882 , n13101 , n13102 );
and ( n13883 , n13102 , n13104 );
and ( n13884 , n13101 , n13104 );
or ( n13885 , n13882 , n13883 , n13884 );
xor ( n13886 , n13881 , n13885 );
and ( n13887 , n7385 , n1134 );
and ( n13888 , n7808 , n1034 );
xor ( n13889 , n13887 , n13888 );
and ( n13890 , n8079 , n940 );
xor ( n13891 , n13889 , n13890 );
xor ( n13892 , n13886 , n13891 );
xor ( n13893 , n13877 , n13892 );
and ( n13894 , n13107 , n13108 );
and ( n13895 , n13108 , n13110 );
and ( n13896 , n13107 , n13110 );
or ( n13897 , n13894 , n13895 , n13896 );
and ( n13898 , n6187 , n1551 );
and ( n13899 , n6569 , n1424 );
xor ( n13900 , n13898 , n13899 );
and ( n13901 , n6816 , n1254 );
xor ( n13902 , n13900 , n13901 );
xor ( n13903 , n13897 , n13902 );
and ( n13904 , n4959 , n2100 );
and ( n13905 , n5459 , n1882 );
xor ( n13906 , n13904 , n13905 );
and ( n13907 , n5819 , n1738 );
xor ( n13908 , n13906 , n13907 );
xor ( n13909 , n13903 , n13908 );
xor ( n13910 , n13893 , n13909 );
xor ( n13911 , n13873 , n13910 );
and ( n13912 , n13127 , n13131 );
and ( n13913 , n13131 , n13137 );
and ( n13914 , n13127 , n13137 );
or ( n13915 , n13912 , n13913 , n13914 );
and ( n13916 , n13163 , n13168 );
and ( n13917 , n13168 , n13174 );
and ( n13918 , n13163 , n13174 );
or ( n13919 , n13916 , n13917 , n13918 );
xor ( n13920 , n13915 , n13919 );
and ( n13921 , n13133 , n13134 );
and ( n13922 , n13134 , n13136 );
and ( n13923 , n13133 , n13136 );
or ( n13924 , n13921 , n13922 , n13923 );
and ( n13925 , n13164 , n13165 );
and ( n13926 , n13165 , n13167 );
and ( n13927 , n13164 , n13167 );
or ( n13928 , n13925 , n13926 , n13927 );
xor ( n13929 , n13924 , n13928 );
and ( n13930 , n4132 , n2739 );
and ( n13931 , n4438 , n2544 );
xor ( n13932 , n13930 , n13931 );
and ( n13933 , n4766 , n2298 );
xor ( n13934 , n13932 , n13933 );
xor ( n13935 , n13929 , n13934 );
xor ( n13936 , n13920 , n13935 );
xor ( n13937 , n13911 , n13936 );
xor ( n13938 , n13869 , n13937 );
xor ( n13939 , n13860 , n13938 );
and ( n13940 , n13198 , n13224 );
and ( n13941 , n13224 , n13263 );
and ( n13942 , n13198 , n13263 );
or ( n13943 , n13940 , n13941 , n13942 );
and ( n13944 , n13159 , n13175 );
and ( n13945 , n13175 , n13191 );
and ( n13946 , n13159 , n13191 );
or ( n13947 , n13944 , n13945 , n13946 );
and ( n13948 , n13202 , n13206 );
and ( n13949 , n13206 , n13223 );
and ( n13950 , n13202 , n13223 );
or ( n13951 , n13948 , n13949 , n13950 );
xor ( n13952 , n13947 , n13951 );
and ( n13953 , n13180 , n13184 );
and ( n13954 , n13184 , n13190 );
and ( n13955 , n13180 , n13190 );
or ( n13956 , n13953 , n13954 , n13955 );
and ( n13957 , n13170 , n13171 );
and ( n13958 , n13171 , n13173 );
and ( n13959 , n13170 , n13173 );
or ( n13960 , n13957 , n13958 , n13959 );
and ( n13961 , n3801 , n2981 );
buf ( n13962 , n13961 );
xor ( n13963 , n13960 , n13962 );
and ( n13964 , n2462 , n4403 );
and ( n13965 , n2779 , n4102 );
xor ( n13966 , n13964 , n13965 );
and ( n13967 , n3024 , n3749 );
xor ( n13968 , n13966 , n13967 );
xor ( n13969 , n13963 , n13968 );
xor ( n13970 , n13956 , n13969 );
and ( n13971 , n13186 , n13187 );
and ( n13972 , n13187 , n13189 );
and ( n13973 , n13186 , n13189 );
or ( n13974 , n13971 , n13972 , n13973 );
and ( n13975 , n13212 , n13213 );
and ( n13976 , n13213 , n13215 );
and ( n13977 , n13212 , n13215 );
or ( n13978 , n13975 , n13976 , n13977 );
xor ( n13979 , n13974 , n13978 );
and ( n13980 , n1933 , n5408 );
and ( n13981 , n2120 , n5103 );
xor ( n13982 , n13980 , n13981 );
and ( n13983 , n2324 , n4730 );
xor ( n13984 , n13982 , n13983 );
xor ( n13985 , n13979 , n13984 );
xor ( n13986 , n13970 , n13985 );
xor ( n13987 , n13952 , n13986 );
xor ( n13988 , n13943 , n13987 );
and ( n13989 , n13229 , n13244 );
and ( n13990 , n13244 , n13262 );
and ( n13991 , n13229 , n13262 );
or ( n13992 , n13989 , n13990 , n13991 );
and ( n13993 , n13211 , n13216 );
and ( n13994 , n13216 , n13222 );
and ( n13995 , n13211 , n13222 );
or ( n13996 , n13993 , n13994 , n13995 );
and ( n13997 , n13233 , n13237 );
and ( n13998 , n13237 , n13243 );
and ( n13999 , n13233 , n13243 );
or ( n14000 , n13997 , n13998 , n13999 );
xor ( n14001 , n13996 , n14000 );
and ( n14002 , n13218 , n13219 );
and ( n14003 , n13219 , n13221 );
and ( n14004 , n13218 , n13221 );
or ( n14005 , n14002 , n14003 , n14004 );
and ( n14006 , n1383 , n6504 );
and ( n14007 , n1580 , n6132 );
xor ( n14008 , n14006 , n14007 );
and ( n14009 , n1694 , n5765 );
xor ( n14010 , n14008 , n14009 );
xor ( n14011 , n14005 , n14010 );
and ( n14012 , n1047 , n7662 );
and ( n14013 , n1164 , n7310 );
xor ( n14014 , n14012 , n14013 );
and ( n14015 , n1287 , n6971 );
xor ( n14016 , n14014 , n14015 );
xor ( n14017 , n14011 , n14016 );
xor ( n14018 , n14001 , n14017 );
xor ( n14019 , n13992 , n14018 );
and ( n14020 , n13249 , n13254 );
and ( n14021 , n13254 , n13261 );
and ( n14022 , n13249 , n13261 );
or ( n14023 , n14020 , n14021 , n14022 );
and ( n14024 , n13239 , n13240 );
and ( n14025 , n13240 , n13242 );
and ( n14026 , n13239 , n13242 );
or ( n14027 , n14024 , n14025 , n14026 );
and ( n14028 , n13250 , n13251 );
and ( n14029 , n13251 , n13253 );
and ( n14030 , n13250 , n13253 );
or ( n14031 , n14028 , n14029 , n14030 );
xor ( n14032 , n14027 , n14031 );
and ( n14033 , n783 , n9348 );
and ( n14034 , n856 , n8669 );
xor ( n14035 , n14033 , n14034 );
and ( n14036 , n925 , n8243 );
xor ( n14037 , n14035 , n14036 );
xor ( n14038 , n14032 , n14037 );
xor ( n14039 , n14023 , n14038 );
and ( n14040 , n13257 , n13258 );
and ( n14041 , n13258 , n13260 );
and ( n14042 , n13257 , n13260 );
or ( n14043 , n14040 , n14041 , n14042 );
buf ( n14044 , n427 );
and ( n14045 , n599 , n14044 );
and ( n14046 , n608 , n13256 );
xor ( n14047 , n14045 , n14046 );
and ( n14048 , n611 , n12531 );
xor ( n14049 , n14047 , n14048 );
xor ( n14050 , n14043 , n14049 );
and ( n14051 , n632 , n11718 );
and ( n14052 , n671 , n10977 );
xor ( n14053 , n14051 , n14052 );
and ( n14054 , n715 , n10239 );
xor ( n14055 , n14053 , n14054 );
xor ( n14056 , n14050 , n14055 );
xor ( n14057 , n14039 , n14056 );
xor ( n14058 , n14019 , n14057 );
xor ( n14059 , n13988 , n14058 );
xor ( n14060 , n13939 , n14059 );
xor ( n14061 , n13856 , n14060 );
and ( n14062 , n13067 , n13071 );
and ( n14063 , n13071 , n13140 );
and ( n14064 , n13067 , n13140 );
or ( n14065 , n14062 , n14063 , n14064 );
and ( n14066 , n13280 , n13316 );
and ( n14067 , n13316 , n13324 );
and ( n14068 , n13280 , n13324 );
or ( n14069 , n14066 , n14067 , n14068 );
xor ( n14070 , n14065 , n14069 );
and ( n14071 , n13284 , n13288 );
and ( n14072 , n13288 , n13315 );
and ( n14073 , n13284 , n13315 );
or ( n14074 , n14071 , n14072 , n14073 );
and ( n14075 , n13293 , n13297 );
and ( n14076 , n13297 , n13314 );
and ( n14077 , n13293 , n13314 );
or ( n14078 , n14075 , n14076 , n14077 );
and ( n14079 , n13080 , n13095 );
and ( n14080 , n13095 , n13112 );
and ( n14081 , n13080 , n13112 );
or ( n14082 , n14079 , n14080 , n14081 );
xor ( n14083 , n14078 , n14082 );
and ( n14084 , n13302 , n13307 );
and ( n14085 , n13307 , n13313 );
and ( n14086 , n13302 , n13313 );
or ( n14087 , n14084 , n14085 , n14086 );
and ( n14088 , n13084 , n13088 );
and ( n14089 , n13088 , n13094 );
and ( n14090 , n13084 , n13094 );
or ( n14091 , n14088 , n14089 , n14090 );
xor ( n14092 , n14087 , n14091 );
and ( n14093 , n13309 , n13310 );
and ( n14094 , n13310 , n13312 );
and ( n14095 , n13309 , n13312 );
or ( n14096 , n14093 , n14094 , n14095 );
and ( n14097 , n11015 , n663 );
and ( n14098 , n11769 , n635 );
xor ( n14099 , n14097 , n14098 );
and ( n14100 , n12320 , n606 );
xor ( n14101 , n14099 , n14100 );
xor ( n14102 , n14096 , n14101 );
and ( n14103 , n8718 , n840 );
and ( n14104 , n9400 , n771 );
xor ( n14105 , n14103 , n14104 );
and ( n14106 , n10291 , n719 );
xor ( n14107 , n14105 , n14106 );
xor ( n14108 , n14102 , n14107 );
xor ( n14109 , n14092 , n14108 );
xor ( n14110 , n14083 , n14109 );
xor ( n14111 , n14074 , n14110 );
and ( n14112 , n13321 , n13323 );
and ( n14113 , n13303 , n13304 );
and ( n14114 , n13304 , n13306 );
and ( n14115 , n13303 , n13306 );
or ( n14116 , n14113 , n14114 , n14115 );
and ( n14117 , n13322 , n615 );
buf ( n14118 , n427 );
and ( n14119 , n14118 , n612 );
xor ( n14120 , n14117 , n14119 );
xor ( n14121 , n14116 , n14120 );
xor ( n14122 , n14112 , n14121 );
xor ( n14123 , n14111 , n14122 );
xor ( n14124 , n14070 , n14123 );
xor ( n14125 , n14061 , n14124 );
xor ( n14126 , n13852 , n14125 );
and ( n14127 , n13050 , n13054 );
and ( n14128 , n13054 , n13327 );
and ( n14129 , n13050 , n13327 );
or ( n14130 , n14127 , n14128 , n14129 );
xor ( n14131 , n14126 , n14130 );
and ( n14132 , n13328 , n13332 );
and ( n14133 , n13333 , n13336 );
or ( n14134 , n14132 , n14133 );
xor ( n14135 , n14131 , n14134 );
buf ( n14136 , n14135 );
buf ( n14137 , n14136 );
not ( n14138 , n14137 );
nor ( n14139 , n14138 , n8739 );
xor ( n14140 , n13843 , n14139 );
and ( n14141 , n13046 , n13341 );
and ( n14142 , n13342 , n13345 );
or ( n14143 , n14141 , n14142 );
xor ( n14144 , n14140 , n14143 );
buf ( n14145 , n14144 );
buf ( n14146 , n14145 );
not ( n14147 , n14146 );
buf ( n14148 , n542 );
not ( n14149 , n14148 );
nor ( n14150 , n14147 , n14149 );
xor ( n14151 , n13597 , n14150 );
xor ( n14152 , n13357 , n13594 );
nor ( n14153 , n13349 , n14149 );
and ( n14154 , n14152 , n14153 );
xor ( n14155 , n14152 , n14153 );
xor ( n14156 , n13361 , n13592 );
nor ( n14157 , n12564 , n14149 );
and ( n14158 , n14156 , n14157 );
xor ( n14159 , n14156 , n14157 );
xor ( n14160 , n13365 , n13590 );
nor ( n14161 , n11799 , n14149 );
and ( n14162 , n14160 , n14161 );
xor ( n14163 , n14160 , n14161 );
xor ( n14164 , n13369 , n13588 );
nor ( n14165 , n11050 , n14149 );
and ( n14166 , n14164 , n14165 );
xor ( n14167 , n14164 , n14165 );
xor ( n14168 , n13373 , n13586 );
nor ( n14169 , n10321 , n14149 );
and ( n14170 , n14168 , n14169 );
xor ( n14171 , n14168 , n14169 );
xor ( n14172 , n13377 , n13584 );
nor ( n14173 , n9429 , n14149 );
and ( n14174 , n14172 , n14173 );
xor ( n14175 , n14172 , n14173 );
xor ( n14176 , n13381 , n13582 );
nor ( n14177 , n8949 , n14149 );
and ( n14178 , n14176 , n14177 );
xor ( n14179 , n14176 , n14177 );
xor ( n14180 , n13385 , n13580 );
nor ( n14181 , n9437 , n14149 );
and ( n14182 , n14180 , n14181 );
xor ( n14183 , n14180 , n14181 );
xor ( n14184 , n13389 , n13578 );
nor ( n14185 , n9446 , n14149 );
and ( n14186 , n14184 , n14185 );
xor ( n14187 , n14184 , n14185 );
xor ( n14188 , n13393 , n13576 );
nor ( n14189 , n9455 , n14149 );
and ( n14190 , n14188 , n14189 );
xor ( n14191 , n14188 , n14189 );
xor ( n14192 , n13397 , n13574 );
nor ( n14193 , n9464 , n14149 );
and ( n14194 , n14192 , n14193 );
xor ( n14195 , n14192 , n14193 );
xor ( n14196 , n13401 , n13572 );
nor ( n14197 , n9473 , n14149 );
and ( n14198 , n14196 , n14197 );
xor ( n14199 , n14196 , n14197 );
xor ( n14200 , n13405 , n13570 );
nor ( n14201 , n9482 , n14149 );
and ( n14202 , n14200 , n14201 );
xor ( n14203 , n14200 , n14201 );
xor ( n14204 , n13409 , n13568 );
nor ( n14205 , n9491 , n14149 );
and ( n14206 , n14204 , n14205 );
xor ( n14207 , n14204 , n14205 );
xor ( n14208 , n13413 , n13566 );
nor ( n14209 , n9500 , n14149 );
and ( n14210 , n14208 , n14209 );
xor ( n14211 , n14208 , n14209 );
xor ( n14212 , n13417 , n13564 );
nor ( n14213 , n9509 , n14149 );
and ( n14214 , n14212 , n14213 );
xor ( n14215 , n14212 , n14213 );
xor ( n14216 , n13421 , n13562 );
nor ( n14217 , n9518 , n14149 );
and ( n14218 , n14216 , n14217 );
xor ( n14219 , n14216 , n14217 );
xor ( n14220 , n13425 , n13560 );
nor ( n14221 , n9527 , n14149 );
and ( n14222 , n14220 , n14221 );
xor ( n14223 , n14220 , n14221 );
xor ( n14224 , n13429 , n13558 );
nor ( n14225 , n9536 , n14149 );
and ( n14226 , n14224 , n14225 );
xor ( n14227 , n14224 , n14225 );
xor ( n14228 , n13433 , n13556 );
nor ( n14229 , n9545 , n14149 );
and ( n14230 , n14228 , n14229 );
xor ( n14231 , n14228 , n14229 );
xor ( n14232 , n13437 , n13554 );
nor ( n14233 , n9554 , n14149 );
and ( n14234 , n14232 , n14233 );
xor ( n14235 , n14232 , n14233 );
xor ( n14236 , n13441 , n13552 );
nor ( n14237 , n9563 , n14149 );
and ( n14238 , n14236 , n14237 );
xor ( n14239 , n14236 , n14237 );
xor ( n14240 , n13445 , n13550 );
nor ( n14241 , n9572 , n14149 );
and ( n14242 , n14240 , n14241 );
xor ( n14243 , n14240 , n14241 );
xor ( n14244 , n13449 , n13548 );
nor ( n14245 , n9581 , n14149 );
and ( n14246 , n14244 , n14245 );
xor ( n14247 , n14244 , n14245 );
xor ( n14248 , n13453 , n13546 );
nor ( n14249 , n9590 , n14149 );
and ( n14250 , n14248 , n14249 );
xor ( n14251 , n14248 , n14249 );
xor ( n14252 , n13457 , n13544 );
nor ( n14253 , n9599 , n14149 );
and ( n14254 , n14252 , n14253 );
xor ( n14255 , n14252 , n14253 );
xor ( n14256 , n13461 , n13542 );
nor ( n14257 , n9608 , n14149 );
and ( n14258 , n14256 , n14257 );
xor ( n14259 , n14256 , n14257 );
xor ( n14260 , n13465 , n13540 );
nor ( n14261 , n9617 , n14149 );
and ( n14262 , n14260 , n14261 );
xor ( n14263 , n14260 , n14261 );
xor ( n14264 , n13469 , n13538 );
nor ( n14265 , n9626 , n14149 );
and ( n14266 , n14264 , n14265 );
xor ( n14267 , n14264 , n14265 );
xor ( n14268 , n13473 , n13536 );
nor ( n14269 , n9635 , n14149 );
and ( n14270 , n14268 , n14269 );
xor ( n14271 , n14268 , n14269 );
xor ( n14272 , n13477 , n13534 );
nor ( n14273 , n9644 , n14149 );
and ( n14274 , n14272 , n14273 );
xor ( n14275 , n14272 , n14273 );
xor ( n14276 , n13481 , n13532 );
nor ( n14277 , n9653 , n14149 );
and ( n14278 , n14276 , n14277 );
xor ( n14279 , n14276 , n14277 );
xor ( n14280 , n13485 , n13530 );
nor ( n14281 , n9662 , n14149 );
and ( n14282 , n14280 , n14281 );
xor ( n14283 , n14280 , n14281 );
xor ( n14284 , n13489 , n13528 );
nor ( n14285 , n9671 , n14149 );
and ( n14286 , n14284 , n14285 );
xor ( n14287 , n14284 , n14285 );
xor ( n14288 , n13493 , n13526 );
nor ( n14289 , n9680 , n14149 );
and ( n14290 , n14288 , n14289 );
xor ( n14291 , n14288 , n14289 );
xor ( n14292 , n13497 , n13524 );
nor ( n14293 , n9689 , n14149 );
and ( n14294 , n14292 , n14293 );
xor ( n14295 , n14292 , n14293 );
xor ( n14296 , n13501 , n13522 );
nor ( n14297 , n9698 , n14149 );
and ( n14298 , n14296 , n14297 );
xor ( n14299 , n14296 , n14297 );
xor ( n14300 , n13505 , n13520 );
nor ( n14301 , n9707 , n14149 );
and ( n14302 , n14300 , n14301 );
xor ( n14303 , n14300 , n14301 );
xor ( n14304 , n13509 , n13518 );
nor ( n14305 , n9716 , n14149 );
and ( n14306 , n14304 , n14305 );
xor ( n14307 , n14304 , n14305 );
xor ( n14308 , n13513 , n13516 );
nor ( n14309 , n9725 , n14149 );
and ( n14310 , n14308 , n14309 );
xor ( n14311 , n14308 , n14309 );
xor ( n14312 , n13514 , n13515 );
nor ( n14313 , n9734 , n14149 );
and ( n14314 , n14312 , n14313 );
xor ( n14315 , n14312 , n14313 );
nor ( n14316 , n9752 , n13351 );
nor ( n14317 , n9743 , n14149 );
and ( n14318 , n14316 , n14317 );
and ( n14319 , n14315 , n14318 );
or ( n14320 , n14314 , n14319 );
and ( n14321 , n14311 , n14320 );
or ( n14322 , n14310 , n14321 );
and ( n14323 , n14307 , n14322 );
or ( n14324 , n14306 , n14323 );
and ( n14325 , n14303 , n14324 );
or ( n14326 , n14302 , n14325 );
and ( n14327 , n14299 , n14326 );
or ( n14328 , n14298 , n14327 );
and ( n14329 , n14295 , n14328 );
or ( n14330 , n14294 , n14329 );
and ( n14331 , n14291 , n14330 );
or ( n14332 , n14290 , n14331 );
and ( n14333 , n14287 , n14332 );
or ( n14334 , n14286 , n14333 );
and ( n14335 , n14283 , n14334 );
or ( n14336 , n14282 , n14335 );
and ( n14337 , n14279 , n14336 );
or ( n14338 , n14278 , n14337 );
and ( n14339 , n14275 , n14338 );
or ( n14340 , n14274 , n14339 );
and ( n14341 , n14271 , n14340 );
or ( n14342 , n14270 , n14341 );
and ( n14343 , n14267 , n14342 );
or ( n14344 , n14266 , n14343 );
and ( n14345 , n14263 , n14344 );
or ( n14346 , n14262 , n14345 );
and ( n14347 , n14259 , n14346 );
or ( n14348 , n14258 , n14347 );
and ( n14349 , n14255 , n14348 );
or ( n14350 , n14254 , n14349 );
and ( n14351 , n14251 , n14350 );
or ( n14352 , n14250 , n14351 );
and ( n14353 , n14247 , n14352 );
or ( n14354 , n14246 , n14353 );
and ( n14355 , n14243 , n14354 );
or ( n14356 , n14242 , n14355 );
and ( n14357 , n14239 , n14356 );
or ( n14358 , n14238 , n14357 );
and ( n14359 , n14235 , n14358 );
or ( n14360 , n14234 , n14359 );
and ( n14361 , n14231 , n14360 );
or ( n14362 , n14230 , n14361 );
and ( n14363 , n14227 , n14362 );
or ( n14364 , n14226 , n14363 );
and ( n14365 , n14223 , n14364 );
or ( n14366 , n14222 , n14365 );
and ( n14367 , n14219 , n14366 );
or ( n14368 , n14218 , n14367 );
and ( n14369 , n14215 , n14368 );
or ( n14370 , n14214 , n14369 );
and ( n14371 , n14211 , n14370 );
or ( n14372 , n14210 , n14371 );
and ( n14373 , n14207 , n14372 );
or ( n14374 , n14206 , n14373 );
and ( n14375 , n14203 , n14374 );
or ( n14376 , n14202 , n14375 );
and ( n14377 , n14199 , n14376 );
or ( n14378 , n14198 , n14377 );
and ( n14379 , n14195 , n14378 );
or ( n14380 , n14194 , n14379 );
and ( n14381 , n14191 , n14380 );
or ( n14382 , n14190 , n14381 );
and ( n14383 , n14187 , n14382 );
or ( n14384 , n14186 , n14383 );
and ( n14385 , n14183 , n14384 );
or ( n14386 , n14182 , n14385 );
and ( n14387 , n14179 , n14386 );
or ( n14388 , n14178 , n14387 );
and ( n14389 , n14175 , n14388 );
or ( n14390 , n14174 , n14389 );
and ( n14391 , n14171 , n14390 );
or ( n14392 , n14170 , n14391 );
and ( n14393 , n14167 , n14392 );
or ( n14394 , n14166 , n14393 );
and ( n14395 , n14163 , n14394 );
or ( n14396 , n14162 , n14395 );
and ( n14397 , n14159 , n14396 );
or ( n14398 , n14158 , n14397 );
and ( n14399 , n14155 , n14398 );
or ( n14400 , n14154 , n14399 );
xor ( n14401 , n14151 , n14400 );
buf ( n14402 , n490 );
not ( n14403 , n14402 );
nor ( n14404 , n601 , n14403 );
buf ( n14405 , n14404 );
nor ( n14406 , n622 , n12808 );
xor ( n14407 , n14405 , n14406 );
buf ( n14408 , n14407 );
nor ( n14409 , n646 , n12037 );
xor ( n14410 , n14408 , n14409 );
and ( n14411 , n13601 , n13602 );
buf ( n14412 , n14411 );
xor ( n14413 , n14410 , n14412 );
nor ( n14414 , n684 , n11282 );
xor ( n14415 , n14413 , n14414 );
and ( n14416 , n13604 , n13605 );
and ( n14417 , n13606 , n13608 );
or ( n14418 , n14416 , n14417 );
xor ( n14419 , n14415 , n14418 );
nor ( n14420 , n733 , n10547 );
xor ( n14421 , n14419 , n14420 );
and ( n14422 , n13609 , n13610 );
and ( n14423 , n13611 , n13614 );
or ( n14424 , n14422 , n14423 );
xor ( n14425 , n14421 , n14424 );
nor ( n14426 , n796 , n9829 );
xor ( n14427 , n14425 , n14426 );
and ( n14428 , n13615 , n13616 );
and ( n14429 , n13617 , n13620 );
or ( n14430 , n14428 , n14429 );
xor ( n14431 , n14427 , n14430 );
nor ( n14432 , n868 , n8955 );
xor ( n14433 , n14431 , n14432 );
and ( n14434 , n13621 , n13622 );
and ( n14435 , n13623 , n13626 );
or ( n14436 , n14434 , n14435 );
xor ( n14437 , n14433 , n14436 );
nor ( n14438 , n958 , n603 );
xor ( n14439 , n14437 , n14438 );
and ( n14440 , n13627 , n13628 );
and ( n14441 , n13629 , n13632 );
or ( n14442 , n14440 , n14441 );
xor ( n14443 , n14439 , n14442 );
nor ( n14444 , n1062 , n652 );
xor ( n14445 , n14443 , n14444 );
and ( n14446 , n13633 , n13634 );
and ( n14447 , n13635 , n13638 );
or ( n14448 , n14446 , n14447 );
xor ( n14449 , n14445 , n14448 );
nor ( n14450 , n1176 , n624 );
xor ( n14451 , n14449 , n14450 );
and ( n14452 , n13639 , n13640 );
and ( n14453 , n13641 , n13644 );
or ( n14454 , n14452 , n14453 );
xor ( n14455 , n14451 , n14454 );
nor ( n14456 , n1303 , n648 );
xor ( n14457 , n14455 , n14456 );
and ( n14458 , n13645 , n13646 );
and ( n14459 , n13647 , n13650 );
or ( n14460 , n14458 , n14459 );
xor ( n14461 , n14457 , n14460 );
nor ( n14462 , n1445 , n686 );
xor ( n14463 , n14461 , n14462 );
and ( n14464 , n13651 , n13652 );
and ( n14465 , n13653 , n13656 );
or ( n14466 , n14464 , n14465 );
xor ( n14467 , n14463 , n14466 );
nor ( n14468 , n1598 , n735 );
xor ( n14469 , n14467 , n14468 );
and ( n14470 , n13657 , n13658 );
and ( n14471 , n13659 , n13662 );
or ( n14472 , n14470 , n14471 );
xor ( n14473 , n14469 , n14472 );
nor ( n14474 , n1766 , n798 );
xor ( n14475 , n14473 , n14474 );
and ( n14476 , n13663 , n13664 );
and ( n14477 , n13665 , n13668 );
or ( n14478 , n14476 , n14477 );
xor ( n14479 , n14475 , n14478 );
nor ( n14480 , n1945 , n870 );
xor ( n14481 , n14479 , n14480 );
and ( n14482 , n13669 , n13670 );
and ( n14483 , n13671 , n13674 );
or ( n14484 , n14482 , n14483 );
xor ( n14485 , n14481 , n14484 );
nor ( n14486 , n2137 , n960 );
xor ( n14487 , n14485 , n14486 );
and ( n14488 , n13675 , n13676 );
and ( n14489 , n13677 , n13680 );
or ( n14490 , n14488 , n14489 );
xor ( n14491 , n14487 , n14490 );
nor ( n14492 , n2343 , n1064 );
xor ( n14493 , n14491 , n14492 );
and ( n14494 , n13681 , n13682 );
and ( n14495 , n13683 , n13686 );
or ( n14496 , n14494 , n14495 );
xor ( n14497 , n14493 , n14496 );
nor ( n14498 , n2566 , n1178 );
xor ( n14499 , n14497 , n14498 );
and ( n14500 , n13687 , n13688 );
and ( n14501 , n13689 , n13692 );
or ( n14502 , n14500 , n14501 );
xor ( n14503 , n14499 , n14502 );
nor ( n14504 , n2797 , n1305 );
xor ( n14505 , n14503 , n14504 );
and ( n14506 , n13693 , n13694 );
and ( n14507 , n13695 , n13698 );
or ( n14508 , n14506 , n14507 );
xor ( n14509 , n14505 , n14508 );
nor ( n14510 , n3043 , n1447 );
xor ( n14511 , n14509 , n14510 );
and ( n14512 , n13699 , n13700 );
and ( n14513 , n13701 , n13704 );
or ( n14514 , n14512 , n14513 );
xor ( n14515 , n14511 , n14514 );
nor ( n14516 , n3300 , n1600 );
xor ( n14517 , n14515 , n14516 );
and ( n14518 , n13705 , n13706 );
and ( n14519 , n13707 , n13710 );
or ( n14520 , n14518 , n14519 );
xor ( n14521 , n14517 , n14520 );
nor ( n14522 , n3570 , n1768 );
xor ( n14523 , n14521 , n14522 );
and ( n14524 , n13711 , n13712 );
and ( n14525 , n13713 , n13716 );
or ( n14526 , n14524 , n14525 );
xor ( n14527 , n14523 , n14526 );
nor ( n14528 , n3853 , n1947 );
xor ( n14529 , n14527 , n14528 );
and ( n14530 , n13717 , n13718 );
and ( n14531 , n13719 , n13722 );
or ( n14532 , n14530 , n14531 );
xor ( n14533 , n14529 , n14532 );
nor ( n14534 , n4151 , n2139 );
xor ( n14535 , n14533 , n14534 );
and ( n14536 , n13723 , n13724 );
and ( n14537 , n13725 , n13728 );
or ( n14538 , n14536 , n14537 );
xor ( n14539 , n14535 , n14538 );
nor ( n14540 , n4458 , n2345 );
xor ( n14541 , n14539 , n14540 );
and ( n14542 , n13729 , n13730 );
and ( n14543 , n13731 , n13734 );
or ( n14544 , n14542 , n14543 );
xor ( n14545 , n14541 , n14544 );
nor ( n14546 , n4786 , n2568 );
xor ( n14547 , n14545 , n14546 );
and ( n14548 , n13735 , n13736 );
and ( n14549 , n13737 , n13740 );
or ( n14550 , n14548 , n14549 );
xor ( n14551 , n14547 , n14550 );
nor ( n14552 , n5126 , n2799 );
xor ( n14553 , n14551 , n14552 );
and ( n14554 , n13741 , n13742 );
and ( n14555 , n13743 , n13746 );
or ( n14556 , n14554 , n14555 );
xor ( n14557 , n14553 , n14556 );
nor ( n14558 , n5477 , n3045 );
xor ( n14559 , n14557 , n14558 );
and ( n14560 , n13747 , n13748 );
and ( n14561 , n13749 , n13752 );
or ( n14562 , n14560 , n14561 );
xor ( n14563 , n14559 , n14562 );
nor ( n14564 , n5838 , n3302 );
xor ( n14565 , n14563 , n14564 );
and ( n14566 , n13753 , n13754 );
and ( n14567 , n13755 , n13758 );
or ( n14568 , n14566 , n14567 );
xor ( n14569 , n14565 , n14568 );
nor ( n14570 , n6212 , n3572 );
xor ( n14571 , n14569 , n14570 );
and ( n14572 , n13759 , n13760 );
and ( n14573 , n13761 , n13764 );
or ( n14574 , n14572 , n14573 );
xor ( n14575 , n14571 , n14574 );
nor ( n14576 , n6596 , n3855 );
xor ( n14577 , n14575 , n14576 );
and ( n14578 , n13765 , n13766 );
and ( n14579 , n13767 , n13770 );
or ( n14580 , n14578 , n14579 );
xor ( n14581 , n14577 , n14580 );
nor ( n14582 , n6997 , n4153 );
xor ( n14583 , n14581 , n14582 );
and ( n14584 , n13771 , n13772 );
and ( n14585 , n13773 , n13776 );
or ( n14586 , n14584 , n14585 );
xor ( n14587 , n14583 , n14586 );
nor ( n14588 , n7413 , n4460 );
xor ( n14589 , n14587 , n14588 );
and ( n14590 , n13777 , n13778 );
and ( n14591 , n13779 , n13782 );
or ( n14592 , n14590 , n14591 );
xor ( n14593 , n14589 , n14592 );
nor ( n14594 , n7841 , n4788 );
xor ( n14595 , n14593 , n14594 );
and ( n14596 , n13783 , n13784 );
and ( n14597 , n13785 , n13788 );
or ( n14598 , n14596 , n14597 );
xor ( n14599 , n14595 , n14598 );
nor ( n14600 , n8281 , n5128 );
xor ( n14601 , n14599 , n14600 );
and ( n14602 , n13789 , n13790 );
and ( n14603 , n13791 , n13794 );
or ( n14604 , n14602 , n14603 );
xor ( n14605 , n14601 , n14604 );
nor ( n14606 , n8737 , n5479 );
xor ( n14607 , n14605 , n14606 );
and ( n14608 , n13795 , n13796 );
and ( n14609 , n13797 , n13800 );
or ( n14610 , n14608 , n14609 );
xor ( n14611 , n14607 , n14610 );
nor ( n14612 , n9420 , n5840 );
xor ( n14613 , n14611 , n14612 );
and ( n14614 , n13801 , n13802 );
and ( n14615 , n13803 , n13806 );
or ( n14616 , n14614 , n14615 );
xor ( n14617 , n14613 , n14616 );
nor ( n14618 , n10312 , n6214 );
xor ( n14619 , n14617 , n14618 );
and ( n14620 , n13807 , n13808 );
and ( n14621 , n13809 , n13812 );
or ( n14622 , n14620 , n14621 );
xor ( n14623 , n14619 , n14622 );
nor ( n14624 , n11041 , n6598 );
xor ( n14625 , n14623 , n14624 );
and ( n14626 , n13813 , n13814 );
and ( n14627 , n13815 , n13818 );
or ( n14628 , n14626 , n14627 );
xor ( n14629 , n14625 , n14628 );
nor ( n14630 , n11790 , n6999 );
xor ( n14631 , n14629 , n14630 );
and ( n14632 , n13819 , n13820 );
and ( n14633 , n13821 , n13824 );
or ( n14634 , n14632 , n14633 );
xor ( n14635 , n14631 , n14634 );
nor ( n14636 , n12555 , n7415 );
xor ( n14637 , n14635 , n14636 );
and ( n14638 , n13825 , n13826 );
and ( n14639 , n13827 , n13830 );
or ( n14640 , n14638 , n14639 );
xor ( n14641 , n14637 , n14640 );
nor ( n14642 , n13340 , n7843 );
xor ( n14643 , n14641 , n14642 );
and ( n14644 , n13831 , n13832 );
and ( n14645 , n13833 , n13836 );
or ( n14646 , n14644 , n14645 );
xor ( n14647 , n14643 , n14646 );
nor ( n14648 , n14138 , n8283 );
xor ( n14649 , n14647 , n14648 );
and ( n14650 , n13837 , n13838 );
and ( n14651 , n13839 , n13842 );
or ( n14652 , n14650 , n14651 );
xor ( n14653 , n14649 , n14652 );
and ( n14654 , n14065 , n14069 );
and ( n14655 , n14069 , n14123 );
and ( n14656 , n14065 , n14123 );
or ( n14657 , n14654 , n14655 , n14656 );
and ( n14658 , n13856 , n14060 );
and ( n14659 , n14060 , n14124 );
and ( n14660 , n13856 , n14124 );
or ( n14661 , n14658 , n14659 , n14660 );
xor ( n14662 , n14657 , n14661 );
and ( n14663 , n13860 , n13938 );
and ( n14664 , n13938 , n14059 );
and ( n14665 , n13860 , n14059 );
or ( n14666 , n14663 , n14664 , n14665 );
and ( n14667 , n13943 , n13987 );
and ( n14668 , n13987 , n14058 );
and ( n14669 , n13943 , n14058 );
or ( n14670 , n14667 , n14668 , n14669 );
and ( n14671 , n13873 , n13910 );
and ( n14672 , n13910 , n13936 );
and ( n14673 , n13873 , n13936 );
or ( n14674 , n14671 , n14672 , n14673 );
and ( n14675 , n13947 , n13951 );
and ( n14676 , n13951 , n13986 );
and ( n14677 , n13947 , n13986 );
or ( n14678 , n14675 , n14676 , n14677 );
xor ( n14679 , n14674 , n14678 );
and ( n14680 , n13915 , n13919 );
and ( n14681 , n13919 , n13935 );
and ( n14682 , n13915 , n13935 );
or ( n14683 , n14680 , n14681 , n14682 );
and ( n14684 , n13897 , n13902 );
and ( n14685 , n13902 , n13908 );
and ( n14686 , n13897 , n13908 );
or ( n14687 , n14684 , n14685 , n14686 );
and ( n14688 , n13887 , n13888 );
and ( n14689 , n13888 , n13890 );
and ( n14690 , n13887 , n13890 );
or ( n14691 , n14688 , n14689 , n14690 );
and ( n14692 , n13898 , n13899 );
and ( n14693 , n13899 , n13901 );
and ( n14694 , n13898 , n13901 );
or ( n14695 , n14692 , n14693 , n14694 );
xor ( n14696 , n14691 , n14695 );
and ( n14697 , n7385 , n1254 );
and ( n14698 , n7808 , n1134 );
xor ( n14699 , n14697 , n14698 );
and ( n14700 , n8079 , n1034 );
xor ( n14701 , n14699 , n14700 );
xor ( n14702 , n14696 , n14701 );
xor ( n14703 , n14687 , n14702 );
and ( n14704 , n13904 , n13905 );
and ( n14705 , n13905 , n13907 );
and ( n14706 , n13904 , n13907 );
or ( n14707 , n14704 , n14705 , n14706 );
and ( n14708 , n6187 , n1738 );
and ( n14709 , n6569 , n1551 );
xor ( n14710 , n14708 , n14709 );
and ( n14711 , n6816 , n1424 );
xor ( n14712 , n14710 , n14711 );
xor ( n14713 , n14707 , n14712 );
and ( n14714 , n4959 , n2298 );
and ( n14715 , n5459 , n2100 );
xor ( n14716 , n14714 , n14715 );
and ( n14717 , n5819 , n1882 );
xor ( n14718 , n14716 , n14717 );
xor ( n14719 , n14713 , n14718 );
xor ( n14720 , n14703 , n14719 );
xor ( n14721 , n14683 , n14720 );
and ( n14722 , n13924 , n13928 );
and ( n14723 , n13928 , n13934 );
and ( n14724 , n13924 , n13934 );
or ( n14725 , n14722 , n14723 , n14724 );
and ( n14726 , n13960 , n13962 );
and ( n14727 , n13962 , n13968 );
and ( n14728 , n13960 , n13968 );
or ( n14729 , n14726 , n14727 , n14728 );
xor ( n14730 , n14725 , n14729 );
and ( n14731 , n13930 , n13931 );
and ( n14732 , n13931 , n13933 );
and ( n14733 , n13930 , n13933 );
or ( n14734 , n14731 , n14732 , n14733 );
and ( n14735 , n3182 , n3495 );
and ( n14736 , n3545 , n3271 );
and ( n14737 , n14735 , n14736 );
and ( n14738 , n14736 , n13961 );
and ( n14739 , n14735 , n13961 );
or ( n14740 , n14737 , n14738 , n14739 );
xor ( n14741 , n14734 , n14740 );
and ( n14742 , n4132 , n2981 );
and ( n14743 , n4438 , n2739 );
xor ( n14744 , n14742 , n14743 );
and ( n14745 , n4766 , n2544 );
xor ( n14746 , n14744 , n14745 );
xor ( n14747 , n14741 , n14746 );
xor ( n14748 , n14730 , n14747 );
xor ( n14749 , n14721 , n14748 );
xor ( n14750 , n14679 , n14749 );
xor ( n14751 , n14670 , n14750 );
and ( n14752 , n13992 , n14018 );
and ( n14753 , n14018 , n14057 );
and ( n14754 , n13992 , n14057 );
or ( n14755 , n14752 , n14753 , n14754 );
and ( n14756 , n13956 , n13969 );
and ( n14757 , n13969 , n13985 );
and ( n14758 , n13956 , n13985 );
or ( n14759 , n14756 , n14757 , n14758 );
and ( n14760 , n13996 , n14000 );
and ( n14761 , n14000 , n14017 );
and ( n14762 , n13996 , n14017 );
or ( n14763 , n14760 , n14761 , n14762 );
xor ( n14764 , n14759 , n14763 );
and ( n14765 , n13974 , n13978 );
and ( n14766 , n13978 , n13984 );
and ( n14767 , n13974 , n13984 );
or ( n14768 , n14765 , n14766 , n14767 );
and ( n14769 , n13964 , n13965 );
and ( n14770 , n13965 , n13967 );
and ( n14771 , n13964 , n13967 );
or ( n14772 , n14769 , n14770 , n14771 );
and ( n14773 , n3182 , n3749 );
buf ( n14774 , n3545 );
xor ( n14775 , n14773 , n14774 );
and ( n14776 , n3801 , n3271 );
xor ( n14777 , n14775 , n14776 );
xor ( n14778 , n14772 , n14777 );
and ( n14779 , n2462 , n4730 );
and ( n14780 , n2779 , n4403 );
xor ( n14781 , n14779 , n14780 );
and ( n14782 , n3024 , n4102 );
xor ( n14783 , n14781 , n14782 );
xor ( n14784 , n14778 , n14783 );
xor ( n14785 , n14768 , n14784 );
and ( n14786 , n14006 , n14007 );
and ( n14787 , n14007 , n14009 );
and ( n14788 , n14006 , n14009 );
or ( n14789 , n14786 , n14787 , n14788 );
and ( n14790 , n13980 , n13981 );
and ( n14791 , n13981 , n13983 );
and ( n14792 , n13980 , n13983 );
or ( n14793 , n14790 , n14791 , n14792 );
xor ( n14794 , n14789 , n14793 );
and ( n14795 , n1933 , n5765 );
and ( n14796 , n2120 , n5408 );
xor ( n14797 , n14795 , n14796 );
and ( n14798 , n2324 , n5103 );
xor ( n14799 , n14797 , n14798 );
xor ( n14800 , n14794 , n14799 );
xor ( n14801 , n14785 , n14800 );
xor ( n14802 , n14764 , n14801 );
xor ( n14803 , n14755 , n14802 );
and ( n14804 , n14023 , n14038 );
and ( n14805 , n14038 , n14056 );
and ( n14806 , n14023 , n14056 );
or ( n14807 , n14804 , n14805 , n14806 );
and ( n14808 , n14043 , n14049 );
and ( n14809 , n14049 , n14055 );
and ( n14810 , n14043 , n14055 );
or ( n14811 , n14808 , n14809 , n14810 );
and ( n14812 , n14033 , n14034 );
and ( n14813 , n14034 , n14036 );
and ( n14814 , n14033 , n14036 );
or ( n14815 , n14812 , n14813 , n14814 );
and ( n14816 , n14051 , n14052 );
and ( n14817 , n14052 , n14054 );
and ( n14818 , n14051 , n14054 );
or ( n14819 , n14816 , n14817 , n14818 );
xor ( n14820 , n14815 , n14819 );
and ( n14821 , n783 , n10239 );
and ( n14822 , n856 , n9348 );
xor ( n14823 , n14821 , n14822 );
and ( n14824 , n925 , n8669 );
xor ( n14825 , n14823 , n14824 );
xor ( n14826 , n14820 , n14825 );
xor ( n14827 , n14811 , n14826 );
and ( n14828 , n14045 , n14046 );
and ( n14829 , n14046 , n14048 );
and ( n14830 , n14045 , n14048 );
or ( n14831 , n14828 , n14829 , n14830 );
and ( n14832 , n632 , n12531 );
and ( n14833 , n671 , n11718 );
xor ( n14834 , n14832 , n14833 );
and ( n14835 , n715 , n10977 );
xor ( n14836 , n14834 , n14835 );
xor ( n14837 , n14831 , n14836 );
buf ( n14838 , n426 );
and ( n14839 , n599 , n14838 );
and ( n14840 , n608 , n14044 );
xor ( n14841 , n14839 , n14840 );
and ( n14842 , n611 , n13256 );
xor ( n14843 , n14841 , n14842 );
xor ( n14844 , n14837 , n14843 );
xor ( n14845 , n14827 , n14844 );
xor ( n14846 , n14807 , n14845 );
and ( n14847 , n14005 , n14010 );
and ( n14848 , n14010 , n14016 );
and ( n14849 , n14005 , n14016 );
or ( n14850 , n14847 , n14848 , n14849 );
and ( n14851 , n14027 , n14031 );
and ( n14852 , n14031 , n14037 );
and ( n14853 , n14027 , n14037 );
or ( n14854 , n14851 , n14852 , n14853 );
xor ( n14855 , n14850 , n14854 );
and ( n14856 , n14012 , n14013 );
and ( n14857 , n14013 , n14015 );
and ( n14858 , n14012 , n14015 );
or ( n14859 , n14856 , n14857 , n14858 );
and ( n14860 , n1383 , n6971 );
and ( n14861 , n1580 , n6504 );
xor ( n14862 , n14860 , n14861 );
and ( n14863 , n1694 , n6132 );
xor ( n14864 , n14862 , n14863 );
xor ( n14865 , n14859 , n14864 );
and ( n14866 , n1047 , n8243 );
and ( n14867 , n1164 , n7662 );
xor ( n14868 , n14866 , n14867 );
and ( n14869 , n1287 , n7310 );
xor ( n14870 , n14868 , n14869 );
xor ( n14871 , n14865 , n14870 );
xor ( n14872 , n14855 , n14871 );
xor ( n14873 , n14846 , n14872 );
xor ( n14874 , n14803 , n14873 );
xor ( n14875 , n14751 , n14874 );
xor ( n14876 , n14666 , n14875 );
and ( n14877 , n13864 , n13868 );
and ( n14878 , n13868 , n13937 );
and ( n14879 , n13864 , n13937 );
or ( n14880 , n14877 , n14878 , n14879 );
and ( n14881 , n14074 , n14110 );
and ( n14882 , n14110 , n14122 );
and ( n14883 , n14074 , n14122 );
or ( n14884 , n14881 , n14882 , n14883 );
xor ( n14885 , n14880 , n14884 );
and ( n14886 , n14078 , n14082 );
and ( n14887 , n14082 , n14109 );
and ( n14888 , n14078 , n14109 );
or ( n14889 , n14886 , n14887 , n14888 );
and ( n14890 , n14087 , n14091 );
and ( n14891 , n14091 , n14108 );
and ( n14892 , n14087 , n14108 );
or ( n14893 , n14890 , n14891 , n14892 );
and ( n14894 , n13877 , n13892 );
and ( n14895 , n13892 , n13909 );
and ( n14896 , n13877 , n13909 );
or ( n14897 , n14894 , n14895 , n14896 );
xor ( n14898 , n14893 , n14897 );
and ( n14899 , n14096 , n14101 );
and ( n14900 , n14101 , n14107 );
and ( n14901 , n14096 , n14107 );
or ( n14902 , n14899 , n14900 , n14901 );
and ( n14903 , n13881 , n13885 );
and ( n14904 , n13885 , n13891 );
and ( n14905 , n13881 , n13891 );
or ( n14906 , n14903 , n14904 , n14905 );
xor ( n14907 , n14902 , n14906 );
and ( n14908 , n14103 , n14104 );
and ( n14909 , n14104 , n14106 );
and ( n14910 , n14103 , n14106 );
or ( n14911 , n14908 , n14909 , n14910 );
and ( n14912 , n11015 , n719 );
and ( n14913 , n11769 , n663 );
xor ( n14914 , n14912 , n14913 );
and ( n14915 , n12320 , n635 );
xor ( n14916 , n14914 , n14915 );
xor ( n14917 , n14911 , n14916 );
and ( n14918 , n8718 , n940 );
and ( n14919 , n9400 , n840 );
xor ( n14920 , n14918 , n14919 );
and ( n14921 , n10291 , n771 );
xor ( n14922 , n14920 , n14921 );
xor ( n14923 , n14917 , n14922 );
xor ( n14924 , n14907 , n14923 );
xor ( n14925 , n14898 , n14924 );
xor ( n14926 , n14889 , n14925 );
and ( n14927 , n14112 , n14121 );
and ( n14928 , n14116 , n14120 );
and ( n14929 , n14097 , n14098 );
and ( n14930 , n14098 , n14100 );
and ( n14931 , n14097 , n14100 );
or ( n14932 , n14929 , n14930 , n14931 );
and ( n14933 , n14117 , n14119 );
xor ( n14934 , n14932 , n14933 );
and ( n14935 , n13322 , n606 );
and ( n14936 , n14118 , n615 );
xor ( n14937 , n14935 , n14936 );
buf ( n14938 , n426 );
and ( n14939 , n14938 , n612 );
xor ( n14940 , n14937 , n14939 );
xor ( n14941 , n14934 , n14940 );
xor ( n14942 , n14928 , n14941 );
xor ( n14943 , n14927 , n14942 );
xor ( n14944 , n14926 , n14943 );
xor ( n14945 , n14885 , n14944 );
xor ( n14946 , n14876 , n14945 );
xor ( n14947 , n14662 , n14946 );
and ( n14948 , n13847 , n13851 );
and ( n14949 , n13851 , n14125 );
and ( n14950 , n13847 , n14125 );
or ( n14951 , n14948 , n14949 , n14950 );
xor ( n14952 , n14947 , n14951 );
and ( n14953 , n14126 , n14130 );
and ( n14954 , n14131 , n14134 );
or ( n14955 , n14953 , n14954 );
xor ( n14956 , n14952 , n14955 );
buf ( n14957 , n14956 );
buf ( n14958 , n14957 );
not ( n14959 , n14958 );
nor ( n14960 , n14959 , n8739 );
xor ( n14961 , n14653 , n14960 );
and ( n14962 , n13843 , n14139 );
and ( n14963 , n14140 , n14143 );
or ( n14964 , n14962 , n14963 );
xor ( n14965 , n14961 , n14964 );
buf ( n14966 , n14965 );
buf ( n14967 , n14966 );
not ( n14968 , n14967 );
buf ( n14969 , n543 );
not ( n14970 , n14969 );
nor ( n14971 , n14968 , n14970 );
xor ( n14972 , n14401 , n14971 );
xor ( n14973 , n14155 , n14398 );
nor ( n14974 , n14147 , n14970 );
and ( n14975 , n14973 , n14974 );
xor ( n14976 , n14973 , n14974 );
xor ( n14977 , n14159 , n14396 );
nor ( n14978 , n13349 , n14970 );
and ( n14979 , n14977 , n14978 );
xor ( n14980 , n14977 , n14978 );
xor ( n14981 , n14163 , n14394 );
nor ( n14982 , n12564 , n14970 );
and ( n14983 , n14981 , n14982 );
xor ( n14984 , n14981 , n14982 );
xor ( n14985 , n14167 , n14392 );
nor ( n14986 , n11799 , n14970 );
and ( n14987 , n14985 , n14986 );
xor ( n14988 , n14985 , n14986 );
xor ( n14989 , n14171 , n14390 );
nor ( n14990 , n11050 , n14970 );
and ( n14991 , n14989 , n14990 );
xor ( n14992 , n14989 , n14990 );
xor ( n14993 , n14175 , n14388 );
nor ( n14994 , n10321 , n14970 );
and ( n14995 , n14993 , n14994 );
xor ( n14996 , n14993 , n14994 );
xor ( n14997 , n14179 , n14386 );
nor ( n14998 , n9429 , n14970 );
and ( n14999 , n14997 , n14998 );
xor ( n15000 , n14997 , n14998 );
xor ( n15001 , n14183 , n14384 );
nor ( n15002 , n8949 , n14970 );
and ( n15003 , n15001 , n15002 );
xor ( n15004 , n15001 , n15002 );
xor ( n15005 , n14187 , n14382 );
nor ( n15006 , n9437 , n14970 );
and ( n15007 , n15005 , n15006 );
xor ( n15008 , n15005 , n15006 );
xor ( n15009 , n14191 , n14380 );
nor ( n15010 , n9446 , n14970 );
and ( n15011 , n15009 , n15010 );
xor ( n15012 , n15009 , n15010 );
xor ( n15013 , n14195 , n14378 );
nor ( n15014 , n9455 , n14970 );
and ( n15015 , n15013 , n15014 );
xor ( n15016 , n15013 , n15014 );
xor ( n15017 , n14199 , n14376 );
nor ( n15018 , n9464 , n14970 );
and ( n15019 , n15017 , n15018 );
xor ( n15020 , n15017 , n15018 );
xor ( n15021 , n14203 , n14374 );
nor ( n15022 , n9473 , n14970 );
and ( n15023 , n15021 , n15022 );
xor ( n15024 , n15021 , n15022 );
xor ( n15025 , n14207 , n14372 );
nor ( n15026 , n9482 , n14970 );
and ( n15027 , n15025 , n15026 );
xor ( n15028 , n15025 , n15026 );
xor ( n15029 , n14211 , n14370 );
nor ( n15030 , n9491 , n14970 );
and ( n15031 , n15029 , n15030 );
xor ( n15032 , n15029 , n15030 );
xor ( n15033 , n14215 , n14368 );
nor ( n15034 , n9500 , n14970 );
and ( n15035 , n15033 , n15034 );
xor ( n15036 , n15033 , n15034 );
xor ( n15037 , n14219 , n14366 );
nor ( n15038 , n9509 , n14970 );
and ( n15039 , n15037 , n15038 );
xor ( n15040 , n15037 , n15038 );
xor ( n15041 , n14223 , n14364 );
nor ( n15042 , n9518 , n14970 );
and ( n15043 , n15041 , n15042 );
xor ( n15044 , n15041 , n15042 );
xor ( n15045 , n14227 , n14362 );
nor ( n15046 , n9527 , n14970 );
and ( n15047 , n15045 , n15046 );
xor ( n15048 , n15045 , n15046 );
xor ( n15049 , n14231 , n14360 );
nor ( n15050 , n9536 , n14970 );
and ( n15051 , n15049 , n15050 );
xor ( n15052 , n15049 , n15050 );
xor ( n15053 , n14235 , n14358 );
nor ( n15054 , n9545 , n14970 );
and ( n15055 , n15053 , n15054 );
xor ( n15056 , n15053 , n15054 );
xor ( n15057 , n14239 , n14356 );
nor ( n15058 , n9554 , n14970 );
and ( n15059 , n15057 , n15058 );
xor ( n15060 , n15057 , n15058 );
xor ( n15061 , n14243 , n14354 );
nor ( n15062 , n9563 , n14970 );
and ( n15063 , n15061 , n15062 );
xor ( n15064 , n15061 , n15062 );
xor ( n15065 , n14247 , n14352 );
nor ( n15066 , n9572 , n14970 );
and ( n15067 , n15065 , n15066 );
xor ( n15068 , n15065 , n15066 );
xor ( n15069 , n14251 , n14350 );
nor ( n15070 , n9581 , n14970 );
and ( n15071 , n15069 , n15070 );
xor ( n15072 , n15069 , n15070 );
xor ( n15073 , n14255 , n14348 );
nor ( n15074 , n9590 , n14970 );
and ( n15075 , n15073 , n15074 );
xor ( n15076 , n15073 , n15074 );
xor ( n15077 , n14259 , n14346 );
nor ( n15078 , n9599 , n14970 );
and ( n15079 , n15077 , n15078 );
xor ( n15080 , n15077 , n15078 );
xor ( n15081 , n14263 , n14344 );
nor ( n15082 , n9608 , n14970 );
and ( n15083 , n15081 , n15082 );
xor ( n15084 , n15081 , n15082 );
xor ( n15085 , n14267 , n14342 );
nor ( n15086 , n9617 , n14970 );
and ( n15087 , n15085 , n15086 );
xor ( n15088 , n15085 , n15086 );
xor ( n15089 , n14271 , n14340 );
nor ( n15090 , n9626 , n14970 );
and ( n15091 , n15089 , n15090 );
xor ( n15092 , n15089 , n15090 );
xor ( n15093 , n14275 , n14338 );
nor ( n15094 , n9635 , n14970 );
and ( n15095 , n15093 , n15094 );
xor ( n15096 , n15093 , n15094 );
xor ( n15097 , n14279 , n14336 );
nor ( n15098 , n9644 , n14970 );
and ( n15099 , n15097 , n15098 );
xor ( n15100 , n15097 , n15098 );
xor ( n15101 , n14283 , n14334 );
nor ( n15102 , n9653 , n14970 );
and ( n15103 , n15101 , n15102 );
xor ( n15104 , n15101 , n15102 );
xor ( n15105 , n14287 , n14332 );
nor ( n15106 , n9662 , n14970 );
and ( n15107 , n15105 , n15106 );
xor ( n15108 , n15105 , n15106 );
xor ( n15109 , n14291 , n14330 );
nor ( n15110 , n9671 , n14970 );
and ( n15111 , n15109 , n15110 );
xor ( n15112 , n15109 , n15110 );
xor ( n15113 , n14295 , n14328 );
nor ( n15114 , n9680 , n14970 );
and ( n15115 , n15113 , n15114 );
xor ( n15116 , n15113 , n15114 );
xor ( n15117 , n14299 , n14326 );
nor ( n15118 , n9689 , n14970 );
and ( n15119 , n15117 , n15118 );
xor ( n15120 , n15117 , n15118 );
xor ( n15121 , n14303 , n14324 );
nor ( n15122 , n9698 , n14970 );
and ( n15123 , n15121 , n15122 );
xor ( n15124 , n15121 , n15122 );
xor ( n15125 , n14307 , n14322 );
nor ( n15126 , n9707 , n14970 );
and ( n15127 , n15125 , n15126 );
xor ( n15128 , n15125 , n15126 );
xor ( n15129 , n14311 , n14320 );
nor ( n15130 , n9716 , n14970 );
and ( n15131 , n15129 , n15130 );
xor ( n15132 , n15129 , n15130 );
xor ( n15133 , n14315 , n14318 );
nor ( n15134 , n9725 , n14970 );
and ( n15135 , n15133 , n15134 );
xor ( n15136 , n15133 , n15134 );
xor ( n15137 , n14316 , n14317 );
nor ( n15138 , n9734 , n14970 );
and ( n15139 , n15137 , n15138 );
xor ( n15140 , n15137 , n15138 );
nor ( n15141 , n9752 , n14149 );
nor ( n15142 , n9743 , n14970 );
and ( n15143 , n15141 , n15142 );
and ( n15144 , n15140 , n15143 );
or ( n15145 , n15139 , n15144 );
and ( n15146 , n15136 , n15145 );
or ( n15147 , n15135 , n15146 );
and ( n15148 , n15132 , n15147 );
or ( n15149 , n15131 , n15148 );
and ( n15150 , n15128 , n15149 );
or ( n15151 , n15127 , n15150 );
and ( n15152 , n15124 , n15151 );
or ( n15153 , n15123 , n15152 );
and ( n15154 , n15120 , n15153 );
or ( n15155 , n15119 , n15154 );
and ( n15156 , n15116 , n15155 );
or ( n15157 , n15115 , n15156 );
and ( n15158 , n15112 , n15157 );
or ( n15159 , n15111 , n15158 );
and ( n15160 , n15108 , n15159 );
or ( n15161 , n15107 , n15160 );
and ( n15162 , n15104 , n15161 );
or ( n15163 , n15103 , n15162 );
and ( n15164 , n15100 , n15163 );
or ( n15165 , n15099 , n15164 );
and ( n15166 , n15096 , n15165 );
or ( n15167 , n15095 , n15166 );
and ( n15168 , n15092 , n15167 );
or ( n15169 , n15091 , n15168 );
and ( n15170 , n15088 , n15169 );
or ( n15171 , n15087 , n15170 );
and ( n15172 , n15084 , n15171 );
or ( n15173 , n15083 , n15172 );
and ( n15174 , n15080 , n15173 );
or ( n15175 , n15079 , n15174 );
and ( n15176 , n15076 , n15175 );
or ( n15177 , n15075 , n15176 );
and ( n15178 , n15072 , n15177 );
or ( n15179 , n15071 , n15178 );
and ( n15180 , n15068 , n15179 );
or ( n15181 , n15067 , n15180 );
and ( n15182 , n15064 , n15181 );
or ( n15183 , n15063 , n15182 );
and ( n15184 , n15060 , n15183 );
or ( n15185 , n15059 , n15184 );
and ( n15186 , n15056 , n15185 );
or ( n15187 , n15055 , n15186 );
and ( n15188 , n15052 , n15187 );
or ( n15189 , n15051 , n15188 );
and ( n15190 , n15048 , n15189 );
or ( n15191 , n15047 , n15190 );
and ( n15192 , n15044 , n15191 );
or ( n15193 , n15043 , n15192 );
and ( n15194 , n15040 , n15193 );
or ( n15195 , n15039 , n15194 );
and ( n15196 , n15036 , n15195 );
or ( n15197 , n15035 , n15196 );
and ( n15198 , n15032 , n15197 );
or ( n15199 , n15031 , n15198 );
and ( n15200 , n15028 , n15199 );
or ( n15201 , n15027 , n15200 );
and ( n15202 , n15024 , n15201 );
or ( n15203 , n15023 , n15202 );
and ( n15204 , n15020 , n15203 );
or ( n15205 , n15019 , n15204 );
and ( n15206 , n15016 , n15205 );
or ( n15207 , n15015 , n15206 );
and ( n15208 , n15012 , n15207 );
or ( n15209 , n15011 , n15208 );
and ( n15210 , n15008 , n15209 );
or ( n15211 , n15007 , n15210 );
and ( n15212 , n15004 , n15211 );
or ( n15213 , n15003 , n15212 );
and ( n15214 , n15000 , n15213 );
or ( n15215 , n14999 , n15214 );
and ( n15216 , n14996 , n15215 );
or ( n15217 , n14995 , n15216 );
and ( n15218 , n14992 , n15217 );
or ( n15219 , n14991 , n15218 );
and ( n15220 , n14988 , n15219 );
or ( n15221 , n14987 , n15220 );
and ( n15222 , n14984 , n15221 );
or ( n15223 , n14983 , n15222 );
and ( n15224 , n14980 , n15223 );
or ( n15225 , n14979 , n15224 );
and ( n15226 , n14976 , n15225 );
or ( n15227 , n14975 , n15226 );
xor ( n15228 , n14972 , n15227 );
buf ( n15229 , n489 );
not ( n15230 , n15229 );
nor ( n15231 , n601 , n15230 );
buf ( n15232 , n15231 );
nor ( n15233 , n622 , n13599 );
xor ( n15234 , n15232 , n15233 );
buf ( n15235 , n15234 );
nor ( n15236 , n646 , n12808 );
xor ( n15237 , n15235 , n15236 );
and ( n15238 , n14405 , n14406 );
buf ( n15239 , n15238 );
xor ( n15240 , n15237 , n15239 );
nor ( n15241 , n684 , n12037 );
xor ( n15242 , n15240 , n15241 );
and ( n15243 , n14408 , n14409 );
and ( n15244 , n14410 , n14412 );
or ( n15245 , n15243 , n15244 );
xor ( n15246 , n15242 , n15245 );
nor ( n15247 , n733 , n11282 );
xor ( n15248 , n15246 , n15247 );
and ( n15249 , n14413 , n14414 );
and ( n15250 , n14415 , n14418 );
or ( n15251 , n15249 , n15250 );
xor ( n15252 , n15248 , n15251 );
nor ( n15253 , n796 , n10547 );
xor ( n15254 , n15252 , n15253 );
and ( n15255 , n14419 , n14420 );
and ( n15256 , n14421 , n14424 );
or ( n15257 , n15255 , n15256 );
xor ( n15258 , n15254 , n15257 );
nor ( n15259 , n868 , n9829 );
xor ( n15260 , n15258 , n15259 );
and ( n15261 , n14425 , n14426 );
and ( n15262 , n14427 , n14430 );
or ( n15263 , n15261 , n15262 );
xor ( n15264 , n15260 , n15263 );
nor ( n15265 , n958 , n8955 );
xor ( n15266 , n15264 , n15265 );
and ( n15267 , n14431 , n14432 );
and ( n15268 , n14433 , n14436 );
or ( n15269 , n15267 , n15268 );
xor ( n15270 , n15266 , n15269 );
nor ( n15271 , n1062 , n603 );
xor ( n15272 , n15270 , n15271 );
and ( n15273 , n14437 , n14438 );
and ( n15274 , n14439 , n14442 );
or ( n15275 , n15273 , n15274 );
xor ( n15276 , n15272 , n15275 );
nor ( n15277 , n1176 , n652 );
xor ( n15278 , n15276 , n15277 );
and ( n15279 , n14443 , n14444 );
and ( n15280 , n14445 , n14448 );
or ( n15281 , n15279 , n15280 );
xor ( n15282 , n15278 , n15281 );
nor ( n15283 , n1303 , n624 );
xor ( n15284 , n15282 , n15283 );
and ( n15285 , n14449 , n14450 );
and ( n15286 , n14451 , n14454 );
or ( n15287 , n15285 , n15286 );
xor ( n15288 , n15284 , n15287 );
nor ( n15289 , n1445 , n648 );
xor ( n15290 , n15288 , n15289 );
and ( n15291 , n14455 , n14456 );
and ( n15292 , n14457 , n14460 );
or ( n15293 , n15291 , n15292 );
xor ( n15294 , n15290 , n15293 );
nor ( n15295 , n1598 , n686 );
xor ( n15296 , n15294 , n15295 );
and ( n15297 , n14461 , n14462 );
and ( n15298 , n14463 , n14466 );
or ( n15299 , n15297 , n15298 );
xor ( n15300 , n15296 , n15299 );
nor ( n15301 , n1766 , n735 );
xor ( n15302 , n15300 , n15301 );
and ( n15303 , n14467 , n14468 );
and ( n15304 , n14469 , n14472 );
or ( n15305 , n15303 , n15304 );
xor ( n15306 , n15302 , n15305 );
nor ( n15307 , n1945 , n798 );
xor ( n15308 , n15306 , n15307 );
and ( n15309 , n14473 , n14474 );
and ( n15310 , n14475 , n14478 );
or ( n15311 , n15309 , n15310 );
xor ( n15312 , n15308 , n15311 );
nor ( n15313 , n2137 , n870 );
xor ( n15314 , n15312 , n15313 );
and ( n15315 , n14479 , n14480 );
and ( n15316 , n14481 , n14484 );
or ( n15317 , n15315 , n15316 );
xor ( n15318 , n15314 , n15317 );
nor ( n15319 , n2343 , n960 );
xor ( n15320 , n15318 , n15319 );
and ( n15321 , n14485 , n14486 );
and ( n15322 , n14487 , n14490 );
or ( n15323 , n15321 , n15322 );
xor ( n15324 , n15320 , n15323 );
nor ( n15325 , n2566 , n1064 );
xor ( n15326 , n15324 , n15325 );
and ( n15327 , n14491 , n14492 );
and ( n15328 , n14493 , n14496 );
or ( n15329 , n15327 , n15328 );
xor ( n15330 , n15326 , n15329 );
nor ( n15331 , n2797 , n1178 );
xor ( n15332 , n15330 , n15331 );
and ( n15333 , n14497 , n14498 );
and ( n15334 , n14499 , n14502 );
or ( n15335 , n15333 , n15334 );
xor ( n15336 , n15332 , n15335 );
nor ( n15337 , n3043 , n1305 );
xor ( n15338 , n15336 , n15337 );
and ( n15339 , n14503 , n14504 );
and ( n15340 , n14505 , n14508 );
or ( n15341 , n15339 , n15340 );
xor ( n15342 , n15338 , n15341 );
nor ( n15343 , n3300 , n1447 );
xor ( n15344 , n15342 , n15343 );
and ( n15345 , n14509 , n14510 );
and ( n15346 , n14511 , n14514 );
or ( n15347 , n15345 , n15346 );
xor ( n15348 , n15344 , n15347 );
nor ( n15349 , n3570 , n1600 );
xor ( n15350 , n15348 , n15349 );
and ( n15351 , n14515 , n14516 );
and ( n15352 , n14517 , n14520 );
or ( n15353 , n15351 , n15352 );
xor ( n15354 , n15350 , n15353 );
nor ( n15355 , n3853 , n1768 );
xor ( n15356 , n15354 , n15355 );
and ( n15357 , n14521 , n14522 );
and ( n15358 , n14523 , n14526 );
or ( n15359 , n15357 , n15358 );
xor ( n15360 , n15356 , n15359 );
nor ( n15361 , n4151 , n1947 );
xor ( n15362 , n15360 , n15361 );
and ( n15363 , n14527 , n14528 );
and ( n15364 , n14529 , n14532 );
or ( n15365 , n15363 , n15364 );
xor ( n15366 , n15362 , n15365 );
nor ( n15367 , n4458 , n2139 );
xor ( n15368 , n15366 , n15367 );
and ( n15369 , n14533 , n14534 );
and ( n15370 , n14535 , n14538 );
or ( n15371 , n15369 , n15370 );
xor ( n15372 , n15368 , n15371 );
nor ( n15373 , n4786 , n2345 );
xor ( n15374 , n15372 , n15373 );
and ( n15375 , n14539 , n14540 );
and ( n15376 , n14541 , n14544 );
or ( n15377 , n15375 , n15376 );
xor ( n15378 , n15374 , n15377 );
nor ( n15379 , n5126 , n2568 );
xor ( n15380 , n15378 , n15379 );
and ( n15381 , n14545 , n14546 );
and ( n15382 , n14547 , n14550 );
or ( n15383 , n15381 , n15382 );
xor ( n15384 , n15380 , n15383 );
nor ( n15385 , n5477 , n2799 );
xor ( n15386 , n15384 , n15385 );
and ( n15387 , n14551 , n14552 );
and ( n15388 , n14553 , n14556 );
or ( n15389 , n15387 , n15388 );
xor ( n15390 , n15386 , n15389 );
nor ( n15391 , n5838 , n3045 );
xor ( n15392 , n15390 , n15391 );
and ( n15393 , n14557 , n14558 );
and ( n15394 , n14559 , n14562 );
or ( n15395 , n15393 , n15394 );
xor ( n15396 , n15392 , n15395 );
nor ( n15397 , n6212 , n3302 );
xor ( n15398 , n15396 , n15397 );
and ( n15399 , n14563 , n14564 );
and ( n15400 , n14565 , n14568 );
or ( n15401 , n15399 , n15400 );
xor ( n15402 , n15398 , n15401 );
nor ( n15403 , n6596 , n3572 );
xor ( n15404 , n15402 , n15403 );
and ( n15405 , n14569 , n14570 );
and ( n15406 , n14571 , n14574 );
or ( n15407 , n15405 , n15406 );
xor ( n15408 , n15404 , n15407 );
nor ( n15409 , n6997 , n3855 );
xor ( n15410 , n15408 , n15409 );
and ( n15411 , n14575 , n14576 );
and ( n15412 , n14577 , n14580 );
or ( n15413 , n15411 , n15412 );
xor ( n15414 , n15410 , n15413 );
nor ( n15415 , n7413 , n4153 );
xor ( n15416 , n15414 , n15415 );
and ( n15417 , n14581 , n14582 );
and ( n15418 , n14583 , n14586 );
or ( n15419 , n15417 , n15418 );
xor ( n15420 , n15416 , n15419 );
nor ( n15421 , n7841 , n4460 );
xor ( n15422 , n15420 , n15421 );
and ( n15423 , n14587 , n14588 );
and ( n15424 , n14589 , n14592 );
or ( n15425 , n15423 , n15424 );
xor ( n15426 , n15422 , n15425 );
nor ( n15427 , n8281 , n4788 );
xor ( n15428 , n15426 , n15427 );
and ( n15429 , n14593 , n14594 );
and ( n15430 , n14595 , n14598 );
or ( n15431 , n15429 , n15430 );
xor ( n15432 , n15428 , n15431 );
nor ( n15433 , n8737 , n5128 );
xor ( n15434 , n15432 , n15433 );
and ( n15435 , n14599 , n14600 );
and ( n15436 , n14601 , n14604 );
or ( n15437 , n15435 , n15436 );
xor ( n15438 , n15434 , n15437 );
nor ( n15439 , n9420 , n5479 );
xor ( n15440 , n15438 , n15439 );
and ( n15441 , n14605 , n14606 );
and ( n15442 , n14607 , n14610 );
or ( n15443 , n15441 , n15442 );
xor ( n15444 , n15440 , n15443 );
nor ( n15445 , n10312 , n5840 );
xor ( n15446 , n15444 , n15445 );
and ( n15447 , n14611 , n14612 );
and ( n15448 , n14613 , n14616 );
or ( n15449 , n15447 , n15448 );
xor ( n15450 , n15446 , n15449 );
nor ( n15451 , n11041 , n6214 );
xor ( n15452 , n15450 , n15451 );
and ( n15453 , n14617 , n14618 );
and ( n15454 , n14619 , n14622 );
or ( n15455 , n15453 , n15454 );
xor ( n15456 , n15452 , n15455 );
nor ( n15457 , n11790 , n6598 );
xor ( n15458 , n15456 , n15457 );
and ( n15459 , n14623 , n14624 );
and ( n15460 , n14625 , n14628 );
or ( n15461 , n15459 , n15460 );
xor ( n15462 , n15458 , n15461 );
nor ( n15463 , n12555 , n6999 );
xor ( n15464 , n15462 , n15463 );
and ( n15465 , n14629 , n14630 );
and ( n15466 , n14631 , n14634 );
or ( n15467 , n15465 , n15466 );
xor ( n15468 , n15464 , n15467 );
nor ( n15469 , n13340 , n7415 );
xor ( n15470 , n15468 , n15469 );
and ( n15471 , n14635 , n14636 );
and ( n15472 , n14637 , n14640 );
or ( n15473 , n15471 , n15472 );
xor ( n15474 , n15470 , n15473 );
nor ( n15475 , n14138 , n7843 );
xor ( n15476 , n15474 , n15475 );
and ( n15477 , n14641 , n14642 );
and ( n15478 , n14643 , n14646 );
or ( n15479 , n15477 , n15478 );
xor ( n15480 , n15476 , n15479 );
nor ( n15481 , n14959 , n8283 );
xor ( n15482 , n15480 , n15481 );
and ( n15483 , n14647 , n14648 );
and ( n15484 , n14649 , n14652 );
or ( n15485 , n15483 , n15484 );
xor ( n15486 , n15482 , n15485 );
and ( n15487 , n14666 , n14875 );
and ( n15488 , n14875 , n14945 );
and ( n15489 , n14666 , n14945 );
or ( n15490 , n15487 , n15488 , n15489 );
and ( n15491 , n14670 , n14750 );
and ( n15492 , n14750 , n14874 );
and ( n15493 , n14670 , n14874 );
or ( n15494 , n15491 , n15492 , n15493 );
and ( n15495 , n14755 , n14802 );
and ( n15496 , n14802 , n14873 );
and ( n15497 , n14755 , n14873 );
or ( n15498 , n15495 , n15496 , n15497 );
and ( n15499 , n14683 , n14720 );
and ( n15500 , n14720 , n14748 );
and ( n15501 , n14683 , n14748 );
or ( n15502 , n15499 , n15500 , n15501 );
and ( n15503 , n14759 , n14763 );
and ( n15504 , n14763 , n14801 );
and ( n15505 , n14759 , n14801 );
or ( n15506 , n15503 , n15504 , n15505 );
xor ( n15507 , n15502 , n15506 );
and ( n15508 , n14725 , n14729 );
and ( n15509 , n14729 , n14747 );
and ( n15510 , n14725 , n14747 );
or ( n15511 , n15508 , n15509 , n15510 );
and ( n15512 , n14707 , n14712 );
and ( n15513 , n14712 , n14718 );
and ( n15514 , n14707 , n14718 );
or ( n15515 , n15512 , n15513 , n15514 );
and ( n15516 , n14697 , n14698 );
and ( n15517 , n14698 , n14700 );
and ( n15518 , n14697 , n14700 );
or ( n15519 , n15516 , n15517 , n15518 );
and ( n15520 , n14708 , n14709 );
and ( n15521 , n14709 , n14711 );
and ( n15522 , n14708 , n14711 );
or ( n15523 , n15520 , n15521 , n15522 );
xor ( n15524 , n15519 , n15523 );
and ( n15525 , n7385 , n1424 );
and ( n15526 , n7808 , n1254 );
xor ( n15527 , n15525 , n15526 );
and ( n15528 , n8079 , n1134 );
xor ( n15529 , n15527 , n15528 );
xor ( n15530 , n15524 , n15529 );
xor ( n15531 , n15515 , n15530 );
and ( n15532 , n14714 , n14715 );
and ( n15533 , n14715 , n14717 );
and ( n15534 , n14714 , n14717 );
or ( n15535 , n15532 , n15533 , n15534 );
and ( n15536 , n6187 , n1882 );
and ( n15537 , n6569 , n1738 );
xor ( n15538 , n15536 , n15537 );
and ( n15539 , n6816 , n1551 );
xor ( n15540 , n15538 , n15539 );
xor ( n15541 , n15535 , n15540 );
and ( n15542 , n4959 , n2544 );
and ( n15543 , n5459 , n2298 );
xor ( n15544 , n15542 , n15543 );
and ( n15545 , n5819 , n2100 );
xor ( n15546 , n15544 , n15545 );
xor ( n15547 , n15541 , n15546 );
xor ( n15548 , n15531 , n15547 );
xor ( n15549 , n15511 , n15548 );
and ( n15550 , n14734 , n14740 );
and ( n15551 , n14740 , n14746 );
and ( n15552 , n14734 , n14746 );
or ( n15553 , n15550 , n15551 , n15552 );
and ( n15554 , n14772 , n14777 );
and ( n15555 , n14777 , n14783 );
and ( n15556 , n14772 , n14783 );
or ( n15557 , n15554 , n15555 , n15556 );
xor ( n15558 , n15553 , n15557 );
and ( n15559 , n14742 , n14743 );
and ( n15560 , n14743 , n14745 );
and ( n15561 , n14742 , n14745 );
or ( n15562 , n15559 , n15560 , n15561 );
and ( n15563 , n14773 , n14774 );
and ( n15564 , n14774 , n14776 );
and ( n15565 , n14773 , n14776 );
or ( n15566 , n15563 , n15564 , n15565 );
xor ( n15567 , n15562 , n15566 );
and ( n15568 , n4132 , n3271 );
and ( n15569 , n4438 , n2981 );
xor ( n15570 , n15568 , n15569 );
and ( n15571 , n4766 , n2739 );
xor ( n15572 , n15570 , n15571 );
xor ( n15573 , n15567 , n15572 );
xor ( n15574 , n15558 , n15573 );
xor ( n15575 , n15549 , n15574 );
xor ( n15576 , n15507 , n15575 );
xor ( n15577 , n15498 , n15576 );
and ( n15578 , n14807 , n14845 );
and ( n15579 , n14845 , n14872 );
and ( n15580 , n14807 , n14872 );
or ( n15581 , n15578 , n15579 , n15580 );
and ( n15582 , n14768 , n14784 );
and ( n15583 , n14784 , n14800 );
and ( n15584 , n14768 , n14800 );
or ( n15585 , n15582 , n15583 , n15584 );
and ( n15586 , n14850 , n14854 );
and ( n15587 , n14854 , n14871 );
and ( n15588 , n14850 , n14871 );
or ( n15589 , n15586 , n15587 , n15588 );
xor ( n15590 , n15585 , n15589 );
and ( n15591 , n14789 , n14793 );
and ( n15592 , n14793 , n14799 );
and ( n15593 , n14789 , n14799 );
or ( n15594 , n15591 , n15592 , n15593 );
and ( n15595 , n14779 , n14780 );
and ( n15596 , n14780 , n14782 );
and ( n15597 , n14779 , n14782 );
or ( n15598 , n15595 , n15596 , n15597 );
and ( n15599 , n3182 , n4102 );
and ( n15600 , n3545 , n3749 );
xor ( n15601 , n15599 , n15600 );
and ( n15602 , n3801 , n3495 );
xor ( n15603 , n15601 , n15602 );
xor ( n15604 , n15598 , n15603 );
and ( n15605 , n2462 , n5103 );
and ( n15606 , n2779 , n4730 );
xor ( n15607 , n15605 , n15606 );
and ( n15608 , n3024 , n4403 );
xor ( n15609 , n15607 , n15608 );
xor ( n15610 , n15604 , n15609 );
xor ( n15611 , n15594 , n15610 );
and ( n15612 , n14795 , n14796 );
and ( n15613 , n14796 , n14798 );
and ( n15614 , n14795 , n14798 );
or ( n15615 , n15612 , n15613 , n15614 );
and ( n15616 , n14860 , n14861 );
and ( n15617 , n14861 , n14863 );
and ( n15618 , n14860 , n14863 );
or ( n15619 , n15616 , n15617 , n15618 );
xor ( n15620 , n15615 , n15619 );
and ( n15621 , n1933 , n6132 );
and ( n15622 , n2120 , n5765 );
xor ( n15623 , n15621 , n15622 );
and ( n15624 , n2324 , n5408 );
xor ( n15625 , n15623 , n15624 );
xor ( n15626 , n15620 , n15625 );
xor ( n15627 , n15611 , n15626 );
xor ( n15628 , n15590 , n15627 );
xor ( n15629 , n15581 , n15628 );
and ( n15630 , n14811 , n14826 );
and ( n15631 , n14826 , n14844 );
and ( n15632 , n14811 , n14844 );
or ( n15633 , n15630 , n15631 , n15632 );
and ( n15634 , n14859 , n14864 );
and ( n15635 , n14864 , n14870 );
and ( n15636 , n14859 , n14870 );
or ( n15637 , n15634 , n15635 , n15636 );
and ( n15638 , n14815 , n14819 );
and ( n15639 , n14819 , n14825 );
and ( n15640 , n14815 , n14825 );
or ( n15641 , n15638 , n15639 , n15640 );
xor ( n15642 , n15637 , n15641 );
and ( n15643 , n14866 , n14867 );
and ( n15644 , n14867 , n14869 );
and ( n15645 , n14866 , n14869 );
or ( n15646 , n15643 , n15644 , n15645 );
and ( n15647 , n1383 , n7310 );
and ( n15648 , n1580 , n6971 );
xor ( n15649 , n15647 , n15648 );
and ( n15650 , n1694 , n6504 );
xor ( n15651 , n15649 , n15650 );
xor ( n15652 , n15646 , n15651 );
and ( n15653 , n1047 , n8669 );
and ( n15654 , n1164 , n8243 );
xor ( n15655 , n15653 , n15654 );
and ( n15656 , n1287 , n7662 );
xor ( n15657 , n15655 , n15656 );
xor ( n15658 , n15652 , n15657 );
xor ( n15659 , n15642 , n15658 );
xor ( n15660 , n15633 , n15659 );
and ( n15661 , n14831 , n14836 );
and ( n15662 , n14836 , n14843 );
and ( n15663 , n14831 , n14843 );
or ( n15664 , n15661 , n15662 , n15663 );
and ( n15665 , n14821 , n14822 );
and ( n15666 , n14822 , n14824 );
and ( n15667 , n14821 , n14824 );
or ( n15668 , n15665 , n15666 , n15667 );
and ( n15669 , n14832 , n14833 );
and ( n15670 , n14833 , n14835 );
and ( n15671 , n14832 , n14835 );
or ( n15672 , n15669 , n15670 , n15671 );
xor ( n15673 , n15668 , n15672 );
and ( n15674 , n783 , n10977 );
and ( n15675 , n856 , n10239 );
xor ( n15676 , n15674 , n15675 );
and ( n15677 , n925 , n9348 );
xor ( n15678 , n15676 , n15677 );
xor ( n15679 , n15673 , n15678 );
xor ( n15680 , n15664 , n15679 );
and ( n15681 , n14839 , n14840 );
and ( n15682 , n14840 , n14842 );
and ( n15683 , n14839 , n14842 );
or ( n15684 , n15681 , n15682 , n15683 );
and ( n15685 , n632 , n13256 );
and ( n15686 , n671 , n12531 );
xor ( n15687 , n15685 , n15686 );
and ( n15688 , n715 , n11718 );
xor ( n15689 , n15687 , n15688 );
xor ( n15690 , n15684 , n15689 );
buf ( n15691 , n425 );
and ( n15692 , n599 , n15691 );
and ( n15693 , n608 , n14838 );
xor ( n15694 , n15692 , n15693 );
and ( n15695 , n611 , n14044 );
xor ( n15696 , n15694 , n15695 );
xor ( n15697 , n15690 , n15696 );
xor ( n15698 , n15680 , n15697 );
xor ( n15699 , n15660 , n15698 );
xor ( n15700 , n15629 , n15699 );
xor ( n15701 , n15577 , n15700 );
xor ( n15702 , n15494 , n15701 );
and ( n15703 , n14674 , n14678 );
and ( n15704 , n14678 , n14749 );
and ( n15705 , n14674 , n14749 );
or ( n15706 , n15703 , n15704 , n15705 );
and ( n15707 , n14889 , n14925 );
and ( n15708 , n14925 , n14943 );
and ( n15709 , n14889 , n14943 );
or ( n15710 , n15707 , n15708 , n15709 );
xor ( n15711 , n15706 , n15710 );
and ( n15712 , n14893 , n14897 );
and ( n15713 , n14897 , n14924 );
and ( n15714 , n14893 , n14924 );
or ( n15715 , n15712 , n15713 , n15714 );
and ( n15716 , n14902 , n14906 );
and ( n15717 , n14906 , n14923 );
and ( n15718 , n14902 , n14923 );
or ( n15719 , n15716 , n15717 , n15718 );
and ( n15720 , n14687 , n14702 );
and ( n15721 , n14702 , n14719 );
and ( n15722 , n14687 , n14719 );
or ( n15723 , n15720 , n15721 , n15722 );
xor ( n15724 , n15719 , n15723 );
and ( n15725 , n14911 , n14916 );
and ( n15726 , n14916 , n14922 );
and ( n15727 , n14911 , n14922 );
or ( n15728 , n15725 , n15726 , n15727 );
and ( n15729 , n14691 , n14695 );
and ( n15730 , n14695 , n14701 );
and ( n15731 , n14691 , n14701 );
or ( n15732 , n15729 , n15730 , n15731 );
xor ( n15733 , n15728 , n15732 );
and ( n15734 , n14918 , n14919 );
and ( n15735 , n14919 , n14921 );
and ( n15736 , n14918 , n14921 );
or ( n15737 , n15734 , n15735 , n15736 );
and ( n15738 , n11015 , n771 );
and ( n15739 , n11769 , n719 );
xor ( n15740 , n15738 , n15739 );
and ( n15741 , n12320 , n663 );
xor ( n15742 , n15740 , n15741 );
xor ( n15743 , n15737 , n15742 );
and ( n15744 , n8718 , n1034 );
and ( n15745 , n9400 , n940 );
xor ( n15746 , n15744 , n15745 );
and ( n15747 , n10291 , n840 );
xor ( n15748 , n15746 , n15747 );
xor ( n15749 , n15743 , n15748 );
xor ( n15750 , n15733 , n15749 );
xor ( n15751 , n15724 , n15750 );
xor ( n15752 , n15715 , n15751 );
and ( n15753 , n14928 , n14941 );
and ( n15754 , n14932 , n14933 );
and ( n15755 , n14933 , n14940 );
and ( n15756 , n14932 , n14940 );
or ( n15757 , n15754 , n15755 , n15756 );
buf ( n15758 , n425 );
and ( n15759 , n15758 , n612 );
xor ( n15760 , n15757 , n15759 );
and ( n15761 , n14935 , n14936 );
and ( n15762 , n14936 , n14939 );
and ( n15763 , n14935 , n14939 );
or ( n15764 , n15761 , n15762 , n15763 );
and ( n15765 , n14912 , n14913 );
and ( n15766 , n14913 , n14915 );
and ( n15767 , n14912 , n14915 );
or ( n15768 , n15765 , n15766 , n15767 );
xor ( n15769 , n15764 , n15768 );
and ( n15770 , n13322 , n635 );
and ( n15771 , n14118 , n606 );
xor ( n15772 , n15770 , n15771 );
and ( n15773 , n14938 , n615 );
xor ( n15774 , n15772 , n15773 );
xor ( n15775 , n15769 , n15774 );
xor ( n15776 , n15760 , n15775 );
xor ( n15777 , n15753 , n15776 );
xor ( n15778 , n15752 , n15777 );
xor ( n15779 , n15711 , n15778 );
xor ( n15780 , n15702 , n15779 );
xor ( n15781 , n15490 , n15780 );
and ( n15782 , n14927 , n14942 );
and ( n15783 , n14880 , n14884 );
and ( n15784 , n14884 , n14944 );
and ( n15785 , n14880 , n14944 );
or ( n15786 , n15783 , n15784 , n15785 );
xor ( n15787 , n15782 , n15786 );
xor ( n15788 , n15781 , n15787 );
and ( n15789 , n14657 , n14661 );
and ( n15790 , n14661 , n14946 );
and ( n15791 , n14657 , n14946 );
or ( n15792 , n15789 , n15790 , n15791 );
xor ( n15793 , n15788 , n15792 );
and ( n15794 , n14947 , n14951 );
and ( n15795 , n14952 , n14955 );
or ( n15796 , n15794 , n15795 );
xor ( n15797 , n15793 , n15796 );
buf ( n15798 , n15797 );
buf ( n15799 , n15798 );
not ( n15800 , n15799 );
nor ( n15801 , n15800 , n8739 );
xor ( n15802 , n15486 , n15801 );
and ( n15803 , n14653 , n14960 );
and ( n15804 , n14961 , n14964 );
or ( n15805 , n15803 , n15804 );
xor ( n15806 , n15802 , n15805 );
buf ( n15807 , n15806 );
buf ( n15808 , n15807 );
not ( n15809 , n15808 );
buf ( n15810 , n544 );
not ( n15811 , n15810 );
nor ( n15812 , n15809 , n15811 );
xor ( n15813 , n15228 , n15812 );
xor ( n15814 , n14976 , n15225 );
nor ( n15815 , n14968 , n15811 );
and ( n15816 , n15814 , n15815 );
xor ( n15817 , n15814 , n15815 );
xor ( n15818 , n14980 , n15223 );
nor ( n15819 , n14147 , n15811 );
and ( n15820 , n15818 , n15819 );
xor ( n15821 , n15818 , n15819 );
xor ( n15822 , n14984 , n15221 );
nor ( n15823 , n13349 , n15811 );
and ( n15824 , n15822 , n15823 );
xor ( n15825 , n15822 , n15823 );
xor ( n15826 , n14988 , n15219 );
nor ( n15827 , n12564 , n15811 );
and ( n15828 , n15826 , n15827 );
xor ( n15829 , n15826 , n15827 );
xor ( n15830 , n14992 , n15217 );
nor ( n15831 , n11799 , n15811 );
and ( n15832 , n15830 , n15831 );
xor ( n15833 , n15830 , n15831 );
xor ( n15834 , n14996 , n15215 );
nor ( n15835 , n11050 , n15811 );
and ( n15836 , n15834 , n15835 );
xor ( n15837 , n15834 , n15835 );
xor ( n15838 , n15000 , n15213 );
nor ( n15839 , n10321 , n15811 );
and ( n15840 , n15838 , n15839 );
xor ( n15841 , n15838 , n15839 );
xor ( n15842 , n15004 , n15211 );
nor ( n15843 , n9429 , n15811 );
and ( n15844 , n15842 , n15843 );
xor ( n15845 , n15842 , n15843 );
xor ( n15846 , n15008 , n15209 );
nor ( n15847 , n8949 , n15811 );
and ( n15848 , n15846 , n15847 );
xor ( n15849 , n15846 , n15847 );
xor ( n15850 , n15012 , n15207 );
nor ( n15851 , n9437 , n15811 );
and ( n15852 , n15850 , n15851 );
xor ( n15853 , n15850 , n15851 );
xor ( n15854 , n15016 , n15205 );
nor ( n15855 , n9446 , n15811 );
and ( n15856 , n15854 , n15855 );
xor ( n15857 , n15854 , n15855 );
xor ( n15858 , n15020 , n15203 );
nor ( n15859 , n9455 , n15811 );
and ( n15860 , n15858 , n15859 );
xor ( n15861 , n15858 , n15859 );
xor ( n15862 , n15024 , n15201 );
nor ( n15863 , n9464 , n15811 );
and ( n15864 , n15862 , n15863 );
xor ( n15865 , n15862 , n15863 );
xor ( n15866 , n15028 , n15199 );
nor ( n15867 , n9473 , n15811 );
and ( n15868 , n15866 , n15867 );
xor ( n15869 , n15866 , n15867 );
xor ( n15870 , n15032 , n15197 );
nor ( n15871 , n9482 , n15811 );
and ( n15872 , n15870 , n15871 );
xor ( n15873 , n15870 , n15871 );
xor ( n15874 , n15036 , n15195 );
nor ( n15875 , n9491 , n15811 );
and ( n15876 , n15874 , n15875 );
xor ( n15877 , n15874 , n15875 );
xor ( n15878 , n15040 , n15193 );
nor ( n15879 , n9500 , n15811 );
and ( n15880 , n15878 , n15879 );
xor ( n15881 , n15878 , n15879 );
xor ( n15882 , n15044 , n15191 );
nor ( n15883 , n9509 , n15811 );
and ( n15884 , n15882 , n15883 );
xor ( n15885 , n15882 , n15883 );
xor ( n15886 , n15048 , n15189 );
nor ( n15887 , n9518 , n15811 );
and ( n15888 , n15886 , n15887 );
xor ( n15889 , n15886 , n15887 );
xor ( n15890 , n15052 , n15187 );
nor ( n15891 , n9527 , n15811 );
and ( n15892 , n15890 , n15891 );
xor ( n15893 , n15890 , n15891 );
xor ( n15894 , n15056 , n15185 );
nor ( n15895 , n9536 , n15811 );
and ( n15896 , n15894 , n15895 );
xor ( n15897 , n15894 , n15895 );
xor ( n15898 , n15060 , n15183 );
nor ( n15899 , n9545 , n15811 );
and ( n15900 , n15898 , n15899 );
xor ( n15901 , n15898 , n15899 );
xor ( n15902 , n15064 , n15181 );
nor ( n15903 , n9554 , n15811 );
and ( n15904 , n15902 , n15903 );
xor ( n15905 , n15902 , n15903 );
xor ( n15906 , n15068 , n15179 );
nor ( n15907 , n9563 , n15811 );
and ( n15908 , n15906 , n15907 );
xor ( n15909 , n15906 , n15907 );
xor ( n15910 , n15072 , n15177 );
nor ( n15911 , n9572 , n15811 );
and ( n15912 , n15910 , n15911 );
xor ( n15913 , n15910 , n15911 );
xor ( n15914 , n15076 , n15175 );
nor ( n15915 , n9581 , n15811 );
and ( n15916 , n15914 , n15915 );
xor ( n15917 , n15914 , n15915 );
xor ( n15918 , n15080 , n15173 );
nor ( n15919 , n9590 , n15811 );
and ( n15920 , n15918 , n15919 );
xor ( n15921 , n15918 , n15919 );
xor ( n15922 , n15084 , n15171 );
nor ( n15923 , n9599 , n15811 );
and ( n15924 , n15922 , n15923 );
xor ( n15925 , n15922 , n15923 );
xor ( n15926 , n15088 , n15169 );
nor ( n15927 , n9608 , n15811 );
and ( n15928 , n15926 , n15927 );
xor ( n15929 , n15926 , n15927 );
xor ( n15930 , n15092 , n15167 );
nor ( n15931 , n9617 , n15811 );
and ( n15932 , n15930 , n15931 );
xor ( n15933 , n15930 , n15931 );
xor ( n15934 , n15096 , n15165 );
nor ( n15935 , n9626 , n15811 );
and ( n15936 , n15934 , n15935 );
xor ( n15937 , n15934 , n15935 );
xor ( n15938 , n15100 , n15163 );
nor ( n15939 , n9635 , n15811 );
and ( n15940 , n15938 , n15939 );
xor ( n15941 , n15938 , n15939 );
xor ( n15942 , n15104 , n15161 );
nor ( n15943 , n9644 , n15811 );
and ( n15944 , n15942 , n15943 );
xor ( n15945 , n15942 , n15943 );
xor ( n15946 , n15108 , n15159 );
nor ( n15947 , n9653 , n15811 );
and ( n15948 , n15946 , n15947 );
xor ( n15949 , n15946 , n15947 );
xor ( n15950 , n15112 , n15157 );
nor ( n15951 , n9662 , n15811 );
and ( n15952 , n15950 , n15951 );
xor ( n15953 , n15950 , n15951 );
xor ( n15954 , n15116 , n15155 );
nor ( n15955 , n9671 , n15811 );
and ( n15956 , n15954 , n15955 );
xor ( n15957 , n15954 , n15955 );
xor ( n15958 , n15120 , n15153 );
nor ( n15959 , n9680 , n15811 );
and ( n15960 , n15958 , n15959 );
xor ( n15961 , n15958 , n15959 );
xor ( n15962 , n15124 , n15151 );
nor ( n15963 , n9689 , n15811 );
and ( n15964 , n15962 , n15963 );
xor ( n15965 , n15962 , n15963 );
xor ( n15966 , n15128 , n15149 );
nor ( n15967 , n9698 , n15811 );
and ( n15968 , n15966 , n15967 );
xor ( n15969 , n15966 , n15967 );
xor ( n15970 , n15132 , n15147 );
nor ( n15971 , n9707 , n15811 );
and ( n15972 , n15970 , n15971 );
xor ( n15973 , n15970 , n15971 );
xor ( n15974 , n15136 , n15145 );
nor ( n15975 , n9716 , n15811 );
and ( n15976 , n15974 , n15975 );
xor ( n15977 , n15974 , n15975 );
xor ( n15978 , n15140 , n15143 );
nor ( n15979 , n9725 , n15811 );
and ( n15980 , n15978 , n15979 );
xor ( n15981 , n15978 , n15979 );
xor ( n15982 , n15141 , n15142 );
nor ( n15983 , n9734 , n15811 );
and ( n15984 , n15982 , n15983 );
xor ( n15985 , n15982 , n15983 );
nor ( n15986 , n9752 , n14970 );
nor ( n15987 , n9743 , n15811 );
and ( n15988 , n15986 , n15987 );
and ( n15989 , n15985 , n15988 );
or ( n15990 , n15984 , n15989 );
and ( n15991 , n15981 , n15990 );
or ( n15992 , n15980 , n15991 );
and ( n15993 , n15977 , n15992 );
or ( n15994 , n15976 , n15993 );
and ( n15995 , n15973 , n15994 );
or ( n15996 , n15972 , n15995 );
and ( n15997 , n15969 , n15996 );
or ( n15998 , n15968 , n15997 );
and ( n15999 , n15965 , n15998 );
or ( n16000 , n15964 , n15999 );
and ( n16001 , n15961 , n16000 );
or ( n16002 , n15960 , n16001 );
and ( n16003 , n15957 , n16002 );
or ( n16004 , n15956 , n16003 );
and ( n16005 , n15953 , n16004 );
or ( n16006 , n15952 , n16005 );
and ( n16007 , n15949 , n16006 );
or ( n16008 , n15948 , n16007 );
and ( n16009 , n15945 , n16008 );
or ( n16010 , n15944 , n16009 );
and ( n16011 , n15941 , n16010 );
or ( n16012 , n15940 , n16011 );
and ( n16013 , n15937 , n16012 );
or ( n16014 , n15936 , n16013 );
and ( n16015 , n15933 , n16014 );
or ( n16016 , n15932 , n16015 );
and ( n16017 , n15929 , n16016 );
or ( n16018 , n15928 , n16017 );
and ( n16019 , n15925 , n16018 );
or ( n16020 , n15924 , n16019 );
and ( n16021 , n15921 , n16020 );
or ( n16022 , n15920 , n16021 );
and ( n16023 , n15917 , n16022 );
or ( n16024 , n15916 , n16023 );
and ( n16025 , n15913 , n16024 );
or ( n16026 , n15912 , n16025 );
and ( n16027 , n15909 , n16026 );
or ( n16028 , n15908 , n16027 );
and ( n16029 , n15905 , n16028 );
or ( n16030 , n15904 , n16029 );
and ( n16031 , n15901 , n16030 );
or ( n16032 , n15900 , n16031 );
and ( n16033 , n15897 , n16032 );
or ( n16034 , n15896 , n16033 );
and ( n16035 , n15893 , n16034 );
or ( n16036 , n15892 , n16035 );
and ( n16037 , n15889 , n16036 );
or ( n16038 , n15888 , n16037 );
and ( n16039 , n15885 , n16038 );
or ( n16040 , n15884 , n16039 );
and ( n16041 , n15881 , n16040 );
or ( n16042 , n15880 , n16041 );
and ( n16043 , n15877 , n16042 );
or ( n16044 , n15876 , n16043 );
and ( n16045 , n15873 , n16044 );
or ( n16046 , n15872 , n16045 );
and ( n16047 , n15869 , n16046 );
or ( n16048 , n15868 , n16047 );
and ( n16049 , n15865 , n16048 );
or ( n16050 , n15864 , n16049 );
and ( n16051 , n15861 , n16050 );
or ( n16052 , n15860 , n16051 );
and ( n16053 , n15857 , n16052 );
or ( n16054 , n15856 , n16053 );
and ( n16055 , n15853 , n16054 );
or ( n16056 , n15852 , n16055 );
and ( n16057 , n15849 , n16056 );
or ( n16058 , n15848 , n16057 );
and ( n16059 , n15845 , n16058 );
or ( n16060 , n15844 , n16059 );
and ( n16061 , n15841 , n16060 );
or ( n16062 , n15840 , n16061 );
and ( n16063 , n15837 , n16062 );
or ( n16064 , n15836 , n16063 );
and ( n16065 , n15833 , n16064 );
or ( n16066 , n15832 , n16065 );
and ( n16067 , n15829 , n16066 );
or ( n16068 , n15828 , n16067 );
and ( n16069 , n15825 , n16068 );
or ( n16070 , n15824 , n16069 );
and ( n16071 , n15821 , n16070 );
or ( n16072 , n15820 , n16071 );
and ( n16073 , n15817 , n16072 );
or ( n16074 , n15816 , n16073 );
xor ( n16075 , n15813 , n16074 );
buf ( n16076 , n488 );
not ( n16077 , n16076 );
nor ( n16078 , n601 , n16077 );
buf ( n16079 , n16078 );
nor ( n16080 , n622 , n14403 );
xor ( n16081 , n16079 , n16080 );
buf ( n16082 , n16081 );
nor ( n16083 , n646 , n13599 );
xor ( n16084 , n16082 , n16083 );
and ( n16085 , n15232 , n15233 );
buf ( n16086 , n16085 );
xor ( n16087 , n16084 , n16086 );
nor ( n16088 , n684 , n12808 );
xor ( n16089 , n16087 , n16088 );
and ( n16090 , n15235 , n15236 );
and ( n16091 , n15237 , n15239 );
or ( n16092 , n16090 , n16091 );
xor ( n16093 , n16089 , n16092 );
nor ( n16094 , n733 , n12037 );
xor ( n16095 , n16093 , n16094 );
and ( n16096 , n15240 , n15241 );
and ( n16097 , n15242 , n15245 );
or ( n16098 , n16096 , n16097 );
xor ( n16099 , n16095 , n16098 );
nor ( n16100 , n796 , n11282 );
xor ( n16101 , n16099 , n16100 );
and ( n16102 , n15246 , n15247 );
and ( n16103 , n15248 , n15251 );
or ( n16104 , n16102 , n16103 );
xor ( n16105 , n16101 , n16104 );
nor ( n16106 , n868 , n10547 );
xor ( n16107 , n16105 , n16106 );
and ( n16108 , n15252 , n15253 );
and ( n16109 , n15254 , n15257 );
or ( n16110 , n16108 , n16109 );
xor ( n16111 , n16107 , n16110 );
nor ( n16112 , n958 , n9829 );
xor ( n16113 , n16111 , n16112 );
and ( n16114 , n15258 , n15259 );
and ( n16115 , n15260 , n15263 );
or ( n16116 , n16114 , n16115 );
xor ( n16117 , n16113 , n16116 );
nor ( n16118 , n1062 , n8955 );
xor ( n16119 , n16117 , n16118 );
and ( n16120 , n15264 , n15265 );
and ( n16121 , n15266 , n15269 );
or ( n16122 , n16120 , n16121 );
xor ( n16123 , n16119 , n16122 );
nor ( n16124 , n1176 , n603 );
xor ( n16125 , n16123 , n16124 );
and ( n16126 , n15270 , n15271 );
and ( n16127 , n15272 , n15275 );
or ( n16128 , n16126 , n16127 );
xor ( n16129 , n16125 , n16128 );
nor ( n16130 , n1303 , n652 );
xor ( n16131 , n16129 , n16130 );
and ( n16132 , n15276 , n15277 );
and ( n16133 , n15278 , n15281 );
or ( n16134 , n16132 , n16133 );
xor ( n16135 , n16131 , n16134 );
nor ( n16136 , n1445 , n624 );
xor ( n16137 , n16135 , n16136 );
and ( n16138 , n15282 , n15283 );
and ( n16139 , n15284 , n15287 );
or ( n16140 , n16138 , n16139 );
xor ( n16141 , n16137 , n16140 );
nor ( n16142 , n1598 , n648 );
xor ( n16143 , n16141 , n16142 );
and ( n16144 , n15288 , n15289 );
and ( n16145 , n15290 , n15293 );
or ( n16146 , n16144 , n16145 );
xor ( n16147 , n16143 , n16146 );
nor ( n16148 , n1766 , n686 );
xor ( n16149 , n16147 , n16148 );
and ( n16150 , n15294 , n15295 );
and ( n16151 , n15296 , n15299 );
or ( n16152 , n16150 , n16151 );
xor ( n16153 , n16149 , n16152 );
nor ( n16154 , n1945 , n735 );
xor ( n16155 , n16153 , n16154 );
and ( n16156 , n15300 , n15301 );
and ( n16157 , n15302 , n15305 );
or ( n16158 , n16156 , n16157 );
xor ( n16159 , n16155 , n16158 );
nor ( n16160 , n2137 , n798 );
xor ( n16161 , n16159 , n16160 );
and ( n16162 , n15306 , n15307 );
and ( n16163 , n15308 , n15311 );
or ( n16164 , n16162 , n16163 );
xor ( n16165 , n16161 , n16164 );
nor ( n16166 , n2343 , n870 );
xor ( n16167 , n16165 , n16166 );
and ( n16168 , n15312 , n15313 );
and ( n16169 , n15314 , n15317 );
or ( n16170 , n16168 , n16169 );
xor ( n16171 , n16167 , n16170 );
nor ( n16172 , n2566 , n960 );
xor ( n16173 , n16171 , n16172 );
and ( n16174 , n15318 , n15319 );
and ( n16175 , n15320 , n15323 );
or ( n16176 , n16174 , n16175 );
xor ( n16177 , n16173 , n16176 );
nor ( n16178 , n2797 , n1064 );
xor ( n16179 , n16177 , n16178 );
and ( n16180 , n15324 , n15325 );
and ( n16181 , n15326 , n15329 );
or ( n16182 , n16180 , n16181 );
xor ( n16183 , n16179 , n16182 );
nor ( n16184 , n3043 , n1178 );
xor ( n16185 , n16183 , n16184 );
and ( n16186 , n15330 , n15331 );
and ( n16187 , n15332 , n15335 );
or ( n16188 , n16186 , n16187 );
xor ( n16189 , n16185 , n16188 );
nor ( n16190 , n3300 , n1305 );
xor ( n16191 , n16189 , n16190 );
and ( n16192 , n15336 , n15337 );
and ( n16193 , n15338 , n15341 );
or ( n16194 , n16192 , n16193 );
xor ( n16195 , n16191 , n16194 );
nor ( n16196 , n3570 , n1447 );
xor ( n16197 , n16195 , n16196 );
and ( n16198 , n15342 , n15343 );
and ( n16199 , n15344 , n15347 );
or ( n16200 , n16198 , n16199 );
xor ( n16201 , n16197 , n16200 );
nor ( n16202 , n3853 , n1600 );
xor ( n16203 , n16201 , n16202 );
and ( n16204 , n15348 , n15349 );
and ( n16205 , n15350 , n15353 );
or ( n16206 , n16204 , n16205 );
xor ( n16207 , n16203 , n16206 );
nor ( n16208 , n4151 , n1768 );
xor ( n16209 , n16207 , n16208 );
and ( n16210 , n15354 , n15355 );
and ( n16211 , n15356 , n15359 );
or ( n16212 , n16210 , n16211 );
xor ( n16213 , n16209 , n16212 );
nor ( n16214 , n4458 , n1947 );
xor ( n16215 , n16213 , n16214 );
and ( n16216 , n15360 , n15361 );
and ( n16217 , n15362 , n15365 );
or ( n16218 , n16216 , n16217 );
xor ( n16219 , n16215 , n16218 );
nor ( n16220 , n4786 , n2139 );
xor ( n16221 , n16219 , n16220 );
and ( n16222 , n15366 , n15367 );
and ( n16223 , n15368 , n15371 );
or ( n16224 , n16222 , n16223 );
xor ( n16225 , n16221 , n16224 );
nor ( n16226 , n5126 , n2345 );
xor ( n16227 , n16225 , n16226 );
and ( n16228 , n15372 , n15373 );
and ( n16229 , n15374 , n15377 );
or ( n16230 , n16228 , n16229 );
xor ( n16231 , n16227 , n16230 );
nor ( n16232 , n5477 , n2568 );
xor ( n16233 , n16231 , n16232 );
and ( n16234 , n15378 , n15379 );
and ( n16235 , n15380 , n15383 );
or ( n16236 , n16234 , n16235 );
xor ( n16237 , n16233 , n16236 );
nor ( n16238 , n5838 , n2799 );
xor ( n16239 , n16237 , n16238 );
and ( n16240 , n15384 , n15385 );
and ( n16241 , n15386 , n15389 );
or ( n16242 , n16240 , n16241 );
xor ( n16243 , n16239 , n16242 );
nor ( n16244 , n6212 , n3045 );
xor ( n16245 , n16243 , n16244 );
and ( n16246 , n15390 , n15391 );
and ( n16247 , n15392 , n15395 );
or ( n16248 , n16246 , n16247 );
xor ( n16249 , n16245 , n16248 );
nor ( n16250 , n6596 , n3302 );
xor ( n16251 , n16249 , n16250 );
and ( n16252 , n15396 , n15397 );
and ( n16253 , n15398 , n15401 );
or ( n16254 , n16252 , n16253 );
xor ( n16255 , n16251 , n16254 );
nor ( n16256 , n6997 , n3572 );
xor ( n16257 , n16255 , n16256 );
and ( n16258 , n15402 , n15403 );
and ( n16259 , n15404 , n15407 );
or ( n16260 , n16258 , n16259 );
xor ( n16261 , n16257 , n16260 );
nor ( n16262 , n7413 , n3855 );
xor ( n16263 , n16261 , n16262 );
and ( n16264 , n15408 , n15409 );
and ( n16265 , n15410 , n15413 );
or ( n16266 , n16264 , n16265 );
xor ( n16267 , n16263 , n16266 );
nor ( n16268 , n7841 , n4153 );
xor ( n16269 , n16267 , n16268 );
and ( n16270 , n15414 , n15415 );
and ( n16271 , n15416 , n15419 );
or ( n16272 , n16270 , n16271 );
xor ( n16273 , n16269 , n16272 );
nor ( n16274 , n8281 , n4460 );
xor ( n16275 , n16273 , n16274 );
and ( n16276 , n15420 , n15421 );
and ( n16277 , n15422 , n15425 );
or ( n16278 , n16276 , n16277 );
xor ( n16279 , n16275 , n16278 );
nor ( n16280 , n8737 , n4788 );
xor ( n16281 , n16279 , n16280 );
and ( n16282 , n15426 , n15427 );
and ( n16283 , n15428 , n15431 );
or ( n16284 , n16282 , n16283 );
xor ( n16285 , n16281 , n16284 );
nor ( n16286 , n9420 , n5128 );
xor ( n16287 , n16285 , n16286 );
and ( n16288 , n15432 , n15433 );
and ( n16289 , n15434 , n15437 );
or ( n16290 , n16288 , n16289 );
xor ( n16291 , n16287 , n16290 );
nor ( n16292 , n10312 , n5479 );
xor ( n16293 , n16291 , n16292 );
and ( n16294 , n15438 , n15439 );
and ( n16295 , n15440 , n15443 );
or ( n16296 , n16294 , n16295 );
xor ( n16297 , n16293 , n16296 );
nor ( n16298 , n11041 , n5840 );
xor ( n16299 , n16297 , n16298 );
and ( n16300 , n15444 , n15445 );
and ( n16301 , n15446 , n15449 );
or ( n16302 , n16300 , n16301 );
xor ( n16303 , n16299 , n16302 );
nor ( n16304 , n11790 , n6214 );
xor ( n16305 , n16303 , n16304 );
and ( n16306 , n15450 , n15451 );
and ( n16307 , n15452 , n15455 );
or ( n16308 , n16306 , n16307 );
xor ( n16309 , n16305 , n16308 );
nor ( n16310 , n12555 , n6598 );
xor ( n16311 , n16309 , n16310 );
and ( n16312 , n15456 , n15457 );
and ( n16313 , n15458 , n15461 );
or ( n16314 , n16312 , n16313 );
xor ( n16315 , n16311 , n16314 );
nor ( n16316 , n13340 , n6999 );
xor ( n16317 , n16315 , n16316 );
and ( n16318 , n15462 , n15463 );
and ( n16319 , n15464 , n15467 );
or ( n16320 , n16318 , n16319 );
xor ( n16321 , n16317 , n16320 );
nor ( n16322 , n14138 , n7415 );
xor ( n16323 , n16321 , n16322 );
and ( n16324 , n15468 , n15469 );
and ( n16325 , n15470 , n15473 );
or ( n16326 , n16324 , n16325 );
xor ( n16327 , n16323 , n16326 );
nor ( n16328 , n14959 , n7843 );
xor ( n16329 , n16327 , n16328 );
and ( n16330 , n15474 , n15475 );
and ( n16331 , n15476 , n15479 );
or ( n16332 , n16330 , n16331 );
xor ( n16333 , n16329 , n16332 );
nor ( n16334 , n15800 , n8283 );
xor ( n16335 , n16333 , n16334 );
and ( n16336 , n15480 , n15481 );
and ( n16337 , n15482 , n15485 );
or ( n16338 , n16336 , n16337 );
xor ( n16339 , n16335 , n16338 );
and ( n16340 , n15782 , n15786 );
and ( n16341 , n15490 , n15780 );
and ( n16342 , n15780 , n15787 );
and ( n16343 , n15490 , n15787 );
or ( n16344 , n16341 , n16342 , n16343 );
xor ( n16345 , n16340 , n16344 );
and ( n16346 , n15494 , n15701 );
and ( n16347 , n15701 , n15779 );
and ( n16348 , n15494 , n15779 );
or ( n16349 , n16346 , n16347 , n16348 );
and ( n16350 , n15498 , n15576 );
and ( n16351 , n15576 , n15700 );
and ( n16352 , n15498 , n15700 );
or ( n16353 , n16350 , n16351 , n16352 );
and ( n16354 , n15581 , n15628 );
and ( n16355 , n15628 , n15699 );
and ( n16356 , n15581 , n15699 );
or ( n16357 , n16354 , n16355 , n16356 );
and ( n16358 , n15511 , n15548 );
and ( n16359 , n15548 , n15574 );
and ( n16360 , n15511 , n15574 );
or ( n16361 , n16358 , n16359 , n16360 );
and ( n16362 , n15585 , n15589 );
and ( n16363 , n15589 , n15627 );
and ( n16364 , n15585 , n15627 );
or ( n16365 , n16362 , n16363 , n16364 );
xor ( n16366 , n16361 , n16365 );
and ( n16367 , n15553 , n15557 );
and ( n16368 , n15557 , n15573 );
and ( n16369 , n15553 , n15573 );
or ( n16370 , n16367 , n16368 , n16369 );
and ( n16371 , n15535 , n15540 );
and ( n16372 , n15540 , n15546 );
and ( n16373 , n15535 , n15546 );
or ( n16374 , n16371 , n16372 , n16373 );
and ( n16375 , n15525 , n15526 );
and ( n16376 , n15526 , n15528 );
and ( n16377 , n15525 , n15528 );
or ( n16378 , n16375 , n16376 , n16377 );
and ( n16379 , n15536 , n15537 );
and ( n16380 , n15537 , n15539 );
and ( n16381 , n15536 , n15539 );
or ( n16382 , n16379 , n16380 , n16381 );
xor ( n16383 , n16378 , n16382 );
and ( n16384 , n7385 , n1551 );
and ( n16385 , n7808 , n1424 );
xor ( n16386 , n16384 , n16385 );
and ( n16387 , n8079 , n1254 );
xor ( n16388 , n16386 , n16387 );
xor ( n16389 , n16383 , n16388 );
xor ( n16390 , n16374 , n16389 );
and ( n16391 , n15542 , n15543 );
and ( n16392 , n15543 , n15545 );
and ( n16393 , n15542 , n15545 );
or ( n16394 , n16391 , n16392 , n16393 );
and ( n16395 , n6187 , n2100 );
and ( n16396 , n6569 , n1882 );
xor ( n16397 , n16395 , n16396 );
and ( n16398 , n6816 , n1738 );
xor ( n16399 , n16397 , n16398 );
xor ( n16400 , n16394 , n16399 );
and ( n16401 , n4959 , n2739 );
and ( n16402 , n5459 , n2544 );
xor ( n16403 , n16401 , n16402 );
and ( n16404 , n5819 , n2298 );
xor ( n16405 , n16403 , n16404 );
xor ( n16406 , n16400 , n16405 );
xor ( n16407 , n16390 , n16406 );
xor ( n16408 , n16370 , n16407 );
and ( n16409 , n15562 , n15566 );
and ( n16410 , n15566 , n15572 );
and ( n16411 , n15562 , n15572 );
or ( n16412 , n16409 , n16410 , n16411 );
and ( n16413 , n15598 , n15603 );
and ( n16414 , n15603 , n15609 );
and ( n16415 , n15598 , n15609 );
or ( n16416 , n16413 , n16414 , n16415 );
xor ( n16417 , n16412 , n16416 );
and ( n16418 , n15568 , n15569 );
and ( n16419 , n15569 , n15571 );
and ( n16420 , n15568 , n15571 );
or ( n16421 , n16418 , n16419 , n16420 );
and ( n16422 , n15599 , n15600 );
and ( n16423 , n15600 , n15602 );
and ( n16424 , n15599 , n15602 );
or ( n16425 , n16422 , n16423 , n16424 );
xor ( n16426 , n16421 , n16425 );
and ( n16427 , n4132 , n3495 );
and ( n16428 , n4438 , n3271 );
xor ( n16429 , n16427 , n16428 );
and ( n16430 , n4766 , n2981 );
xor ( n16431 , n16429 , n16430 );
xor ( n16432 , n16426 , n16431 );
xor ( n16433 , n16417 , n16432 );
xor ( n16434 , n16408 , n16433 );
xor ( n16435 , n16366 , n16434 );
xor ( n16436 , n16357 , n16435 );
and ( n16437 , n15633 , n15659 );
and ( n16438 , n15659 , n15698 );
and ( n16439 , n15633 , n15698 );
or ( n16440 , n16437 , n16438 , n16439 );
and ( n16441 , n15594 , n15610 );
and ( n16442 , n15610 , n15626 );
and ( n16443 , n15594 , n15626 );
or ( n16444 , n16441 , n16442 , n16443 );
and ( n16445 , n15637 , n15641 );
and ( n16446 , n15641 , n15658 );
and ( n16447 , n15637 , n15658 );
or ( n16448 , n16445 , n16446 , n16447 );
xor ( n16449 , n16444 , n16448 );
and ( n16450 , n15615 , n15619 );
and ( n16451 , n15619 , n15625 );
and ( n16452 , n15615 , n15625 );
or ( n16453 , n16450 , n16451 , n16452 );
and ( n16454 , n15605 , n15606 );
and ( n16455 , n15606 , n15608 );
and ( n16456 , n15605 , n15608 );
or ( n16457 , n16454 , n16455 , n16456 );
and ( n16458 , n3182 , n4403 );
and ( n16459 , n3545 , n4102 );
xor ( n16460 , n16458 , n16459 );
buf ( n16461 , n3801 );
xor ( n16462 , n16460 , n16461 );
xor ( n16463 , n16457 , n16462 );
and ( n16464 , n2462 , n5408 );
and ( n16465 , n2779 , n5103 );
xor ( n16466 , n16464 , n16465 );
and ( n16467 , n3024 , n4730 );
xor ( n16468 , n16466 , n16467 );
xor ( n16469 , n16463 , n16468 );
xor ( n16470 , n16453 , n16469 );
and ( n16471 , n15621 , n15622 );
and ( n16472 , n15622 , n15624 );
and ( n16473 , n15621 , n15624 );
or ( n16474 , n16471 , n16472 , n16473 );
and ( n16475 , n15647 , n15648 );
and ( n16476 , n15648 , n15650 );
and ( n16477 , n15647 , n15650 );
or ( n16478 , n16475 , n16476 , n16477 );
xor ( n16479 , n16474 , n16478 );
and ( n16480 , n1933 , n6504 );
and ( n16481 , n2120 , n6132 );
xor ( n16482 , n16480 , n16481 );
and ( n16483 , n2324 , n5765 );
xor ( n16484 , n16482 , n16483 );
xor ( n16485 , n16479 , n16484 );
xor ( n16486 , n16470 , n16485 );
xor ( n16487 , n16449 , n16486 );
xor ( n16488 , n16440 , n16487 );
and ( n16489 , n15664 , n15679 );
and ( n16490 , n15679 , n15697 );
and ( n16491 , n15664 , n15697 );
or ( n16492 , n16489 , n16490 , n16491 );
and ( n16493 , n15646 , n15651 );
and ( n16494 , n15651 , n15657 );
and ( n16495 , n15646 , n15657 );
or ( n16496 , n16493 , n16494 , n16495 );
and ( n16497 , n15668 , n15672 );
and ( n16498 , n15672 , n15678 );
and ( n16499 , n15668 , n15678 );
or ( n16500 , n16497 , n16498 , n16499 );
xor ( n16501 , n16496 , n16500 );
and ( n16502 , n15653 , n15654 );
and ( n16503 , n15654 , n15656 );
and ( n16504 , n15653 , n15656 );
or ( n16505 , n16502 , n16503 , n16504 );
and ( n16506 , n1383 , n7662 );
and ( n16507 , n1580 , n7310 );
xor ( n16508 , n16506 , n16507 );
and ( n16509 , n1694 , n6971 );
xor ( n16510 , n16508 , n16509 );
xor ( n16511 , n16505 , n16510 );
and ( n16512 , n1047 , n9348 );
and ( n16513 , n1164 , n8669 );
xor ( n16514 , n16512 , n16513 );
and ( n16515 , n1287 , n8243 );
xor ( n16516 , n16514 , n16515 );
xor ( n16517 , n16511 , n16516 );
xor ( n16518 , n16501 , n16517 );
xor ( n16519 , n16492 , n16518 );
and ( n16520 , n15684 , n15689 );
and ( n16521 , n15689 , n15696 );
and ( n16522 , n15684 , n15696 );
or ( n16523 , n16520 , n16521 , n16522 );
and ( n16524 , n15674 , n15675 );
and ( n16525 , n15675 , n15677 );
and ( n16526 , n15674 , n15677 );
or ( n16527 , n16524 , n16525 , n16526 );
and ( n16528 , n15685 , n15686 );
and ( n16529 , n15686 , n15688 );
and ( n16530 , n15685 , n15688 );
or ( n16531 , n16528 , n16529 , n16530 );
xor ( n16532 , n16527 , n16531 );
and ( n16533 , n783 , n11718 );
and ( n16534 , n856 , n10977 );
xor ( n16535 , n16533 , n16534 );
and ( n16536 , n925 , n10239 );
xor ( n16537 , n16535 , n16536 );
xor ( n16538 , n16532 , n16537 );
xor ( n16539 , n16523 , n16538 );
and ( n16540 , n15692 , n15693 );
and ( n16541 , n15693 , n15695 );
and ( n16542 , n15692 , n15695 );
or ( n16543 , n16540 , n16541 , n16542 );
and ( n16544 , n632 , n14044 );
and ( n16545 , n671 , n13256 );
xor ( n16546 , n16544 , n16545 );
and ( n16547 , n715 , n12531 );
xor ( n16548 , n16546 , n16547 );
xor ( n16549 , n16543 , n16548 );
buf ( n16550 , n424 );
and ( n16551 , n599 , n16550 );
and ( n16552 , n608 , n15691 );
xor ( n16553 , n16551 , n16552 );
and ( n16554 , n611 , n14838 );
xor ( n16555 , n16553 , n16554 );
xor ( n16556 , n16549 , n16555 );
xor ( n16557 , n16539 , n16556 );
xor ( n16558 , n16519 , n16557 );
xor ( n16559 , n16488 , n16558 );
xor ( n16560 , n16436 , n16559 );
xor ( n16561 , n16353 , n16560 );
and ( n16562 , n15502 , n15506 );
and ( n16563 , n15506 , n15575 );
and ( n16564 , n15502 , n15575 );
or ( n16565 , n16562 , n16563 , n16564 );
and ( n16566 , n15715 , n15751 );
and ( n16567 , n15751 , n15777 );
and ( n16568 , n15715 , n15777 );
or ( n16569 , n16566 , n16567 , n16568 );
xor ( n16570 , n16565 , n16569 );
and ( n16571 , n15719 , n15723 );
and ( n16572 , n15723 , n15750 );
and ( n16573 , n15719 , n15750 );
or ( n16574 , n16571 , n16572 , n16573 );
and ( n16575 , n15728 , n15732 );
and ( n16576 , n15732 , n15749 );
and ( n16577 , n15728 , n15749 );
or ( n16578 , n16575 , n16576 , n16577 );
and ( n16579 , n15515 , n15530 );
and ( n16580 , n15530 , n15547 );
and ( n16581 , n15515 , n15547 );
or ( n16582 , n16579 , n16580 , n16581 );
xor ( n16583 , n16578 , n16582 );
and ( n16584 , n15737 , n15742 );
and ( n16585 , n15742 , n15748 );
and ( n16586 , n15737 , n15748 );
or ( n16587 , n16584 , n16585 , n16586 );
and ( n16588 , n15519 , n15523 );
and ( n16589 , n15523 , n15529 );
and ( n16590 , n15519 , n15529 );
or ( n16591 , n16588 , n16589 , n16590 );
xor ( n16592 , n16587 , n16591 );
and ( n16593 , n15744 , n15745 );
and ( n16594 , n15745 , n15747 );
and ( n16595 , n15744 , n15747 );
or ( n16596 , n16593 , n16594 , n16595 );
and ( n16597 , n11015 , n840 );
and ( n16598 , n11769 , n771 );
xor ( n16599 , n16597 , n16598 );
and ( n16600 , n12320 , n719 );
xor ( n16601 , n16599 , n16600 );
xor ( n16602 , n16596 , n16601 );
and ( n16603 , n8718 , n1134 );
and ( n16604 , n9400 , n1034 );
xor ( n16605 , n16603 , n16604 );
and ( n16606 , n10291 , n940 );
xor ( n16607 , n16605 , n16606 );
xor ( n16608 , n16602 , n16607 );
xor ( n16609 , n16592 , n16608 );
xor ( n16610 , n16583 , n16609 );
xor ( n16611 , n16574 , n16610 );
and ( n16612 , n15757 , n15759 );
and ( n16613 , n15759 , n15775 );
and ( n16614 , n15757 , n15775 );
or ( n16615 , n16612 , n16613 , n16614 );
and ( n16616 , n15764 , n15768 );
and ( n16617 , n15768 , n15774 );
and ( n16618 , n15764 , n15774 );
or ( n16619 , n16616 , n16617 , n16618 );
and ( n16620 , n15770 , n15771 );
and ( n16621 , n15771 , n15773 );
and ( n16622 , n15770 , n15773 );
or ( n16623 , n16620 , n16621 , n16622 );
and ( n16624 , n15738 , n15739 );
and ( n16625 , n15739 , n15741 );
and ( n16626 , n15738 , n15741 );
or ( n16627 , n16624 , n16625 , n16626 );
xor ( n16628 , n16623 , n16627 );
and ( n16629 , n13322 , n663 );
and ( n16630 , n14118 , n635 );
xor ( n16631 , n16629 , n16630 );
and ( n16632 , n14938 , n606 );
xor ( n16633 , n16631 , n16632 );
xor ( n16634 , n16628 , n16633 );
xor ( n16635 , n16619 , n16634 );
and ( n16636 , n15758 , n615 );
buf ( n16637 , n424 );
and ( n16638 , n16637 , n612 );
xor ( n16639 , n16636 , n16638 );
xor ( n16640 , n16635 , n16639 );
xor ( n16641 , n16615 , n16640 );
xor ( n16642 , n16611 , n16641 );
xor ( n16643 , n16570 , n16642 );
xor ( n16644 , n16561 , n16643 );
xor ( n16645 , n16349 , n16644 );
and ( n16646 , n15753 , n15776 );
and ( n16647 , n15706 , n15710 );
and ( n16648 , n15710 , n15778 );
and ( n16649 , n15706 , n15778 );
or ( n16650 , n16647 , n16648 , n16649 );
xor ( n16651 , n16646 , n16650 );
xor ( n16652 , n16645 , n16651 );
xor ( n16653 , n16345 , n16652 );
and ( n16654 , n15788 , n15792 );
and ( n16655 , n15793 , n15796 );
or ( n16656 , n16654 , n16655 );
xor ( n16657 , n16653 , n16656 );
buf ( n16658 , n16657 );
buf ( n16659 , n16658 );
not ( n16660 , n16659 );
nor ( n16661 , n16660 , n8739 );
xor ( n16662 , n16339 , n16661 );
and ( n16663 , n15486 , n15801 );
and ( n16664 , n15802 , n15805 );
or ( n16665 , n16663 , n16664 );
xor ( n16666 , n16662 , n16665 );
buf ( n16667 , n16666 );
buf ( n16668 , n16667 );
not ( n16669 , n16668 );
buf ( n16670 , n545 );
not ( n16671 , n16670 );
nor ( n16672 , n16669 , n16671 );
xor ( n16673 , n16075 , n16672 );
xor ( n16674 , n15817 , n16072 );
nor ( n16675 , n15809 , n16671 );
and ( n16676 , n16674 , n16675 );
xor ( n16677 , n16674 , n16675 );
xor ( n16678 , n15821 , n16070 );
nor ( n16679 , n14968 , n16671 );
and ( n16680 , n16678 , n16679 );
xor ( n16681 , n16678 , n16679 );
xor ( n16682 , n15825 , n16068 );
nor ( n16683 , n14147 , n16671 );
and ( n16684 , n16682 , n16683 );
xor ( n16685 , n16682 , n16683 );
xor ( n16686 , n15829 , n16066 );
nor ( n16687 , n13349 , n16671 );
and ( n16688 , n16686 , n16687 );
xor ( n16689 , n16686 , n16687 );
xor ( n16690 , n15833 , n16064 );
nor ( n16691 , n12564 , n16671 );
and ( n16692 , n16690 , n16691 );
xor ( n16693 , n16690 , n16691 );
xor ( n16694 , n15837 , n16062 );
nor ( n16695 , n11799 , n16671 );
and ( n16696 , n16694 , n16695 );
xor ( n16697 , n16694 , n16695 );
xor ( n16698 , n15841 , n16060 );
nor ( n16699 , n11050 , n16671 );
and ( n16700 , n16698 , n16699 );
xor ( n16701 , n16698 , n16699 );
xor ( n16702 , n15845 , n16058 );
nor ( n16703 , n10321 , n16671 );
and ( n16704 , n16702 , n16703 );
xor ( n16705 , n16702 , n16703 );
xor ( n16706 , n15849 , n16056 );
nor ( n16707 , n9429 , n16671 );
and ( n16708 , n16706 , n16707 );
xor ( n16709 , n16706 , n16707 );
xor ( n16710 , n15853 , n16054 );
nor ( n16711 , n8949 , n16671 );
and ( n16712 , n16710 , n16711 );
xor ( n16713 , n16710 , n16711 );
xor ( n16714 , n15857 , n16052 );
nor ( n16715 , n9437 , n16671 );
and ( n16716 , n16714 , n16715 );
xor ( n16717 , n16714 , n16715 );
xor ( n16718 , n15861 , n16050 );
nor ( n16719 , n9446 , n16671 );
and ( n16720 , n16718 , n16719 );
xor ( n16721 , n16718 , n16719 );
xor ( n16722 , n15865 , n16048 );
nor ( n16723 , n9455 , n16671 );
and ( n16724 , n16722 , n16723 );
xor ( n16725 , n16722 , n16723 );
xor ( n16726 , n15869 , n16046 );
nor ( n16727 , n9464 , n16671 );
and ( n16728 , n16726 , n16727 );
xor ( n16729 , n16726 , n16727 );
xor ( n16730 , n15873 , n16044 );
nor ( n16731 , n9473 , n16671 );
and ( n16732 , n16730 , n16731 );
xor ( n16733 , n16730 , n16731 );
xor ( n16734 , n15877 , n16042 );
nor ( n16735 , n9482 , n16671 );
and ( n16736 , n16734 , n16735 );
xor ( n16737 , n16734 , n16735 );
xor ( n16738 , n15881 , n16040 );
nor ( n16739 , n9491 , n16671 );
and ( n16740 , n16738 , n16739 );
xor ( n16741 , n16738 , n16739 );
xor ( n16742 , n15885 , n16038 );
nor ( n16743 , n9500 , n16671 );
and ( n16744 , n16742 , n16743 );
xor ( n16745 , n16742 , n16743 );
xor ( n16746 , n15889 , n16036 );
nor ( n16747 , n9509 , n16671 );
and ( n16748 , n16746 , n16747 );
xor ( n16749 , n16746 , n16747 );
xor ( n16750 , n15893 , n16034 );
nor ( n16751 , n9518 , n16671 );
and ( n16752 , n16750 , n16751 );
xor ( n16753 , n16750 , n16751 );
xor ( n16754 , n15897 , n16032 );
nor ( n16755 , n9527 , n16671 );
and ( n16756 , n16754 , n16755 );
xor ( n16757 , n16754 , n16755 );
xor ( n16758 , n15901 , n16030 );
nor ( n16759 , n9536 , n16671 );
and ( n16760 , n16758 , n16759 );
xor ( n16761 , n16758 , n16759 );
xor ( n16762 , n15905 , n16028 );
nor ( n16763 , n9545 , n16671 );
and ( n16764 , n16762 , n16763 );
xor ( n16765 , n16762 , n16763 );
xor ( n16766 , n15909 , n16026 );
nor ( n16767 , n9554 , n16671 );
and ( n16768 , n16766 , n16767 );
xor ( n16769 , n16766 , n16767 );
xor ( n16770 , n15913 , n16024 );
nor ( n16771 , n9563 , n16671 );
and ( n16772 , n16770 , n16771 );
xor ( n16773 , n16770 , n16771 );
xor ( n16774 , n15917 , n16022 );
nor ( n16775 , n9572 , n16671 );
and ( n16776 , n16774 , n16775 );
xor ( n16777 , n16774 , n16775 );
xor ( n16778 , n15921 , n16020 );
nor ( n16779 , n9581 , n16671 );
and ( n16780 , n16778 , n16779 );
xor ( n16781 , n16778 , n16779 );
xor ( n16782 , n15925 , n16018 );
nor ( n16783 , n9590 , n16671 );
and ( n16784 , n16782 , n16783 );
xor ( n16785 , n16782 , n16783 );
xor ( n16786 , n15929 , n16016 );
nor ( n16787 , n9599 , n16671 );
and ( n16788 , n16786 , n16787 );
xor ( n16789 , n16786 , n16787 );
xor ( n16790 , n15933 , n16014 );
nor ( n16791 , n9608 , n16671 );
and ( n16792 , n16790 , n16791 );
xor ( n16793 , n16790 , n16791 );
xor ( n16794 , n15937 , n16012 );
nor ( n16795 , n9617 , n16671 );
and ( n16796 , n16794 , n16795 );
xor ( n16797 , n16794 , n16795 );
xor ( n16798 , n15941 , n16010 );
nor ( n16799 , n9626 , n16671 );
and ( n16800 , n16798 , n16799 );
xor ( n16801 , n16798 , n16799 );
xor ( n16802 , n15945 , n16008 );
nor ( n16803 , n9635 , n16671 );
and ( n16804 , n16802 , n16803 );
xor ( n16805 , n16802 , n16803 );
xor ( n16806 , n15949 , n16006 );
nor ( n16807 , n9644 , n16671 );
and ( n16808 , n16806 , n16807 );
xor ( n16809 , n16806 , n16807 );
xor ( n16810 , n15953 , n16004 );
nor ( n16811 , n9653 , n16671 );
and ( n16812 , n16810 , n16811 );
xor ( n16813 , n16810 , n16811 );
xor ( n16814 , n15957 , n16002 );
nor ( n16815 , n9662 , n16671 );
and ( n16816 , n16814 , n16815 );
xor ( n16817 , n16814 , n16815 );
xor ( n16818 , n15961 , n16000 );
nor ( n16819 , n9671 , n16671 );
and ( n16820 , n16818 , n16819 );
xor ( n16821 , n16818 , n16819 );
xor ( n16822 , n15965 , n15998 );
nor ( n16823 , n9680 , n16671 );
and ( n16824 , n16822 , n16823 );
xor ( n16825 , n16822 , n16823 );
xor ( n16826 , n15969 , n15996 );
nor ( n16827 , n9689 , n16671 );
and ( n16828 , n16826 , n16827 );
xor ( n16829 , n16826 , n16827 );
xor ( n16830 , n15973 , n15994 );
nor ( n16831 , n9698 , n16671 );
and ( n16832 , n16830 , n16831 );
xor ( n16833 , n16830 , n16831 );
xor ( n16834 , n15977 , n15992 );
nor ( n16835 , n9707 , n16671 );
and ( n16836 , n16834 , n16835 );
xor ( n16837 , n16834 , n16835 );
xor ( n16838 , n15981 , n15990 );
nor ( n16839 , n9716 , n16671 );
and ( n16840 , n16838 , n16839 );
xor ( n16841 , n16838 , n16839 );
xor ( n16842 , n15985 , n15988 );
nor ( n16843 , n9725 , n16671 );
and ( n16844 , n16842 , n16843 );
xor ( n16845 , n16842 , n16843 );
xor ( n16846 , n15986 , n15987 );
nor ( n16847 , n9734 , n16671 );
and ( n16848 , n16846 , n16847 );
xor ( n16849 , n16846 , n16847 );
nor ( n16850 , n9752 , n15811 );
nor ( n16851 , n9743 , n16671 );
and ( n16852 , n16850 , n16851 );
and ( n16853 , n16849 , n16852 );
or ( n16854 , n16848 , n16853 );
and ( n16855 , n16845 , n16854 );
or ( n16856 , n16844 , n16855 );
and ( n16857 , n16841 , n16856 );
or ( n16858 , n16840 , n16857 );
and ( n16859 , n16837 , n16858 );
or ( n16860 , n16836 , n16859 );
and ( n16861 , n16833 , n16860 );
or ( n16862 , n16832 , n16861 );
and ( n16863 , n16829 , n16862 );
or ( n16864 , n16828 , n16863 );
and ( n16865 , n16825 , n16864 );
or ( n16866 , n16824 , n16865 );
and ( n16867 , n16821 , n16866 );
or ( n16868 , n16820 , n16867 );
and ( n16869 , n16817 , n16868 );
or ( n16870 , n16816 , n16869 );
and ( n16871 , n16813 , n16870 );
or ( n16872 , n16812 , n16871 );
and ( n16873 , n16809 , n16872 );
or ( n16874 , n16808 , n16873 );
and ( n16875 , n16805 , n16874 );
or ( n16876 , n16804 , n16875 );
and ( n16877 , n16801 , n16876 );
or ( n16878 , n16800 , n16877 );
and ( n16879 , n16797 , n16878 );
or ( n16880 , n16796 , n16879 );
and ( n16881 , n16793 , n16880 );
or ( n16882 , n16792 , n16881 );
and ( n16883 , n16789 , n16882 );
or ( n16884 , n16788 , n16883 );
and ( n16885 , n16785 , n16884 );
or ( n16886 , n16784 , n16885 );
and ( n16887 , n16781 , n16886 );
or ( n16888 , n16780 , n16887 );
and ( n16889 , n16777 , n16888 );
or ( n16890 , n16776 , n16889 );
and ( n16891 , n16773 , n16890 );
or ( n16892 , n16772 , n16891 );
and ( n16893 , n16769 , n16892 );
or ( n16894 , n16768 , n16893 );
and ( n16895 , n16765 , n16894 );
or ( n16896 , n16764 , n16895 );
and ( n16897 , n16761 , n16896 );
or ( n16898 , n16760 , n16897 );
and ( n16899 , n16757 , n16898 );
or ( n16900 , n16756 , n16899 );
and ( n16901 , n16753 , n16900 );
or ( n16902 , n16752 , n16901 );
and ( n16903 , n16749 , n16902 );
or ( n16904 , n16748 , n16903 );
and ( n16905 , n16745 , n16904 );
or ( n16906 , n16744 , n16905 );
and ( n16907 , n16741 , n16906 );
or ( n16908 , n16740 , n16907 );
and ( n16909 , n16737 , n16908 );
or ( n16910 , n16736 , n16909 );
and ( n16911 , n16733 , n16910 );
or ( n16912 , n16732 , n16911 );
and ( n16913 , n16729 , n16912 );
or ( n16914 , n16728 , n16913 );
and ( n16915 , n16725 , n16914 );
or ( n16916 , n16724 , n16915 );
and ( n16917 , n16721 , n16916 );
or ( n16918 , n16720 , n16917 );
and ( n16919 , n16717 , n16918 );
or ( n16920 , n16716 , n16919 );
and ( n16921 , n16713 , n16920 );
or ( n16922 , n16712 , n16921 );
and ( n16923 , n16709 , n16922 );
or ( n16924 , n16708 , n16923 );
and ( n16925 , n16705 , n16924 );
or ( n16926 , n16704 , n16925 );
and ( n16927 , n16701 , n16926 );
or ( n16928 , n16700 , n16927 );
and ( n16929 , n16697 , n16928 );
or ( n16930 , n16696 , n16929 );
and ( n16931 , n16693 , n16930 );
or ( n16932 , n16692 , n16931 );
and ( n16933 , n16689 , n16932 );
or ( n16934 , n16688 , n16933 );
and ( n16935 , n16685 , n16934 );
or ( n16936 , n16684 , n16935 );
and ( n16937 , n16681 , n16936 );
or ( n16938 , n16680 , n16937 );
and ( n16939 , n16677 , n16938 );
or ( n16940 , n16676 , n16939 );
xor ( n16941 , n16673 , n16940 );
buf ( n16942 , n487 );
not ( n16943 , n16942 );
nor ( n16944 , n601 , n16943 );
buf ( n16945 , n16944 );
nor ( n16946 , n622 , n15230 );
xor ( n16947 , n16945 , n16946 );
buf ( n16948 , n16947 );
nor ( n16949 , n646 , n14403 );
xor ( n16950 , n16948 , n16949 );
and ( n16951 , n16079 , n16080 );
buf ( n16952 , n16951 );
xor ( n16953 , n16950 , n16952 );
nor ( n16954 , n684 , n13599 );
xor ( n16955 , n16953 , n16954 );
and ( n16956 , n16082 , n16083 );
and ( n16957 , n16084 , n16086 );
or ( n16958 , n16956 , n16957 );
xor ( n16959 , n16955 , n16958 );
nor ( n16960 , n733 , n12808 );
xor ( n16961 , n16959 , n16960 );
and ( n16962 , n16087 , n16088 );
and ( n16963 , n16089 , n16092 );
or ( n16964 , n16962 , n16963 );
xor ( n16965 , n16961 , n16964 );
nor ( n16966 , n796 , n12037 );
xor ( n16967 , n16965 , n16966 );
and ( n16968 , n16093 , n16094 );
and ( n16969 , n16095 , n16098 );
or ( n16970 , n16968 , n16969 );
xor ( n16971 , n16967 , n16970 );
nor ( n16972 , n868 , n11282 );
xor ( n16973 , n16971 , n16972 );
and ( n16974 , n16099 , n16100 );
and ( n16975 , n16101 , n16104 );
or ( n16976 , n16974 , n16975 );
xor ( n16977 , n16973 , n16976 );
nor ( n16978 , n958 , n10547 );
xor ( n16979 , n16977 , n16978 );
and ( n16980 , n16105 , n16106 );
and ( n16981 , n16107 , n16110 );
or ( n16982 , n16980 , n16981 );
xor ( n16983 , n16979 , n16982 );
nor ( n16984 , n1062 , n9829 );
xor ( n16985 , n16983 , n16984 );
and ( n16986 , n16111 , n16112 );
and ( n16987 , n16113 , n16116 );
or ( n16988 , n16986 , n16987 );
xor ( n16989 , n16985 , n16988 );
nor ( n16990 , n1176 , n8955 );
xor ( n16991 , n16989 , n16990 );
and ( n16992 , n16117 , n16118 );
and ( n16993 , n16119 , n16122 );
or ( n16994 , n16992 , n16993 );
xor ( n16995 , n16991 , n16994 );
nor ( n16996 , n1303 , n603 );
xor ( n16997 , n16995 , n16996 );
and ( n16998 , n16123 , n16124 );
and ( n16999 , n16125 , n16128 );
or ( n17000 , n16998 , n16999 );
xor ( n17001 , n16997 , n17000 );
nor ( n17002 , n1445 , n652 );
xor ( n17003 , n17001 , n17002 );
and ( n17004 , n16129 , n16130 );
and ( n17005 , n16131 , n16134 );
or ( n17006 , n17004 , n17005 );
xor ( n17007 , n17003 , n17006 );
nor ( n17008 , n1598 , n624 );
xor ( n17009 , n17007 , n17008 );
and ( n17010 , n16135 , n16136 );
and ( n17011 , n16137 , n16140 );
or ( n17012 , n17010 , n17011 );
xor ( n17013 , n17009 , n17012 );
nor ( n17014 , n1766 , n648 );
xor ( n17015 , n17013 , n17014 );
and ( n17016 , n16141 , n16142 );
and ( n17017 , n16143 , n16146 );
or ( n17018 , n17016 , n17017 );
xor ( n17019 , n17015 , n17018 );
nor ( n17020 , n1945 , n686 );
xor ( n17021 , n17019 , n17020 );
and ( n17022 , n16147 , n16148 );
and ( n17023 , n16149 , n16152 );
or ( n17024 , n17022 , n17023 );
xor ( n17025 , n17021 , n17024 );
nor ( n17026 , n2137 , n735 );
xor ( n17027 , n17025 , n17026 );
and ( n17028 , n16153 , n16154 );
and ( n17029 , n16155 , n16158 );
or ( n17030 , n17028 , n17029 );
xor ( n17031 , n17027 , n17030 );
nor ( n17032 , n2343 , n798 );
xor ( n17033 , n17031 , n17032 );
and ( n17034 , n16159 , n16160 );
and ( n17035 , n16161 , n16164 );
or ( n17036 , n17034 , n17035 );
xor ( n17037 , n17033 , n17036 );
nor ( n17038 , n2566 , n870 );
xor ( n17039 , n17037 , n17038 );
and ( n17040 , n16165 , n16166 );
and ( n17041 , n16167 , n16170 );
or ( n17042 , n17040 , n17041 );
xor ( n17043 , n17039 , n17042 );
nor ( n17044 , n2797 , n960 );
xor ( n17045 , n17043 , n17044 );
and ( n17046 , n16171 , n16172 );
and ( n17047 , n16173 , n16176 );
or ( n17048 , n17046 , n17047 );
xor ( n17049 , n17045 , n17048 );
nor ( n17050 , n3043 , n1064 );
xor ( n17051 , n17049 , n17050 );
and ( n17052 , n16177 , n16178 );
and ( n17053 , n16179 , n16182 );
or ( n17054 , n17052 , n17053 );
xor ( n17055 , n17051 , n17054 );
nor ( n17056 , n3300 , n1178 );
xor ( n17057 , n17055 , n17056 );
and ( n17058 , n16183 , n16184 );
and ( n17059 , n16185 , n16188 );
or ( n17060 , n17058 , n17059 );
xor ( n17061 , n17057 , n17060 );
nor ( n17062 , n3570 , n1305 );
xor ( n17063 , n17061 , n17062 );
and ( n17064 , n16189 , n16190 );
and ( n17065 , n16191 , n16194 );
or ( n17066 , n17064 , n17065 );
xor ( n17067 , n17063 , n17066 );
nor ( n17068 , n3853 , n1447 );
xor ( n17069 , n17067 , n17068 );
and ( n17070 , n16195 , n16196 );
and ( n17071 , n16197 , n16200 );
or ( n17072 , n17070 , n17071 );
xor ( n17073 , n17069 , n17072 );
nor ( n17074 , n4151 , n1600 );
xor ( n17075 , n17073 , n17074 );
and ( n17076 , n16201 , n16202 );
and ( n17077 , n16203 , n16206 );
or ( n17078 , n17076 , n17077 );
xor ( n17079 , n17075 , n17078 );
nor ( n17080 , n4458 , n1768 );
xor ( n17081 , n17079 , n17080 );
and ( n17082 , n16207 , n16208 );
and ( n17083 , n16209 , n16212 );
or ( n17084 , n17082 , n17083 );
xor ( n17085 , n17081 , n17084 );
nor ( n17086 , n4786 , n1947 );
xor ( n17087 , n17085 , n17086 );
and ( n17088 , n16213 , n16214 );
and ( n17089 , n16215 , n16218 );
or ( n17090 , n17088 , n17089 );
xor ( n17091 , n17087 , n17090 );
nor ( n17092 , n5126 , n2139 );
xor ( n17093 , n17091 , n17092 );
and ( n17094 , n16219 , n16220 );
and ( n17095 , n16221 , n16224 );
or ( n17096 , n17094 , n17095 );
xor ( n17097 , n17093 , n17096 );
nor ( n17098 , n5477 , n2345 );
xor ( n17099 , n17097 , n17098 );
and ( n17100 , n16225 , n16226 );
and ( n17101 , n16227 , n16230 );
or ( n17102 , n17100 , n17101 );
xor ( n17103 , n17099 , n17102 );
nor ( n17104 , n5838 , n2568 );
xor ( n17105 , n17103 , n17104 );
and ( n17106 , n16231 , n16232 );
and ( n17107 , n16233 , n16236 );
or ( n17108 , n17106 , n17107 );
xor ( n17109 , n17105 , n17108 );
nor ( n17110 , n6212 , n2799 );
xor ( n17111 , n17109 , n17110 );
and ( n17112 , n16237 , n16238 );
and ( n17113 , n16239 , n16242 );
or ( n17114 , n17112 , n17113 );
xor ( n17115 , n17111 , n17114 );
nor ( n17116 , n6596 , n3045 );
xor ( n17117 , n17115 , n17116 );
and ( n17118 , n16243 , n16244 );
and ( n17119 , n16245 , n16248 );
or ( n17120 , n17118 , n17119 );
xor ( n17121 , n17117 , n17120 );
nor ( n17122 , n6997 , n3302 );
xor ( n17123 , n17121 , n17122 );
and ( n17124 , n16249 , n16250 );
and ( n17125 , n16251 , n16254 );
or ( n17126 , n17124 , n17125 );
xor ( n17127 , n17123 , n17126 );
nor ( n17128 , n7413 , n3572 );
xor ( n17129 , n17127 , n17128 );
and ( n17130 , n16255 , n16256 );
and ( n17131 , n16257 , n16260 );
or ( n17132 , n17130 , n17131 );
xor ( n17133 , n17129 , n17132 );
nor ( n17134 , n7841 , n3855 );
xor ( n17135 , n17133 , n17134 );
and ( n17136 , n16261 , n16262 );
and ( n17137 , n16263 , n16266 );
or ( n17138 , n17136 , n17137 );
xor ( n17139 , n17135 , n17138 );
nor ( n17140 , n8281 , n4153 );
xor ( n17141 , n17139 , n17140 );
and ( n17142 , n16267 , n16268 );
and ( n17143 , n16269 , n16272 );
or ( n17144 , n17142 , n17143 );
xor ( n17145 , n17141 , n17144 );
nor ( n17146 , n8737 , n4460 );
xor ( n17147 , n17145 , n17146 );
and ( n17148 , n16273 , n16274 );
and ( n17149 , n16275 , n16278 );
or ( n17150 , n17148 , n17149 );
xor ( n17151 , n17147 , n17150 );
nor ( n17152 , n9420 , n4788 );
xor ( n17153 , n17151 , n17152 );
and ( n17154 , n16279 , n16280 );
and ( n17155 , n16281 , n16284 );
or ( n17156 , n17154 , n17155 );
xor ( n17157 , n17153 , n17156 );
nor ( n17158 , n10312 , n5128 );
xor ( n17159 , n17157 , n17158 );
and ( n17160 , n16285 , n16286 );
and ( n17161 , n16287 , n16290 );
or ( n17162 , n17160 , n17161 );
xor ( n17163 , n17159 , n17162 );
nor ( n17164 , n11041 , n5479 );
xor ( n17165 , n17163 , n17164 );
and ( n17166 , n16291 , n16292 );
and ( n17167 , n16293 , n16296 );
or ( n17168 , n17166 , n17167 );
xor ( n17169 , n17165 , n17168 );
nor ( n17170 , n11790 , n5840 );
xor ( n17171 , n17169 , n17170 );
and ( n17172 , n16297 , n16298 );
and ( n17173 , n16299 , n16302 );
or ( n17174 , n17172 , n17173 );
xor ( n17175 , n17171 , n17174 );
nor ( n17176 , n12555 , n6214 );
xor ( n17177 , n17175 , n17176 );
and ( n17178 , n16303 , n16304 );
and ( n17179 , n16305 , n16308 );
or ( n17180 , n17178 , n17179 );
xor ( n17181 , n17177 , n17180 );
nor ( n17182 , n13340 , n6598 );
xor ( n17183 , n17181 , n17182 );
and ( n17184 , n16309 , n16310 );
and ( n17185 , n16311 , n16314 );
or ( n17186 , n17184 , n17185 );
xor ( n17187 , n17183 , n17186 );
nor ( n17188 , n14138 , n6999 );
xor ( n17189 , n17187 , n17188 );
and ( n17190 , n16315 , n16316 );
and ( n17191 , n16317 , n16320 );
or ( n17192 , n17190 , n17191 );
xor ( n17193 , n17189 , n17192 );
nor ( n17194 , n14959 , n7415 );
xor ( n17195 , n17193 , n17194 );
and ( n17196 , n16321 , n16322 );
and ( n17197 , n16323 , n16326 );
or ( n17198 , n17196 , n17197 );
xor ( n17199 , n17195 , n17198 );
nor ( n17200 , n15800 , n7843 );
xor ( n17201 , n17199 , n17200 );
and ( n17202 , n16327 , n16328 );
and ( n17203 , n16329 , n16332 );
or ( n17204 , n17202 , n17203 );
xor ( n17205 , n17201 , n17204 );
nor ( n17206 , n16660 , n8283 );
xor ( n17207 , n17205 , n17206 );
and ( n17208 , n16333 , n16334 );
and ( n17209 , n16335 , n16338 );
or ( n17210 , n17208 , n17209 );
xor ( n17211 , n17207 , n17210 );
and ( n17212 , n16646 , n16650 );
and ( n17213 , n16349 , n16644 );
and ( n17214 , n16644 , n16651 );
and ( n17215 , n16349 , n16651 );
or ( n17216 , n17213 , n17214 , n17215 );
xor ( n17217 , n17212 , n17216 );
and ( n17218 , n16353 , n16560 );
and ( n17219 , n16560 , n16643 );
and ( n17220 , n16353 , n16643 );
or ( n17221 , n17218 , n17219 , n17220 );
and ( n17222 , n16357 , n16435 );
and ( n17223 , n16435 , n16559 );
and ( n17224 , n16357 , n16559 );
or ( n17225 , n17222 , n17223 , n17224 );
and ( n17226 , n16440 , n16487 );
and ( n17227 , n16487 , n16558 );
and ( n17228 , n16440 , n16558 );
or ( n17229 , n17226 , n17227 , n17228 );
and ( n17230 , n16370 , n16407 );
and ( n17231 , n16407 , n16433 );
and ( n17232 , n16370 , n16433 );
or ( n17233 , n17230 , n17231 , n17232 );
and ( n17234 , n16444 , n16448 );
and ( n17235 , n16448 , n16486 );
and ( n17236 , n16444 , n16486 );
or ( n17237 , n17234 , n17235 , n17236 );
xor ( n17238 , n17233 , n17237 );
and ( n17239 , n16412 , n16416 );
and ( n17240 , n16416 , n16432 );
and ( n17241 , n16412 , n16432 );
or ( n17242 , n17239 , n17240 , n17241 );
and ( n17243 , n16394 , n16399 );
and ( n17244 , n16399 , n16405 );
and ( n17245 , n16394 , n16405 );
or ( n17246 , n17243 , n17244 , n17245 );
and ( n17247 , n16384 , n16385 );
and ( n17248 , n16385 , n16387 );
and ( n17249 , n16384 , n16387 );
or ( n17250 , n17247 , n17248 , n17249 );
and ( n17251 , n16395 , n16396 );
and ( n17252 , n16396 , n16398 );
and ( n17253 , n16395 , n16398 );
or ( n17254 , n17251 , n17252 , n17253 );
xor ( n17255 , n17250 , n17254 );
and ( n17256 , n7385 , n1738 );
and ( n17257 , n7808 , n1551 );
xor ( n17258 , n17256 , n17257 );
and ( n17259 , n8079 , n1424 );
xor ( n17260 , n17258 , n17259 );
xor ( n17261 , n17255 , n17260 );
xor ( n17262 , n17246 , n17261 );
and ( n17263 , n16401 , n16402 );
and ( n17264 , n16402 , n16404 );
and ( n17265 , n16401 , n16404 );
or ( n17266 , n17263 , n17264 , n17265 );
and ( n17267 , n6187 , n2298 );
and ( n17268 , n6569 , n2100 );
xor ( n17269 , n17267 , n17268 );
and ( n17270 , n6816 , n1882 );
xor ( n17271 , n17269 , n17270 );
xor ( n17272 , n17266 , n17271 );
and ( n17273 , n4959 , n2981 );
and ( n17274 , n5459 , n2739 );
xor ( n17275 , n17273 , n17274 );
and ( n17276 , n5819 , n2544 );
xor ( n17277 , n17275 , n17276 );
xor ( n17278 , n17272 , n17277 );
xor ( n17279 , n17262 , n17278 );
xor ( n17280 , n17242 , n17279 );
and ( n17281 , n16421 , n16425 );
and ( n17282 , n16425 , n16431 );
and ( n17283 , n16421 , n16431 );
or ( n17284 , n17281 , n17282 , n17283 );
and ( n17285 , n16457 , n16462 );
and ( n17286 , n16462 , n16468 );
and ( n17287 , n16457 , n16468 );
or ( n17288 , n17285 , n17286 , n17287 );
xor ( n17289 , n17284 , n17288 );
and ( n17290 , n16427 , n16428 );
and ( n17291 , n16428 , n16430 );
and ( n17292 , n16427 , n16430 );
or ( n17293 , n17290 , n17291 , n17292 );
and ( n17294 , n16458 , n16459 );
and ( n17295 , n16459 , n16461 );
and ( n17296 , n16458 , n16461 );
or ( n17297 , n17294 , n17295 , n17296 );
xor ( n17298 , n17293 , n17297 );
and ( n17299 , n4132 , n3749 );
and ( n17300 , n4438 , n3495 );
xor ( n17301 , n17299 , n17300 );
and ( n17302 , n4766 , n3271 );
xor ( n17303 , n17301 , n17302 );
xor ( n17304 , n17298 , n17303 );
xor ( n17305 , n17289 , n17304 );
xor ( n17306 , n17280 , n17305 );
xor ( n17307 , n17238 , n17306 );
xor ( n17308 , n17229 , n17307 );
and ( n17309 , n16492 , n16518 );
and ( n17310 , n16518 , n16557 );
and ( n17311 , n16492 , n16557 );
or ( n17312 , n17309 , n17310 , n17311 );
and ( n17313 , n16453 , n16469 );
and ( n17314 , n16469 , n16485 );
and ( n17315 , n16453 , n16485 );
or ( n17316 , n17313 , n17314 , n17315 );
and ( n17317 , n16496 , n16500 );
and ( n17318 , n16500 , n16517 );
and ( n17319 , n16496 , n16517 );
or ( n17320 , n17317 , n17318 , n17319 );
xor ( n17321 , n17316 , n17320 );
and ( n17322 , n16474 , n16478 );
and ( n17323 , n16478 , n16484 );
and ( n17324 , n16474 , n16484 );
or ( n17325 , n17322 , n17323 , n17324 );
and ( n17326 , n16464 , n16465 );
and ( n17327 , n16465 , n16467 );
and ( n17328 , n16464 , n16467 );
or ( n17329 , n17326 , n17327 , n17328 );
and ( n17330 , n3182 , n4730 );
and ( n17331 , n3545 , n4403 );
xor ( n17332 , n17330 , n17331 );
and ( n17333 , n3801 , n4102 );
xor ( n17334 , n17332 , n17333 );
xor ( n17335 , n17329 , n17334 );
and ( n17336 , n2462 , n5765 );
and ( n17337 , n2779 , n5408 );
xor ( n17338 , n17336 , n17337 );
and ( n17339 , n3024 , n5103 );
xor ( n17340 , n17338 , n17339 );
xor ( n17341 , n17335 , n17340 );
xor ( n17342 , n17325 , n17341 );
and ( n17343 , n16480 , n16481 );
and ( n17344 , n16481 , n16483 );
and ( n17345 , n16480 , n16483 );
or ( n17346 , n17343 , n17344 , n17345 );
and ( n17347 , n16506 , n16507 );
and ( n17348 , n16507 , n16509 );
and ( n17349 , n16506 , n16509 );
or ( n17350 , n17347 , n17348 , n17349 );
xor ( n17351 , n17346 , n17350 );
and ( n17352 , n1933 , n6971 );
and ( n17353 , n2120 , n6504 );
xor ( n17354 , n17352 , n17353 );
and ( n17355 , n2324 , n6132 );
xor ( n17356 , n17354 , n17355 );
xor ( n17357 , n17351 , n17356 );
xor ( n17358 , n17342 , n17357 );
xor ( n17359 , n17321 , n17358 );
xor ( n17360 , n17312 , n17359 );
and ( n17361 , n16523 , n16538 );
and ( n17362 , n16538 , n16556 );
and ( n17363 , n16523 , n16556 );
or ( n17364 , n17361 , n17362 , n17363 );
and ( n17365 , n16505 , n16510 );
and ( n17366 , n16510 , n16516 );
and ( n17367 , n16505 , n16516 );
or ( n17368 , n17365 , n17366 , n17367 );
and ( n17369 , n16527 , n16531 );
and ( n17370 , n16531 , n16537 );
and ( n17371 , n16527 , n16537 );
or ( n17372 , n17369 , n17370 , n17371 );
xor ( n17373 , n17368 , n17372 );
and ( n17374 , n16512 , n16513 );
and ( n17375 , n16513 , n16515 );
and ( n17376 , n16512 , n16515 );
or ( n17377 , n17374 , n17375 , n17376 );
and ( n17378 , n1383 , n8243 );
and ( n17379 , n1580 , n7662 );
xor ( n17380 , n17378 , n17379 );
and ( n17381 , n1694 , n7310 );
xor ( n17382 , n17380 , n17381 );
xor ( n17383 , n17377 , n17382 );
and ( n17384 , n1047 , n10239 );
and ( n17385 , n1164 , n9348 );
xor ( n17386 , n17384 , n17385 );
and ( n17387 , n1287 , n8669 );
xor ( n17388 , n17386 , n17387 );
xor ( n17389 , n17383 , n17388 );
xor ( n17390 , n17373 , n17389 );
xor ( n17391 , n17364 , n17390 );
and ( n17392 , n16543 , n16548 );
and ( n17393 , n16548 , n16555 );
and ( n17394 , n16543 , n16555 );
or ( n17395 , n17392 , n17393 , n17394 );
and ( n17396 , n16533 , n16534 );
and ( n17397 , n16534 , n16536 );
and ( n17398 , n16533 , n16536 );
or ( n17399 , n17396 , n17397 , n17398 );
and ( n17400 , n16544 , n16545 );
and ( n17401 , n16545 , n16547 );
and ( n17402 , n16544 , n16547 );
or ( n17403 , n17400 , n17401 , n17402 );
xor ( n17404 , n17399 , n17403 );
and ( n17405 , n783 , n12531 );
and ( n17406 , n856 , n11718 );
xor ( n17407 , n17405 , n17406 );
and ( n17408 , n925 , n10977 );
xor ( n17409 , n17407 , n17408 );
xor ( n17410 , n17404 , n17409 );
xor ( n17411 , n17395 , n17410 );
and ( n17412 , n16551 , n16552 );
and ( n17413 , n16552 , n16554 );
and ( n17414 , n16551 , n16554 );
or ( n17415 , n17412 , n17413 , n17414 );
and ( n17416 , n632 , n14838 );
and ( n17417 , n671 , n14044 );
xor ( n17418 , n17416 , n17417 );
and ( n17419 , n715 , n13256 );
xor ( n17420 , n17418 , n17419 );
xor ( n17421 , n17415 , n17420 );
buf ( n17422 , n423 );
and ( n17423 , n599 , n17422 );
and ( n17424 , n608 , n16550 );
xor ( n17425 , n17423 , n17424 );
and ( n17426 , n611 , n15691 );
xor ( n17427 , n17425 , n17426 );
xor ( n17428 , n17421 , n17427 );
xor ( n17429 , n17411 , n17428 );
xor ( n17430 , n17391 , n17429 );
xor ( n17431 , n17360 , n17430 );
xor ( n17432 , n17308 , n17431 );
xor ( n17433 , n17225 , n17432 );
and ( n17434 , n16361 , n16365 );
and ( n17435 , n16365 , n16434 );
and ( n17436 , n16361 , n16434 );
or ( n17437 , n17434 , n17435 , n17436 );
and ( n17438 , n16574 , n16610 );
and ( n17439 , n16610 , n16641 );
and ( n17440 , n16574 , n16641 );
or ( n17441 , n17438 , n17439 , n17440 );
xor ( n17442 , n17437 , n17441 );
and ( n17443 , n16578 , n16582 );
and ( n17444 , n16582 , n16609 );
and ( n17445 , n16578 , n16609 );
or ( n17446 , n17443 , n17444 , n17445 );
and ( n17447 , n16587 , n16591 );
and ( n17448 , n16591 , n16608 );
and ( n17449 , n16587 , n16608 );
or ( n17450 , n17447 , n17448 , n17449 );
and ( n17451 , n16374 , n16389 );
and ( n17452 , n16389 , n16406 );
and ( n17453 , n16374 , n16406 );
or ( n17454 , n17451 , n17452 , n17453 );
xor ( n17455 , n17450 , n17454 );
and ( n17456 , n16596 , n16601 );
and ( n17457 , n16601 , n16607 );
and ( n17458 , n16596 , n16607 );
or ( n17459 , n17456 , n17457 , n17458 );
and ( n17460 , n16378 , n16382 );
and ( n17461 , n16382 , n16388 );
and ( n17462 , n16378 , n16388 );
or ( n17463 , n17460 , n17461 , n17462 );
xor ( n17464 , n17459 , n17463 );
and ( n17465 , n16603 , n16604 );
and ( n17466 , n16604 , n16606 );
and ( n17467 , n16603 , n16606 );
or ( n17468 , n17465 , n17466 , n17467 );
and ( n17469 , n11015 , n940 );
and ( n17470 , n11769 , n840 );
xor ( n17471 , n17469 , n17470 );
and ( n17472 , n12320 , n771 );
xor ( n17473 , n17471 , n17472 );
xor ( n17474 , n17468 , n17473 );
and ( n17475 , n8718 , n1254 );
and ( n17476 , n9400 , n1134 );
xor ( n17477 , n17475 , n17476 );
and ( n17478 , n10291 , n1034 );
xor ( n17479 , n17477 , n17478 );
xor ( n17480 , n17474 , n17479 );
xor ( n17481 , n17464 , n17480 );
xor ( n17482 , n17455 , n17481 );
xor ( n17483 , n17446 , n17482 );
and ( n17484 , n16619 , n16634 );
and ( n17485 , n16634 , n16639 );
and ( n17486 , n16619 , n16639 );
or ( n17487 , n17484 , n17485 , n17486 );
and ( n17488 , n16623 , n16627 );
and ( n17489 , n16627 , n16633 );
and ( n17490 , n16623 , n16633 );
or ( n17491 , n17488 , n17489 , n17490 );
and ( n17492 , n16629 , n16630 );
and ( n17493 , n16630 , n16632 );
and ( n17494 , n16629 , n16632 );
or ( n17495 , n17492 , n17493 , n17494 );
and ( n17496 , n16597 , n16598 );
and ( n17497 , n16598 , n16600 );
and ( n17498 , n16597 , n16600 );
or ( n17499 , n17496 , n17497 , n17498 );
xor ( n17500 , n17495 , n17499 );
and ( n17501 , n13322 , n719 );
and ( n17502 , n14118 , n663 );
xor ( n17503 , n17501 , n17502 );
and ( n17504 , n14938 , n635 );
xor ( n17505 , n17503 , n17504 );
xor ( n17506 , n17500 , n17505 );
xor ( n17507 , n17491 , n17506 );
and ( n17508 , n16636 , n16638 );
and ( n17509 , n15758 , n606 );
and ( n17510 , n16637 , n615 );
xor ( n17511 , n17509 , n17510 );
buf ( n17512 , n423 );
and ( n17513 , n17512 , n612 );
xor ( n17514 , n17511 , n17513 );
xor ( n17515 , n17508 , n17514 );
xor ( n17516 , n17507 , n17515 );
xor ( n17517 , n17487 , n17516 );
xor ( n17518 , n17483 , n17517 );
xor ( n17519 , n17442 , n17518 );
xor ( n17520 , n17433 , n17519 );
xor ( n17521 , n17221 , n17520 );
and ( n17522 , n16615 , n16640 );
and ( n17523 , n16565 , n16569 );
and ( n17524 , n16569 , n16642 );
and ( n17525 , n16565 , n16642 );
or ( n17526 , n17523 , n17524 , n17525 );
xor ( n17527 , n17522 , n17526 );
xor ( n17528 , n17521 , n17527 );
xor ( n17529 , n17217 , n17528 );
and ( n17530 , n16340 , n16344 );
and ( n17531 , n16344 , n16652 );
and ( n17532 , n16340 , n16652 );
or ( n17533 , n17530 , n17531 , n17532 );
xor ( n17534 , n17529 , n17533 );
and ( n17535 , n16653 , n16656 );
xor ( n17536 , n17534 , n17535 );
buf ( n17537 , n17536 );
buf ( n17538 , n17537 );
not ( n17539 , n17538 );
nor ( n17540 , n17539 , n8739 );
xor ( n17541 , n17211 , n17540 );
and ( n17542 , n16339 , n16661 );
and ( n17543 , n16662 , n16665 );
or ( n17544 , n17542 , n17543 );
xor ( n17545 , n17541 , n17544 );
buf ( n17546 , n17545 );
buf ( n17547 , n17546 );
not ( n17548 , n17547 );
buf ( n17549 , n546 );
not ( n17550 , n17549 );
nor ( n17551 , n17548 , n17550 );
xor ( n17552 , n16941 , n17551 );
xor ( n17553 , n16677 , n16938 );
nor ( n17554 , n16669 , n17550 );
and ( n17555 , n17553 , n17554 );
xor ( n17556 , n17553 , n17554 );
xor ( n17557 , n16681 , n16936 );
nor ( n17558 , n15809 , n17550 );
and ( n17559 , n17557 , n17558 );
xor ( n17560 , n17557 , n17558 );
xor ( n17561 , n16685 , n16934 );
nor ( n17562 , n14968 , n17550 );
and ( n17563 , n17561 , n17562 );
xor ( n17564 , n17561 , n17562 );
xor ( n17565 , n16689 , n16932 );
nor ( n17566 , n14147 , n17550 );
and ( n17567 , n17565 , n17566 );
xor ( n17568 , n17565 , n17566 );
xor ( n17569 , n16693 , n16930 );
nor ( n17570 , n13349 , n17550 );
and ( n17571 , n17569 , n17570 );
xor ( n17572 , n17569 , n17570 );
xor ( n17573 , n16697 , n16928 );
nor ( n17574 , n12564 , n17550 );
and ( n17575 , n17573 , n17574 );
xor ( n17576 , n17573 , n17574 );
xor ( n17577 , n16701 , n16926 );
nor ( n17578 , n11799 , n17550 );
and ( n17579 , n17577 , n17578 );
xor ( n17580 , n17577 , n17578 );
xor ( n17581 , n16705 , n16924 );
nor ( n17582 , n11050 , n17550 );
and ( n17583 , n17581 , n17582 );
xor ( n17584 , n17581 , n17582 );
xor ( n17585 , n16709 , n16922 );
nor ( n17586 , n10321 , n17550 );
and ( n17587 , n17585 , n17586 );
xor ( n17588 , n17585 , n17586 );
xor ( n17589 , n16713 , n16920 );
nor ( n17590 , n9429 , n17550 );
and ( n17591 , n17589 , n17590 );
xor ( n17592 , n17589 , n17590 );
xor ( n17593 , n16717 , n16918 );
nor ( n17594 , n8949 , n17550 );
and ( n17595 , n17593 , n17594 );
xor ( n17596 , n17593 , n17594 );
xor ( n17597 , n16721 , n16916 );
nor ( n17598 , n9437 , n17550 );
and ( n17599 , n17597 , n17598 );
xor ( n17600 , n17597 , n17598 );
xor ( n17601 , n16725 , n16914 );
nor ( n17602 , n9446 , n17550 );
and ( n17603 , n17601 , n17602 );
xor ( n17604 , n17601 , n17602 );
xor ( n17605 , n16729 , n16912 );
nor ( n17606 , n9455 , n17550 );
and ( n17607 , n17605 , n17606 );
xor ( n17608 , n17605 , n17606 );
xor ( n17609 , n16733 , n16910 );
nor ( n17610 , n9464 , n17550 );
and ( n17611 , n17609 , n17610 );
xor ( n17612 , n17609 , n17610 );
xor ( n17613 , n16737 , n16908 );
nor ( n17614 , n9473 , n17550 );
and ( n17615 , n17613 , n17614 );
xor ( n17616 , n17613 , n17614 );
xor ( n17617 , n16741 , n16906 );
nor ( n17618 , n9482 , n17550 );
and ( n17619 , n17617 , n17618 );
xor ( n17620 , n17617 , n17618 );
xor ( n17621 , n16745 , n16904 );
nor ( n17622 , n9491 , n17550 );
and ( n17623 , n17621 , n17622 );
xor ( n17624 , n17621 , n17622 );
xor ( n17625 , n16749 , n16902 );
nor ( n17626 , n9500 , n17550 );
and ( n17627 , n17625 , n17626 );
xor ( n17628 , n17625 , n17626 );
xor ( n17629 , n16753 , n16900 );
nor ( n17630 , n9509 , n17550 );
and ( n17631 , n17629 , n17630 );
xor ( n17632 , n17629 , n17630 );
xor ( n17633 , n16757 , n16898 );
nor ( n17634 , n9518 , n17550 );
and ( n17635 , n17633 , n17634 );
xor ( n17636 , n17633 , n17634 );
xor ( n17637 , n16761 , n16896 );
nor ( n17638 , n9527 , n17550 );
and ( n17639 , n17637 , n17638 );
xor ( n17640 , n17637 , n17638 );
xor ( n17641 , n16765 , n16894 );
nor ( n17642 , n9536 , n17550 );
and ( n17643 , n17641 , n17642 );
xor ( n17644 , n17641 , n17642 );
xor ( n17645 , n16769 , n16892 );
nor ( n17646 , n9545 , n17550 );
and ( n17647 , n17645 , n17646 );
xor ( n17648 , n17645 , n17646 );
xor ( n17649 , n16773 , n16890 );
nor ( n17650 , n9554 , n17550 );
and ( n17651 , n17649 , n17650 );
xor ( n17652 , n17649 , n17650 );
xor ( n17653 , n16777 , n16888 );
nor ( n17654 , n9563 , n17550 );
and ( n17655 , n17653 , n17654 );
xor ( n17656 , n17653 , n17654 );
xor ( n17657 , n16781 , n16886 );
nor ( n17658 , n9572 , n17550 );
and ( n17659 , n17657 , n17658 );
xor ( n17660 , n17657 , n17658 );
xor ( n17661 , n16785 , n16884 );
nor ( n17662 , n9581 , n17550 );
and ( n17663 , n17661 , n17662 );
xor ( n17664 , n17661 , n17662 );
xor ( n17665 , n16789 , n16882 );
nor ( n17666 , n9590 , n17550 );
and ( n17667 , n17665 , n17666 );
xor ( n17668 , n17665 , n17666 );
xor ( n17669 , n16793 , n16880 );
nor ( n17670 , n9599 , n17550 );
and ( n17671 , n17669 , n17670 );
xor ( n17672 , n17669 , n17670 );
xor ( n17673 , n16797 , n16878 );
nor ( n17674 , n9608 , n17550 );
and ( n17675 , n17673 , n17674 );
xor ( n17676 , n17673 , n17674 );
xor ( n17677 , n16801 , n16876 );
nor ( n17678 , n9617 , n17550 );
and ( n17679 , n17677 , n17678 );
xor ( n17680 , n17677 , n17678 );
xor ( n17681 , n16805 , n16874 );
nor ( n17682 , n9626 , n17550 );
and ( n17683 , n17681 , n17682 );
xor ( n17684 , n17681 , n17682 );
xor ( n17685 , n16809 , n16872 );
nor ( n17686 , n9635 , n17550 );
and ( n17687 , n17685 , n17686 );
xor ( n17688 , n17685 , n17686 );
xor ( n17689 , n16813 , n16870 );
nor ( n17690 , n9644 , n17550 );
and ( n17691 , n17689 , n17690 );
xor ( n17692 , n17689 , n17690 );
xor ( n17693 , n16817 , n16868 );
nor ( n17694 , n9653 , n17550 );
and ( n17695 , n17693 , n17694 );
xor ( n17696 , n17693 , n17694 );
xor ( n17697 , n16821 , n16866 );
nor ( n17698 , n9662 , n17550 );
and ( n17699 , n17697 , n17698 );
xor ( n17700 , n17697 , n17698 );
xor ( n17701 , n16825 , n16864 );
nor ( n17702 , n9671 , n17550 );
and ( n17703 , n17701 , n17702 );
xor ( n17704 , n17701 , n17702 );
xor ( n17705 , n16829 , n16862 );
nor ( n17706 , n9680 , n17550 );
and ( n17707 , n17705 , n17706 );
xor ( n17708 , n17705 , n17706 );
xor ( n17709 , n16833 , n16860 );
nor ( n17710 , n9689 , n17550 );
and ( n17711 , n17709 , n17710 );
xor ( n17712 , n17709 , n17710 );
xor ( n17713 , n16837 , n16858 );
nor ( n17714 , n9698 , n17550 );
and ( n17715 , n17713 , n17714 );
xor ( n17716 , n17713 , n17714 );
xor ( n17717 , n16841 , n16856 );
nor ( n17718 , n9707 , n17550 );
and ( n17719 , n17717 , n17718 );
xor ( n17720 , n17717 , n17718 );
xor ( n17721 , n16845 , n16854 );
nor ( n17722 , n9716 , n17550 );
and ( n17723 , n17721 , n17722 );
xor ( n17724 , n17721 , n17722 );
xor ( n17725 , n16849 , n16852 );
nor ( n17726 , n9725 , n17550 );
and ( n17727 , n17725 , n17726 );
xor ( n17728 , n17725 , n17726 );
xor ( n17729 , n16850 , n16851 );
nor ( n17730 , n9734 , n17550 );
and ( n17731 , n17729 , n17730 );
xor ( n17732 , n17729 , n17730 );
nor ( n17733 , n9752 , n16671 );
nor ( n17734 , n9743 , n17550 );
and ( n17735 , n17733 , n17734 );
and ( n17736 , n17732 , n17735 );
or ( n17737 , n17731 , n17736 );
and ( n17738 , n17728 , n17737 );
or ( n17739 , n17727 , n17738 );
and ( n17740 , n17724 , n17739 );
or ( n17741 , n17723 , n17740 );
and ( n17742 , n17720 , n17741 );
or ( n17743 , n17719 , n17742 );
and ( n17744 , n17716 , n17743 );
or ( n17745 , n17715 , n17744 );
and ( n17746 , n17712 , n17745 );
or ( n17747 , n17711 , n17746 );
and ( n17748 , n17708 , n17747 );
or ( n17749 , n17707 , n17748 );
and ( n17750 , n17704 , n17749 );
or ( n17751 , n17703 , n17750 );
and ( n17752 , n17700 , n17751 );
or ( n17753 , n17699 , n17752 );
and ( n17754 , n17696 , n17753 );
or ( n17755 , n17695 , n17754 );
and ( n17756 , n17692 , n17755 );
or ( n17757 , n17691 , n17756 );
and ( n17758 , n17688 , n17757 );
or ( n17759 , n17687 , n17758 );
and ( n17760 , n17684 , n17759 );
or ( n17761 , n17683 , n17760 );
and ( n17762 , n17680 , n17761 );
or ( n17763 , n17679 , n17762 );
and ( n17764 , n17676 , n17763 );
or ( n17765 , n17675 , n17764 );
and ( n17766 , n17672 , n17765 );
or ( n17767 , n17671 , n17766 );
and ( n17768 , n17668 , n17767 );
or ( n17769 , n17667 , n17768 );
and ( n17770 , n17664 , n17769 );
or ( n17771 , n17663 , n17770 );
and ( n17772 , n17660 , n17771 );
or ( n17773 , n17659 , n17772 );
and ( n17774 , n17656 , n17773 );
or ( n17775 , n17655 , n17774 );
and ( n17776 , n17652 , n17775 );
or ( n17777 , n17651 , n17776 );
and ( n17778 , n17648 , n17777 );
or ( n17779 , n17647 , n17778 );
and ( n17780 , n17644 , n17779 );
or ( n17781 , n17643 , n17780 );
and ( n17782 , n17640 , n17781 );
or ( n17783 , n17639 , n17782 );
and ( n17784 , n17636 , n17783 );
or ( n17785 , n17635 , n17784 );
and ( n17786 , n17632 , n17785 );
or ( n17787 , n17631 , n17786 );
and ( n17788 , n17628 , n17787 );
or ( n17789 , n17627 , n17788 );
and ( n17790 , n17624 , n17789 );
or ( n17791 , n17623 , n17790 );
and ( n17792 , n17620 , n17791 );
or ( n17793 , n17619 , n17792 );
and ( n17794 , n17616 , n17793 );
or ( n17795 , n17615 , n17794 );
and ( n17796 , n17612 , n17795 );
or ( n17797 , n17611 , n17796 );
and ( n17798 , n17608 , n17797 );
or ( n17799 , n17607 , n17798 );
and ( n17800 , n17604 , n17799 );
or ( n17801 , n17603 , n17800 );
and ( n17802 , n17600 , n17801 );
or ( n17803 , n17599 , n17802 );
and ( n17804 , n17596 , n17803 );
or ( n17805 , n17595 , n17804 );
and ( n17806 , n17592 , n17805 );
or ( n17807 , n17591 , n17806 );
and ( n17808 , n17588 , n17807 );
or ( n17809 , n17587 , n17808 );
and ( n17810 , n17584 , n17809 );
or ( n17811 , n17583 , n17810 );
and ( n17812 , n17580 , n17811 );
or ( n17813 , n17579 , n17812 );
and ( n17814 , n17576 , n17813 );
or ( n17815 , n17575 , n17814 );
and ( n17816 , n17572 , n17815 );
or ( n17817 , n17571 , n17816 );
and ( n17818 , n17568 , n17817 );
or ( n17819 , n17567 , n17818 );
and ( n17820 , n17564 , n17819 );
or ( n17821 , n17563 , n17820 );
and ( n17822 , n17560 , n17821 );
or ( n17823 , n17559 , n17822 );
and ( n17824 , n17556 , n17823 );
or ( n17825 , n17555 , n17824 );
xor ( n17826 , n17552 , n17825 );
buf ( n17827 , n486 );
not ( n17828 , n17827 );
nor ( n17829 , n601 , n17828 );
buf ( n17830 , n17829 );
nor ( n17831 , n622 , n16077 );
xor ( n17832 , n17830 , n17831 );
buf ( n17833 , n17832 );
nor ( n17834 , n646 , n15230 );
xor ( n17835 , n17833 , n17834 );
and ( n17836 , n16945 , n16946 );
buf ( n17837 , n17836 );
xor ( n17838 , n17835 , n17837 );
nor ( n17839 , n684 , n14403 );
xor ( n17840 , n17838 , n17839 );
and ( n17841 , n16948 , n16949 );
and ( n17842 , n16950 , n16952 );
or ( n17843 , n17841 , n17842 );
xor ( n17844 , n17840 , n17843 );
nor ( n17845 , n733 , n13599 );
xor ( n17846 , n17844 , n17845 );
and ( n17847 , n16953 , n16954 );
and ( n17848 , n16955 , n16958 );
or ( n17849 , n17847 , n17848 );
xor ( n17850 , n17846 , n17849 );
nor ( n17851 , n796 , n12808 );
xor ( n17852 , n17850 , n17851 );
and ( n17853 , n16959 , n16960 );
and ( n17854 , n16961 , n16964 );
or ( n17855 , n17853 , n17854 );
xor ( n17856 , n17852 , n17855 );
nor ( n17857 , n868 , n12037 );
xor ( n17858 , n17856 , n17857 );
and ( n17859 , n16965 , n16966 );
and ( n17860 , n16967 , n16970 );
or ( n17861 , n17859 , n17860 );
xor ( n17862 , n17858 , n17861 );
nor ( n17863 , n958 , n11282 );
xor ( n17864 , n17862 , n17863 );
and ( n17865 , n16971 , n16972 );
and ( n17866 , n16973 , n16976 );
or ( n17867 , n17865 , n17866 );
xor ( n17868 , n17864 , n17867 );
nor ( n17869 , n1062 , n10547 );
xor ( n17870 , n17868 , n17869 );
and ( n17871 , n16977 , n16978 );
and ( n17872 , n16979 , n16982 );
or ( n17873 , n17871 , n17872 );
xor ( n17874 , n17870 , n17873 );
nor ( n17875 , n1176 , n9829 );
xor ( n17876 , n17874 , n17875 );
and ( n17877 , n16983 , n16984 );
and ( n17878 , n16985 , n16988 );
or ( n17879 , n17877 , n17878 );
xor ( n17880 , n17876 , n17879 );
nor ( n17881 , n1303 , n8955 );
xor ( n17882 , n17880 , n17881 );
and ( n17883 , n16989 , n16990 );
and ( n17884 , n16991 , n16994 );
or ( n17885 , n17883 , n17884 );
xor ( n17886 , n17882 , n17885 );
nor ( n17887 , n1445 , n603 );
xor ( n17888 , n17886 , n17887 );
and ( n17889 , n16995 , n16996 );
and ( n17890 , n16997 , n17000 );
or ( n17891 , n17889 , n17890 );
xor ( n17892 , n17888 , n17891 );
nor ( n17893 , n1598 , n652 );
xor ( n17894 , n17892 , n17893 );
and ( n17895 , n17001 , n17002 );
and ( n17896 , n17003 , n17006 );
or ( n17897 , n17895 , n17896 );
xor ( n17898 , n17894 , n17897 );
nor ( n17899 , n1766 , n624 );
xor ( n17900 , n17898 , n17899 );
and ( n17901 , n17007 , n17008 );
and ( n17902 , n17009 , n17012 );
or ( n17903 , n17901 , n17902 );
xor ( n17904 , n17900 , n17903 );
nor ( n17905 , n1945 , n648 );
xor ( n17906 , n17904 , n17905 );
and ( n17907 , n17013 , n17014 );
and ( n17908 , n17015 , n17018 );
or ( n17909 , n17907 , n17908 );
xor ( n17910 , n17906 , n17909 );
nor ( n17911 , n2137 , n686 );
xor ( n17912 , n17910 , n17911 );
and ( n17913 , n17019 , n17020 );
and ( n17914 , n17021 , n17024 );
or ( n17915 , n17913 , n17914 );
xor ( n17916 , n17912 , n17915 );
nor ( n17917 , n2343 , n735 );
xor ( n17918 , n17916 , n17917 );
and ( n17919 , n17025 , n17026 );
and ( n17920 , n17027 , n17030 );
or ( n17921 , n17919 , n17920 );
xor ( n17922 , n17918 , n17921 );
nor ( n17923 , n2566 , n798 );
xor ( n17924 , n17922 , n17923 );
and ( n17925 , n17031 , n17032 );
and ( n17926 , n17033 , n17036 );
or ( n17927 , n17925 , n17926 );
xor ( n17928 , n17924 , n17927 );
nor ( n17929 , n2797 , n870 );
xor ( n17930 , n17928 , n17929 );
and ( n17931 , n17037 , n17038 );
and ( n17932 , n17039 , n17042 );
or ( n17933 , n17931 , n17932 );
xor ( n17934 , n17930 , n17933 );
nor ( n17935 , n3043 , n960 );
xor ( n17936 , n17934 , n17935 );
and ( n17937 , n17043 , n17044 );
and ( n17938 , n17045 , n17048 );
or ( n17939 , n17937 , n17938 );
xor ( n17940 , n17936 , n17939 );
nor ( n17941 , n3300 , n1064 );
xor ( n17942 , n17940 , n17941 );
and ( n17943 , n17049 , n17050 );
and ( n17944 , n17051 , n17054 );
or ( n17945 , n17943 , n17944 );
xor ( n17946 , n17942 , n17945 );
nor ( n17947 , n3570 , n1178 );
xor ( n17948 , n17946 , n17947 );
and ( n17949 , n17055 , n17056 );
and ( n17950 , n17057 , n17060 );
or ( n17951 , n17949 , n17950 );
xor ( n17952 , n17948 , n17951 );
nor ( n17953 , n3853 , n1305 );
xor ( n17954 , n17952 , n17953 );
and ( n17955 , n17061 , n17062 );
and ( n17956 , n17063 , n17066 );
or ( n17957 , n17955 , n17956 );
xor ( n17958 , n17954 , n17957 );
nor ( n17959 , n4151 , n1447 );
xor ( n17960 , n17958 , n17959 );
and ( n17961 , n17067 , n17068 );
and ( n17962 , n17069 , n17072 );
or ( n17963 , n17961 , n17962 );
xor ( n17964 , n17960 , n17963 );
nor ( n17965 , n4458 , n1600 );
xor ( n17966 , n17964 , n17965 );
and ( n17967 , n17073 , n17074 );
and ( n17968 , n17075 , n17078 );
or ( n17969 , n17967 , n17968 );
xor ( n17970 , n17966 , n17969 );
nor ( n17971 , n4786 , n1768 );
xor ( n17972 , n17970 , n17971 );
and ( n17973 , n17079 , n17080 );
and ( n17974 , n17081 , n17084 );
or ( n17975 , n17973 , n17974 );
xor ( n17976 , n17972 , n17975 );
nor ( n17977 , n5126 , n1947 );
xor ( n17978 , n17976 , n17977 );
and ( n17979 , n17085 , n17086 );
and ( n17980 , n17087 , n17090 );
or ( n17981 , n17979 , n17980 );
xor ( n17982 , n17978 , n17981 );
nor ( n17983 , n5477 , n2139 );
xor ( n17984 , n17982 , n17983 );
and ( n17985 , n17091 , n17092 );
and ( n17986 , n17093 , n17096 );
or ( n17987 , n17985 , n17986 );
xor ( n17988 , n17984 , n17987 );
nor ( n17989 , n5838 , n2345 );
xor ( n17990 , n17988 , n17989 );
and ( n17991 , n17097 , n17098 );
and ( n17992 , n17099 , n17102 );
or ( n17993 , n17991 , n17992 );
xor ( n17994 , n17990 , n17993 );
nor ( n17995 , n6212 , n2568 );
xor ( n17996 , n17994 , n17995 );
and ( n17997 , n17103 , n17104 );
and ( n17998 , n17105 , n17108 );
or ( n17999 , n17997 , n17998 );
xor ( n18000 , n17996 , n17999 );
nor ( n18001 , n6596 , n2799 );
xor ( n18002 , n18000 , n18001 );
and ( n18003 , n17109 , n17110 );
and ( n18004 , n17111 , n17114 );
or ( n18005 , n18003 , n18004 );
xor ( n18006 , n18002 , n18005 );
nor ( n18007 , n6997 , n3045 );
xor ( n18008 , n18006 , n18007 );
and ( n18009 , n17115 , n17116 );
and ( n18010 , n17117 , n17120 );
or ( n18011 , n18009 , n18010 );
xor ( n18012 , n18008 , n18011 );
nor ( n18013 , n7413 , n3302 );
xor ( n18014 , n18012 , n18013 );
and ( n18015 , n17121 , n17122 );
and ( n18016 , n17123 , n17126 );
or ( n18017 , n18015 , n18016 );
xor ( n18018 , n18014 , n18017 );
nor ( n18019 , n7841 , n3572 );
xor ( n18020 , n18018 , n18019 );
and ( n18021 , n17127 , n17128 );
and ( n18022 , n17129 , n17132 );
or ( n18023 , n18021 , n18022 );
xor ( n18024 , n18020 , n18023 );
nor ( n18025 , n8281 , n3855 );
xor ( n18026 , n18024 , n18025 );
and ( n18027 , n17133 , n17134 );
and ( n18028 , n17135 , n17138 );
or ( n18029 , n18027 , n18028 );
xor ( n18030 , n18026 , n18029 );
nor ( n18031 , n8737 , n4153 );
xor ( n18032 , n18030 , n18031 );
and ( n18033 , n17139 , n17140 );
and ( n18034 , n17141 , n17144 );
or ( n18035 , n18033 , n18034 );
xor ( n18036 , n18032 , n18035 );
nor ( n18037 , n9420 , n4460 );
xor ( n18038 , n18036 , n18037 );
and ( n18039 , n17145 , n17146 );
and ( n18040 , n17147 , n17150 );
or ( n18041 , n18039 , n18040 );
xor ( n18042 , n18038 , n18041 );
nor ( n18043 , n10312 , n4788 );
xor ( n18044 , n18042 , n18043 );
and ( n18045 , n17151 , n17152 );
and ( n18046 , n17153 , n17156 );
or ( n18047 , n18045 , n18046 );
xor ( n18048 , n18044 , n18047 );
nor ( n18049 , n11041 , n5128 );
xor ( n18050 , n18048 , n18049 );
and ( n18051 , n17157 , n17158 );
and ( n18052 , n17159 , n17162 );
or ( n18053 , n18051 , n18052 );
xor ( n18054 , n18050 , n18053 );
nor ( n18055 , n11790 , n5479 );
xor ( n18056 , n18054 , n18055 );
and ( n18057 , n17163 , n17164 );
and ( n18058 , n17165 , n17168 );
or ( n18059 , n18057 , n18058 );
xor ( n18060 , n18056 , n18059 );
nor ( n18061 , n12555 , n5840 );
xor ( n18062 , n18060 , n18061 );
and ( n18063 , n17169 , n17170 );
and ( n18064 , n17171 , n17174 );
or ( n18065 , n18063 , n18064 );
xor ( n18066 , n18062 , n18065 );
nor ( n18067 , n13340 , n6214 );
xor ( n18068 , n18066 , n18067 );
and ( n18069 , n17175 , n17176 );
and ( n18070 , n17177 , n17180 );
or ( n18071 , n18069 , n18070 );
xor ( n18072 , n18068 , n18071 );
nor ( n18073 , n14138 , n6598 );
xor ( n18074 , n18072 , n18073 );
and ( n18075 , n17181 , n17182 );
and ( n18076 , n17183 , n17186 );
or ( n18077 , n18075 , n18076 );
xor ( n18078 , n18074 , n18077 );
nor ( n18079 , n14959 , n6999 );
xor ( n18080 , n18078 , n18079 );
and ( n18081 , n17187 , n17188 );
and ( n18082 , n17189 , n17192 );
or ( n18083 , n18081 , n18082 );
xor ( n18084 , n18080 , n18083 );
nor ( n18085 , n15800 , n7415 );
xor ( n18086 , n18084 , n18085 );
and ( n18087 , n17193 , n17194 );
and ( n18088 , n17195 , n17198 );
or ( n18089 , n18087 , n18088 );
xor ( n18090 , n18086 , n18089 );
nor ( n18091 , n16660 , n7843 );
xor ( n18092 , n18090 , n18091 );
and ( n18093 , n17199 , n17200 );
and ( n18094 , n17201 , n17204 );
or ( n18095 , n18093 , n18094 );
xor ( n18096 , n18092 , n18095 );
nor ( n18097 , n17539 , n8283 );
xor ( n18098 , n18096 , n18097 );
and ( n18099 , n17205 , n17206 );
and ( n18100 , n17207 , n17210 );
or ( n18101 , n18099 , n18100 );
xor ( n18102 , n18098 , n18101 );
and ( n18103 , n17522 , n17526 );
and ( n18104 , n17221 , n17520 );
and ( n18105 , n17520 , n17527 );
and ( n18106 , n17221 , n17527 );
or ( n18107 , n18104 , n18105 , n18106 );
xor ( n18108 , n18103 , n18107 );
and ( n18109 , n17225 , n17432 );
and ( n18110 , n17432 , n17519 );
and ( n18111 , n17225 , n17519 );
or ( n18112 , n18109 , n18110 , n18111 );
and ( n18113 , n17229 , n17307 );
and ( n18114 , n17307 , n17431 );
and ( n18115 , n17229 , n17431 );
or ( n18116 , n18113 , n18114 , n18115 );
and ( n18117 , n17233 , n17237 );
and ( n18118 , n17237 , n17306 );
and ( n18119 , n17233 , n17306 );
or ( n18120 , n18117 , n18118 , n18119 );
and ( n18121 , n17446 , n17482 );
and ( n18122 , n17482 , n17517 );
and ( n18123 , n17446 , n17517 );
or ( n18124 , n18121 , n18122 , n18123 );
xor ( n18125 , n18120 , n18124 );
and ( n18126 , n17450 , n17454 );
and ( n18127 , n17454 , n17481 );
and ( n18128 , n17450 , n17481 );
or ( n18129 , n18126 , n18127 , n18128 );
and ( n18130 , n17508 , n17514 );
and ( n18131 , n17491 , n17506 );
and ( n18132 , n17506 , n17515 );
and ( n18133 , n17491 , n17515 );
or ( n18134 , n18131 , n18132 , n18133 );
xor ( n18135 , n18130 , n18134 );
and ( n18136 , n17495 , n17499 );
and ( n18137 , n17499 , n17505 );
and ( n18138 , n17495 , n17505 );
or ( n18139 , n18136 , n18137 , n18138 );
and ( n18140 , n17509 , n17510 );
and ( n18141 , n17510 , n17513 );
and ( n18142 , n17509 , n17513 );
or ( n18143 , n18140 , n18141 , n18142 );
buf ( n18144 , n422 );
and ( n18145 , n18144 , n612 );
xor ( n18146 , n18143 , n18145 );
and ( n18147 , n15758 , n635 );
and ( n18148 , n16637 , n606 );
xor ( n18149 , n18147 , n18148 );
and ( n18150 , n17512 , n615 );
xor ( n18151 , n18149 , n18150 );
xor ( n18152 , n18146 , n18151 );
xor ( n18153 , n18139 , n18152 );
and ( n18154 , n17501 , n17502 );
and ( n18155 , n17502 , n17504 );
and ( n18156 , n17501 , n17504 );
or ( n18157 , n18154 , n18155 , n18156 );
and ( n18158 , n17469 , n17470 );
and ( n18159 , n17470 , n17472 );
and ( n18160 , n17469 , n17472 );
or ( n18161 , n18158 , n18159 , n18160 );
xor ( n18162 , n18157 , n18161 );
and ( n18163 , n13322 , n771 );
and ( n18164 , n14118 , n719 );
xor ( n18165 , n18163 , n18164 );
and ( n18166 , n14938 , n663 );
xor ( n18167 , n18165 , n18166 );
xor ( n18168 , n18162 , n18167 );
xor ( n18169 , n18153 , n18168 );
xor ( n18170 , n18135 , n18169 );
xor ( n18171 , n18129 , n18170 );
and ( n18172 , n17459 , n17463 );
and ( n18173 , n17463 , n17480 );
and ( n18174 , n17459 , n17480 );
or ( n18175 , n18172 , n18173 , n18174 );
and ( n18176 , n17246 , n17261 );
and ( n18177 , n17261 , n17278 );
and ( n18178 , n17246 , n17278 );
or ( n18179 , n18176 , n18177 , n18178 );
xor ( n18180 , n18175 , n18179 );
and ( n18181 , n17468 , n17473 );
and ( n18182 , n17473 , n17479 );
and ( n18183 , n17468 , n17479 );
or ( n18184 , n18181 , n18182 , n18183 );
and ( n18185 , n17250 , n17254 );
and ( n18186 , n17254 , n17260 );
and ( n18187 , n17250 , n17260 );
or ( n18188 , n18185 , n18186 , n18187 );
xor ( n18189 , n18184 , n18188 );
and ( n18190 , n17475 , n17476 );
and ( n18191 , n17476 , n17478 );
and ( n18192 , n17475 , n17478 );
or ( n18193 , n18190 , n18191 , n18192 );
and ( n18194 , n11015 , n1034 );
and ( n18195 , n11769 , n940 );
xor ( n18196 , n18194 , n18195 );
and ( n18197 , n12320 , n840 );
xor ( n18198 , n18196 , n18197 );
xor ( n18199 , n18193 , n18198 );
and ( n18200 , n8718 , n1424 );
and ( n18201 , n9400 , n1254 );
xor ( n18202 , n18200 , n18201 );
and ( n18203 , n10291 , n1134 );
xor ( n18204 , n18202 , n18203 );
xor ( n18205 , n18199 , n18204 );
xor ( n18206 , n18189 , n18205 );
xor ( n18207 , n18180 , n18206 );
xor ( n18208 , n18171 , n18207 );
xor ( n18209 , n18125 , n18208 );
xor ( n18210 , n18116 , n18209 );
and ( n18211 , n17312 , n17359 );
and ( n18212 , n17359 , n17430 );
and ( n18213 , n17312 , n17430 );
or ( n18214 , n18211 , n18212 , n18213 );
and ( n18215 , n17242 , n17279 );
and ( n18216 , n17279 , n17305 );
and ( n18217 , n17242 , n17305 );
or ( n18218 , n18215 , n18216 , n18217 );
and ( n18219 , n17316 , n17320 );
and ( n18220 , n17320 , n17358 );
and ( n18221 , n17316 , n17358 );
or ( n18222 , n18219 , n18220 , n18221 );
xor ( n18223 , n18218 , n18222 );
and ( n18224 , n17284 , n17288 );
and ( n18225 , n17288 , n17304 );
and ( n18226 , n17284 , n17304 );
or ( n18227 , n18224 , n18225 , n18226 );
and ( n18228 , n17266 , n17271 );
and ( n18229 , n17271 , n17277 );
and ( n18230 , n17266 , n17277 );
or ( n18231 , n18228 , n18229 , n18230 );
and ( n18232 , n17256 , n17257 );
and ( n18233 , n17257 , n17259 );
and ( n18234 , n17256 , n17259 );
or ( n18235 , n18232 , n18233 , n18234 );
and ( n18236 , n17267 , n17268 );
and ( n18237 , n17268 , n17270 );
and ( n18238 , n17267 , n17270 );
or ( n18239 , n18236 , n18237 , n18238 );
xor ( n18240 , n18235 , n18239 );
and ( n18241 , n7385 , n1882 );
and ( n18242 , n7808 , n1738 );
xor ( n18243 , n18241 , n18242 );
and ( n18244 , n8079 , n1551 );
xor ( n18245 , n18243 , n18244 );
xor ( n18246 , n18240 , n18245 );
xor ( n18247 , n18231 , n18246 );
and ( n18248 , n17273 , n17274 );
and ( n18249 , n17274 , n17276 );
and ( n18250 , n17273 , n17276 );
or ( n18251 , n18248 , n18249 , n18250 );
and ( n18252 , n6187 , n2544 );
and ( n18253 , n6569 , n2298 );
xor ( n18254 , n18252 , n18253 );
and ( n18255 , n6816 , n2100 );
xor ( n18256 , n18254 , n18255 );
xor ( n18257 , n18251 , n18256 );
and ( n18258 , n4959 , n3271 );
and ( n18259 , n5459 , n2981 );
xor ( n18260 , n18258 , n18259 );
and ( n18261 , n5819 , n2739 );
xor ( n18262 , n18260 , n18261 );
xor ( n18263 , n18257 , n18262 );
xor ( n18264 , n18247 , n18263 );
xor ( n18265 , n18227 , n18264 );
and ( n18266 , n17293 , n17297 );
and ( n18267 , n17297 , n17303 );
and ( n18268 , n17293 , n17303 );
or ( n18269 , n18266 , n18267 , n18268 );
and ( n18270 , n17329 , n17334 );
and ( n18271 , n17334 , n17340 );
and ( n18272 , n17329 , n17340 );
or ( n18273 , n18270 , n18271 , n18272 );
xor ( n18274 , n18269 , n18273 );
and ( n18275 , n17299 , n17300 );
and ( n18276 , n17300 , n17302 );
and ( n18277 , n17299 , n17302 );
or ( n18278 , n18275 , n18276 , n18277 );
and ( n18279 , n17330 , n17331 );
and ( n18280 , n17331 , n17333 );
and ( n18281 , n17330 , n17333 );
or ( n18282 , n18279 , n18280 , n18281 );
xor ( n18283 , n18278 , n18282 );
buf ( n18284 , n4132 );
and ( n18285 , n4438 , n3749 );
xor ( n18286 , n18284 , n18285 );
and ( n18287 , n4766 , n3495 );
xor ( n18288 , n18286 , n18287 );
xor ( n18289 , n18283 , n18288 );
xor ( n18290 , n18274 , n18289 );
xor ( n18291 , n18265 , n18290 );
xor ( n18292 , n18223 , n18291 );
xor ( n18293 , n18214 , n18292 );
and ( n18294 , n17364 , n17390 );
and ( n18295 , n17390 , n17429 );
and ( n18296 , n17364 , n17429 );
or ( n18297 , n18294 , n18295 , n18296 );
and ( n18298 , n17325 , n17341 );
and ( n18299 , n17341 , n17357 );
and ( n18300 , n17325 , n17357 );
or ( n18301 , n18298 , n18299 , n18300 );
and ( n18302 , n17368 , n17372 );
and ( n18303 , n17372 , n17389 );
and ( n18304 , n17368 , n17389 );
or ( n18305 , n18302 , n18303 , n18304 );
xor ( n18306 , n18301 , n18305 );
and ( n18307 , n17346 , n17350 );
and ( n18308 , n17350 , n17356 );
and ( n18309 , n17346 , n17356 );
or ( n18310 , n18307 , n18308 , n18309 );
and ( n18311 , n17336 , n17337 );
and ( n18312 , n17337 , n17339 );
and ( n18313 , n17336 , n17339 );
or ( n18314 , n18311 , n18312 , n18313 );
and ( n18315 , n3182 , n5103 );
and ( n18316 , n3545 , n4730 );
xor ( n18317 , n18315 , n18316 );
and ( n18318 , n3801 , n4403 );
xor ( n18319 , n18317 , n18318 );
xor ( n18320 , n18314 , n18319 );
and ( n18321 , n2462 , n6132 );
and ( n18322 , n2779 , n5765 );
xor ( n18323 , n18321 , n18322 );
and ( n18324 , n3024 , n5408 );
xor ( n18325 , n18323 , n18324 );
xor ( n18326 , n18320 , n18325 );
xor ( n18327 , n18310 , n18326 );
and ( n18328 , n17352 , n17353 );
and ( n18329 , n17353 , n17355 );
and ( n18330 , n17352 , n17355 );
or ( n18331 , n18328 , n18329 , n18330 );
and ( n18332 , n17378 , n17379 );
and ( n18333 , n17379 , n17381 );
and ( n18334 , n17378 , n17381 );
or ( n18335 , n18332 , n18333 , n18334 );
xor ( n18336 , n18331 , n18335 );
and ( n18337 , n1933 , n7310 );
and ( n18338 , n2120 , n6971 );
xor ( n18339 , n18337 , n18338 );
and ( n18340 , n2324 , n6504 );
xor ( n18341 , n18339 , n18340 );
xor ( n18342 , n18336 , n18341 );
xor ( n18343 , n18327 , n18342 );
xor ( n18344 , n18306 , n18343 );
xor ( n18345 , n18297 , n18344 );
and ( n18346 , n17395 , n17410 );
and ( n18347 , n17410 , n17428 );
and ( n18348 , n17395 , n17428 );
or ( n18349 , n18346 , n18347 , n18348 );
and ( n18350 , n17377 , n17382 );
and ( n18351 , n17382 , n17388 );
and ( n18352 , n17377 , n17388 );
or ( n18353 , n18350 , n18351 , n18352 );
and ( n18354 , n17399 , n17403 );
and ( n18355 , n17403 , n17409 );
and ( n18356 , n17399 , n17409 );
or ( n18357 , n18354 , n18355 , n18356 );
xor ( n18358 , n18353 , n18357 );
and ( n18359 , n17384 , n17385 );
and ( n18360 , n17385 , n17387 );
and ( n18361 , n17384 , n17387 );
or ( n18362 , n18359 , n18360 , n18361 );
and ( n18363 , n1383 , n8669 );
and ( n18364 , n1580 , n8243 );
xor ( n18365 , n18363 , n18364 );
and ( n18366 , n1694 , n7662 );
xor ( n18367 , n18365 , n18366 );
xor ( n18368 , n18362 , n18367 );
and ( n18369 , n1047 , n10977 );
and ( n18370 , n1164 , n10239 );
xor ( n18371 , n18369 , n18370 );
and ( n18372 , n1287 , n9348 );
xor ( n18373 , n18371 , n18372 );
xor ( n18374 , n18368 , n18373 );
xor ( n18375 , n18358 , n18374 );
xor ( n18376 , n18349 , n18375 );
and ( n18377 , n17415 , n17420 );
and ( n18378 , n17420 , n17427 );
and ( n18379 , n17415 , n17427 );
or ( n18380 , n18377 , n18378 , n18379 );
and ( n18381 , n17405 , n17406 );
and ( n18382 , n17406 , n17408 );
and ( n18383 , n17405 , n17408 );
or ( n18384 , n18381 , n18382 , n18383 );
and ( n18385 , n17416 , n17417 );
and ( n18386 , n17417 , n17419 );
and ( n18387 , n17416 , n17419 );
or ( n18388 , n18385 , n18386 , n18387 );
xor ( n18389 , n18384 , n18388 );
and ( n18390 , n783 , n13256 );
and ( n18391 , n856 , n12531 );
xor ( n18392 , n18390 , n18391 );
and ( n18393 , n925 , n11718 );
xor ( n18394 , n18392 , n18393 );
xor ( n18395 , n18389 , n18394 );
xor ( n18396 , n18380 , n18395 );
and ( n18397 , n17423 , n17424 );
and ( n18398 , n17424 , n17426 );
and ( n18399 , n17423 , n17426 );
or ( n18400 , n18397 , n18398 , n18399 );
and ( n18401 , n632 , n15691 );
and ( n18402 , n671 , n14838 );
xor ( n18403 , n18401 , n18402 );
and ( n18404 , n715 , n14044 );
xor ( n18405 , n18403 , n18404 );
xor ( n18406 , n18400 , n18405 );
buf ( n18407 , n422 );
and ( n18408 , n599 , n18407 );
and ( n18409 , n608 , n17422 );
xor ( n18410 , n18408 , n18409 );
and ( n18411 , n611 , n16550 );
xor ( n18412 , n18410 , n18411 );
xor ( n18413 , n18406 , n18412 );
xor ( n18414 , n18396 , n18413 );
xor ( n18415 , n18376 , n18414 );
xor ( n18416 , n18345 , n18415 );
xor ( n18417 , n18293 , n18416 );
xor ( n18418 , n18210 , n18417 );
xor ( n18419 , n18112 , n18418 );
and ( n18420 , n17487 , n17516 );
and ( n18421 , n17437 , n17441 );
and ( n18422 , n17441 , n17518 );
and ( n18423 , n17437 , n17518 );
or ( n18424 , n18421 , n18422 , n18423 );
xor ( n18425 , n18420 , n18424 );
xor ( n18426 , n18419 , n18425 );
xor ( n18427 , n18108 , n18426 );
and ( n18428 , n17212 , n17216 );
and ( n18429 , n17216 , n17528 );
and ( n18430 , n17212 , n17528 );
or ( n18431 , n18428 , n18429 , n18430 );
xor ( n18432 , n18427 , n18431 );
and ( n18433 , n17529 , n17533 );
and ( n18434 , n17534 , n17535 );
or ( n18435 , n18433 , n18434 );
xor ( n18436 , n18432 , n18435 );
buf ( n18437 , n18436 );
buf ( n18438 , n18437 );
not ( n18439 , n18438 );
nor ( n18440 , n18439 , n8739 );
xor ( n18441 , n18102 , n18440 );
and ( n18442 , n17211 , n17540 );
and ( n18443 , n17541 , n17544 );
or ( n18444 , n18442 , n18443 );
xor ( n18445 , n18441 , n18444 );
buf ( n18446 , n18445 );
buf ( n18447 , n18446 );
not ( n18448 , n18447 );
buf ( n18449 , n547 );
not ( n18450 , n18449 );
nor ( n18451 , n18448 , n18450 );
xor ( n18452 , n17826 , n18451 );
xor ( n18453 , n17556 , n17823 );
nor ( n18454 , n17548 , n18450 );
and ( n18455 , n18453 , n18454 );
xor ( n18456 , n18453 , n18454 );
xor ( n18457 , n17560 , n17821 );
nor ( n18458 , n16669 , n18450 );
and ( n18459 , n18457 , n18458 );
xor ( n18460 , n18457 , n18458 );
xor ( n18461 , n17564 , n17819 );
nor ( n18462 , n15809 , n18450 );
and ( n18463 , n18461 , n18462 );
xor ( n18464 , n18461 , n18462 );
xor ( n18465 , n17568 , n17817 );
nor ( n18466 , n14968 , n18450 );
and ( n18467 , n18465 , n18466 );
xor ( n18468 , n18465 , n18466 );
xor ( n18469 , n17572 , n17815 );
nor ( n18470 , n14147 , n18450 );
and ( n18471 , n18469 , n18470 );
xor ( n18472 , n18469 , n18470 );
xor ( n18473 , n17576 , n17813 );
nor ( n18474 , n13349 , n18450 );
and ( n18475 , n18473 , n18474 );
xor ( n18476 , n18473 , n18474 );
xor ( n18477 , n17580 , n17811 );
nor ( n18478 , n12564 , n18450 );
and ( n18479 , n18477 , n18478 );
xor ( n18480 , n18477 , n18478 );
xor ( n18481 , n17584 , n17809 );
nor ( n18482 , n11799 , n18450 );
and ( n18483 , n18481 , n18482 );
xor ( n18484 , n18481 , n18482 );
xor ( n18485 , n17588 , n17807 );
nor ( n18486 , n11050 , n18450 );
and ( n18487 , n18485 , n18486 );
xor ( n18488 , n18485 , n18486 );
xor ( n18489 , n17592 , n17805 );
nor ( n18490 , n10321 , n18450 );
and ( n18491 , n18489 , n18490 );
xor ( n18492 , n18489 , n18490 );
xor ( n18493 , n17596 , n17803 );
nor ( n18494 , n9429 , n18450 );
and ( n18495 , n18493 , n18494 );
xor ( n18496 , n18493 , n18494 );
xor ( n18497 , n17600 , n17801 );
nor ( n18498 , n8949 , n18450 );
and ( n18499 , n18497 , n18498 );
xor ( n18500 , n18497 , n18498 );
xor ( n18501 , n17604 , n17799 );
nor ( n18502 , n9437 , n18450 );
and ( n18503 , n18501 , n18502 );
xor ( n18504 , n18501 , n18502 );
xor ( n18505 , n17608 , n17797 );
nor ( n18506 , n9446 , n18450 );
and ( n18507 , n18505 , n18506 );
xor ( n18508 , n18505 , n18506 );
xor ( n18509 , n17612 , n17795 );
nor ( n18510 , n9455 , n18450 );
and ( n18511 , n18509 , n18510 );
xor ( n18512 , n18509 , n18510 );
xor ( n18513 , n17616 , n17793 );
nor ( n18514 , n9464 , n18450 );
and ( n18515 , n18513 , n18514 );
xor ( n18516 , n18513 , n18514 );
xor ( n18517 , n17620 , n17791 );
nor ( n18518 , n9473 , n18450 );
and ( n18519 , n18517 , n18518 );
xor ( n18520 , n18517 , n18518 );
xor ( n18521 , n17624 , n17789 );
nor ( n18522 , n9482 , n18450 );
and ( n18523 , n18521 , n18522 );
xor ( n18524 , n18521 , n18522 );
xor ( n18525 , n17628 , n17787 );
nor ( n18526 , n9491 , n18450 );
and ( n18527 , n18525 , n18526 );
xor ( n18528 , n18525 , n18526 );
xor ( n18529 , n17632 , n17785 );
nor ( n18530 , n9500 , n18450 );
and ( n18531 , n18529 , n18530 );
xor ( n18532 , n18529 , n18530 );
xor ( n18533 , n17636 , n17783 );
nor ( n18534 , n9509 , n18450 );
and ( n18535 , n18533 , n18534 );
xor ( n18536 , n18533 , n18534 );
xor ( n18537 , n17640 , n17781 );
nor ( n18538 , n9518 , n18450 );
and ( n18539 , n18537 , n18538 );
xor ( n18540 , n18537 , n18538 );
xor ( n18541 , n17644 , n17779 );
nor ( n18542 , n9527 , n18450 );
and ( n18543 , n18541 , n18542 );
xor ( n18544 , n18541 , n18542 );
xor ( n18545 , n17648 , n17777 );
nor ( n18546 , n9536 , n18450 );
and ( n18547 , n18545 , n18546 );
xor ( n18548 , n18545 , n18546 );
xor ( n18549 , n17652 , n17775 );
nor ( n18550 , n9545 , n18450 );
and ( n18551 , n18549 , n18550 );
xor ( n18552 , n18549 , n18550 );
xor ( n18553 , n17656 , n17773 );
nor ( n18554 , n9554 , n18450 );
and ( n18555 , n18553 , n18554 );
xor ( n18556 , n18553 , n18554 );
xor ( n18557 , n17660 , n17771 );
nor ( n18558 , n9563 , n18450 );
and ( n18559 , n18557 , n18558 );
xor ( n18560 , n18557 , n18558 );
xor ( n18561 , n17664 , n17769 );
nor ( n18562 , n9572 , n18450 );
and ( n18563 , n18561 , n18562 );
xor ( n18564 , n18561 , n18562 );
xor ( n18565 , n17668 , n17767 );
nor ( n18566 , n9581 , n18450 );
and ( n18567 , n18565 , n18566 );
xor ( n18568 , n18565 , n18566 );
xor ( n18569 , n17672 , n17765 );
nor ( n18570 , n9590 , n18450 );
and ( n18571 , n18569 , n18570 );
xor ( n18572 , n18569 , n18570 );
xor ( n18573 , n17676 , n17763 );
nor ( n18574 , n9599 , n18450 );
and ( n18575 , n18573 , n18574 );
xor ( n18576 , n18573 , n18574 );
xor ( n18577 , n17680 , n17761 );
nor ( n18578 , n9608 , n18450 );
and ( n18579 , n18577 , n18578 );
xor ( n18580 , n18577 , n18578 );
xor ( n18581 , n17684 , n17759 );
nor ( n18582 , n9617 , n18450 );
and ( n18583 , n18581 , n18582 );
xor ( n18584 , n18581 , n18582 );
xor ( n18585 , n17688 , n17757 );
nor ( n18586 , n9626 , n18450 );
and ( n18587 , n18585 , n18586 );
xor ( n18588 , n18585 , n18586 );
xor ( n18589 , n17692 , n17755 );
nor ( n18590 , n9635 , n18450 );
and ( n18591 , n18589 , n18590 );
xor ( n18592 , n18589 , n18590 );
xor ( n18593 , n17696 , n17753 );
nor ( n18594 , n9644 , n18450 );
and ( n18595 , n18593 , n18594 );
xor ( n18596 , n18593 , n18594 );
xor ( n18597 , n17700 , n17751 );
nor ( n18598 , n9653 , n18450 );
and ( n18599 , n18597 , n18598 );
xor ( n18600 , n18597 , n18598 );
xor ( n18601 , n17704 , n17749 );
nor ( n18602 , n9662 , n18450 );
and ( n18603 , n18601 , n18602 );
xor ( n18604 , n18601 , n18602 );
xor ( n18605 , n17708 , n17747 );
nor ( n18606 , n9671 , n18450 );
and ( n18607 , n18605 , n18606 );
xor ( n18608 , n18605 , n18606 );
xor ( n18609 , n17712 , n17745 );
nor ( n18610 , n9680 , n18450 );
and ( n18611 , n18609 , n18610 );
xor ( n18612 , n18609 , n18610 );
xor ( n18613 , n17716 , n17743 );
nor ( n18614 , n9689 , n18450 );
and ( n18615 , n18613 , n18614 );
xor ( n18616 , n18613 , n18614 );
xor ( n18617 , n17720 , n17741 );
nor ( n18618 , n9698 , n18450 );
and ( n18619 , n18617 , n18618 );
xor ( n18620 , n18617 , n18618 );
xor ( n18621 , n17724 , n17739 );
nor ( n18622 , n9707 , n18450 );
and ( n18623 , n18621 , n18622 );
xor ( n18624 , n18621 , n18622 );
xor ( n18625 , n17728 , n17737 );
nor ( n18626 , n9716 , n18450 );
and ( n18627 , n18625 , n18626 );
xor ( n18628 , n18625 , n18626 );
xor ( n18629 , n17732 , n17735 );
nor ( n18630 , n9725 , n18450 );
and ( n18631 , n18629 , n18630 );
xor ( n18632 , n18629 , n18630 );
xor ( n18633 , n17733 , n17734 );
nor ( n18634 , n9734 , n18450 );
and ( n18635 , n18633 , n18634 );
xor ( n18636 , n18633 , n18634 );
nor ( n18637 , n9752 , n17550 );
nor ( n18638 , n9743 , n18450 );
and ( n18639 , n18637 , n18638 );
and ( n18640 , n18636 , n18639 );
or ( n18641 , n18635 , n18640 );
and ( n18642 , n18632 , n18641 );
or ( n18643 , n18631 , n18642 );
and ( n18644 , n18628 , n18643 );
or ( n18645 , n18627 , n18644 );
and ( n18646 , n18624 , n18645 );
or ( n18647 , n18623 , n18646 );
and ( n18648 , n18620 , n18647 );
or ( n18649 , n18619 , n18648 );
and ( n18650 , n18616 , n18649 );
or ( n18651 , n18615 , n18650 );
and ( n18652 , n18612 , n18651 );
or ( n18653 , n18611 , n18652 );
and ( n18654 , n18608 , n18653 );
or ( n18655 , n18607 , n18654 );
and ( n18656 , n18604 , n18655 );
or ( n18657 , n18603 , n18656 );
and ( n18658 , n18600 , n18657 );
or ( n18659 , n18599 , n18658 );
and ( n18660 , n18596 , n18659 );
or ( n18661 , n18595 , n18660 );
and ( n18662 , n18592 , n18661 );
or ( n18663 , n18591 , n18662 );
and ( n18664 , n18588 , n18663 );
or ( n18665 , n18587 , n18664 );
and ( n18666 , n18584 , n18665 );
or ( n18667 , n18583 , n18666 );
and ( n18668 , n18580 , n18667 );
or ( n18669 , n18579 , n18668 );
and ( n18670 , n18576 , n18669 );
or ( n18671 , n18575 , n18670 );
and ( n18672 , n18572 , n18671 );
or ( n18673 , n18571 , n18672 );
and ( n18674 , n18568 , n18673 );
or ( n18675 , n18567 , n18674 );
and ( n18676 , n18564 , n18675 );
or ( n18677 , n18563 , n18676 );
and ( n18678 , n18560 , n18677 );
or ( n18679 , n18559 , n18678 );
and ( n18680 , n18556 , n18679 );
or ( n18681 , n18555 , n18680 );
and ( n18682 , n18552 , n18681 );
or ( n18683 , n18551 , n18682 );
and ( n18684 , n18548 , n18683 );
or ( n18685 , n18547 , n18684 );
and ( n18686 , n18544 , n18685 );
or ( n18687 , n18543 , n18686 );
and ( n18688 , n18540 , n18687 );
or ( n18689 , n18539 , n18688 );
and ( n18690 , n18536 , n18689 );
or ( n18691 , n18535 , n18690 );
and ( n18692 , n18532 , n18691 );
or ( n18693 , n18531 , n18692 );
and ( n18694 , n18528 , n18693 );
or ( n18695 , n18527 , n18694 );
and ( n18696 , n18524 , n18695 );
or ( n18697 , n18523 , n18696 );
and ( n18698 , n18520 , n18697 );
or ( n18699 , n18519 , n18698 );
and ( n18700 , n18516 , n18699 );
or ( n18701 , n18515 , n18700 );
and ( n18702 , n18512 , n18701 );
or ( n18703 , n18511 , n18702 );
and ( n18704 , n18508 , n18703 );
or ( n18705 , n18507 , n18704 );
and ( n18706 , n18504 , n18705 );
or ( n18707 , n18503 , n18706 );
and ( n18708 , n18500 , n18707 );
or ( n18709 , n18499 , n18708 );
and ( n18710 , n18496 , n18709 );
or ( n18711 , n18495 , n18710 );
and ( n18712 , n18492 , n18711 );
or ( n18713 , n18491 , n18712 );
and ( n18714 , n18488 , n18713 );
or ( n18715 , n18487 , n18714 );
and ( n18716 , n18484 , n18715 );
or ( n18717 , n18483 , n18716 );
and ( n18718 , n18480 , n18717 );
or ( n18719 , n18479 , n18718 );
and ( n18720 , n18476 , n18719 );
or ( n18721 , n18475 , n18720 );
and ( n18722 , n18472 , n18721 );
or ( n18723 , n18471 , n18722 );
and ( n18724 , n18468 , n18723 );
or ( n18725 , n18467 , n18724 );
and ( n18726 , n18464 , n18725 );
or ( n18727 , n18463 , n18726 );
and ( n18728 , n18460 , n18727 );
or ( n18729 , n18459 , n18728 );
and ( n18730 , n18456 , n18729 );
or ( n18731 , n18455 , n18730 );
xor ( n18732 , n18452 , n18731 );
buf ( n18733 , n485 );
not ( n18734 , n18733 );
nor ( n18735 , n601 , n18734 );
buf ( n18736 , n18735 );
nor ( n18737 , n622 , n16943 );
xor ( n18738 , n18736 , n18737 );
buf ( n18739 , n18738 );
nor ( n18740 , n646 , n16077 );
xor ( n18741 , n18739 , n18740 );
and ( n18742 , n17830 , n17831 );
buf ( n18743 , n18742 );
xor ( n18744 , n18741 , n18743 );
nor ( n18745 , n684 , n15230 );
xor ( n18746 , n18744 , n18745 );
and ( n18747 , n17833 , n17834 );
and ( n18748 , n17835 , n17837 );
or ( n18749 , n18747 , n18748 );
xor ( n18750 , n18746 , n18749 );
nor ( n18751 , n733 , n14403 );
xor ( n18752 , n18750 , n18751 );
and ( n18753 , n17838 , n17839 );
and ( n18754 , n17840 , n17843 );
or ( n18755 , n18753 , n18754 );
xor ( n18756 , n18752 , n18755 );
nor ( n18757 , n796 , n13599 );
xor ( n18758 , n18756 , n18757 );
and ( n18759 , n17844 , n17845 );
and ( n18760 , n17846 , n17849 );
or ( n18761 , n18759 , n18760 );
xor ( n18762 , n18758 , n18761 );
nor ( n18763 , n868 , n12808 );
xor ( n18764 , n18762 , n18763 );
and ( n18765 , n17850 , n17851 );
and ( n18766 , n17852 , n17855 );
or ( n18767 , n18765 , n18766 );
xor ( n18768 , n18764 , n18767 );
nor ( n18769 , n958 , n12037 );
xor ( n18770 , n18768 , n18769 );
and ( n18771 , n17856 , n17857 );
and ( n18772 , n17858 , n17861 );
or ( n18773 , n18771 , n18772 );
xor ( n18774 , n18770 , n18773 );
nor ( n18775 , n1062 , n11282 );
xor ( n18776 , n18774 , n18775 );
and ( n18777 , n17862 , n17863 );
and ( n18778 , n17864 , n17867 );
or ( n18779 , n18777 , n18778 );
xor ( n18780 , n18776 , n18779 );
nor ( n18781 , n1176 , n10547 );
xor ( n18782 , n18780 , n18781 );
and ( n18783 , n17868 , n17869 );
and ( n18784 , n17870 , n17873 );
or ( n18785 , n18783 , n18784 );
xor ( n18786 , n18782 , n18785 );
nor ( n18787 , n1303 , n9829 );
xor ( n18788 , n18786 , n18787 );
and ( n18789 , n17874 , n17875 );
and ( n18790 , n17876 , n17879 );
or ( n18791 , n18789 , n18790 );
xor ( n18792 , n18788 , n18791 );
nor ( n18793 , n1445 , n8955 );
xor ( n18794 , n18792 , n18793 );
and ( n18795 , n17880 , n17881 );
and ( n18796 , n17882 , n17885 );
or ( n18797 , n18795 , n18796 );
xor ( n18798 , n18794 , n18797 );
nor ( n18799 , n1598 , n603 );
xor ( n18800 , n18798 , n18799 );
and ( n18801 , n17886 , n17887 );
and ( n18802 , n17888 , n17891 );
or ( n18803 , n18801 , n18802 );
xor ( n18804 , n18800 , n18803 );
nor ( n18805 , n1766 , n652 );
xor ( n18806 , n18804 , n18805 );
and ( n18807 , n17892 , n17893 );
and ( n18808 , n17894 , n17897 );
or ( n18809 , n18807 , n18808 );
xor ( n18810 , n18806 , n18809 );
nor ( n18811 , n1945 , n624 );
xor ( n18812 , n18810 , n18811 );
and ( n18813 , n17898 , n17899 );
and ( n18814 , n17900 , n17903 );
or ( n18815 , n18813 , n18814 );
xor ( n18816 , n18812 , n18815 );
nor ( n18817 , n2137 , n648 );
xor ( n18818 , n18816 , n18817 );
and ( n18819 , n17904 , n17905 );
and ( n18820 , n17906 , n17909 );
or ( n18821 , n18819 , n18820 );
xor ( n18822 , n18818 , n18821 );
nor ( n18823 , n2343 , n686 );
xor ( n18824 , n18822 , n18823 );
and ( n18825 , n17910 , n17911 );
and ( n18826 , n17912 , n17915 );
or ( n18827 , n18825 , n18826 );
xor ( n18828 , n18824 , n18827 );
nor ( n18829 , n2566 , n735 );
xor ( n18830 , n18828 , n18829 );
and ( n18831 , n17916 , n17917 );
and ( n18832 , n17918 , n17921 );
or ( n18833 , n18831 , n18832 );
xor ( n18834 , n18830 , n18833 );
nor ( n18835 , n2797 , n798 );
xor ( n18836 , n18834 , n18835 );
and ( n18837 , n17922 , n17923 );
and ( n18838 , n17924 , n17927 );
or ( n18839 , n18837 , n18838 );
xor ( n18840 , n18836 , n18839 );
nor ( n18841 , n3043 , n870 );
xor ( n18842 , n18840 , n18841 );
and ( n18843 , n17928 , n17929 );
and ( n18844 , n17930 , n17933 );
or ( n18845 , n18843 , n18844 );
xor ( n18846 , n18842 , n18845 );
nor ( n18847 , n3300 , n960 );
xor ( n18848 , n18846 , n18847 );
and ( n18849 , n17934 , n17935 );
and ( n18850 , n17936 , n17939 );
or ( n18851 , n18849 , n18850 );
xor ( n18852 , n18848 , n18851 );
nor ( n18853 , n3570 , n1064 );
xor ( n18854 , n18852 , n18853 );
and ( n18855 , n17940 , n17941 );
and ( n18856 , n17942 , n17945 );
or ( n18857 , n18855 , n18856 );
xor ( n18858 , n18854 , n18857 );
nor ( n18859 , n3853 , n1178 );
xor ( n18860 , n18858 , n18859 );
and ( n18861 , n17946 , n17947 );
and ( n18862 , n17948 , n17951 );
or ( n18863 , n18861 , n18862 );
xor ( n18864 , n18860 , n18863 );
nor ( n18865 , n4151 , n1305 );
xor ( n18866 , n18864 , n18865 );
and ( n18867 , n17952 , n17953 );
and ( n18868 , n17954 , n17957 );
or ( n18869 , n18867 , n18868 );
xor ( n18870 , n18866 , n18869 );
nor ( n18871 , n4458 , n1447 );
xor ( n18872 , n18870 , n18871 );
and ( n18873 , n17958 , n17959 );
and ( n18874 , n17960 , n17963 );
or ( n18875 , n18873 , n18874 );
xor ( n18876 , n18872 , n18875 );
nor ( n18877 , n4786 , n1600 );
xor ( n18878 , n18876 , n18877 );
and ( n18879 , n17964 , n17965 );
and ( n18880 , n17966 , n17969 );
or ( n18881 , n18879 , n18880 );
xor ( n18882 , n18878 , n18881 );
nor ( n18883 , n5126 , n1768 );
xor ( n18884 , n18882 , n18883 );
and ( n18885 , n17970 , n17971 );
and ( n18886 , n17972 , n17975 );
or ( n18887 , n18885 , n18886 );
xor ( n18888 , n18884 , n18887 );
nor ( n18889 , n5477 , n1947 );
xor ( n18890 , n18888 , n18889 );
and ( n18891 , n17976 , n17977 );
and ( n18892 , n17978 , n17981 );
or ( n18893 , n18891 , n18892 );
xor ( n18894 , n18890 , n18893 );
nor ( n18895 , n5838 , n2139 );
xor ( n18896 , n18894 , n18895 );
and ( n18897 , n17982 , n17983 );
and ( n18898 , n17984 , n17987 );
or ( n18899 , n18897 , n18898 );
xor ( n18900 , n18896 , n18899 );
nor ( n18901 , n6212 , n2345 );
xor ( n18902 , n18900 , n18901 );
and ( n18903 , n17988 , n17989 );
and ( n18904 , n17990 , n17993 );
or ( n18905 , n18903 , n18904 );
xor ( n18906 , n18902 , n18905 );
nor ( n18907 , n6596 , n2568 );
xor ( n18908 , n18906 , n18907 );
and ( n18909 , n17994 , n17995 );
and ( n18910 , n17996 , n17999 );
or ( n18911 , n18909 , n18910 );
xor ( n18912 , n18908 , n18911 );
nor ( n18913 , n6997 , n2799 );
xor ( n18914 , n18912 , n18913 );
and ( n18915 , n18000 , n18001 );
and ( n18916 , n18002 , n18005 );
or ( n18917 , n18915 , n18916 );
xor ( n18918 , n18914 , n18917 );
nor ( n18919 , n7413 , n3045 );
xor ( n18920 , n18918 , n18919 );
and ( n18921 , n18006 , n18007 );
and ( n18922 , n18008 , n18011 );
or ( n18923 , n18921 , n18922 );
xor ( n18924 , n18920 , n18923 );
nor ( n18925 , n7841 , n3302 );
xor ( n18926 , n18924 , n18925 );
and ( n18927 , n18012 , n18013 );
and ( n18928 , n18014 , n18017 );
or ( n18929 , n18927 , n18928 );
xor ( n18930 , n18926 , n18929 );
nor ( n18931 , n8281 , n3572 );
xor ( n18932 , n18930 , n18931 );
and ( n18933 , n18018 , n18019 );
and ( n18934 , n18020 , n18023 );
or ( n18935 , n18933 , n18934 );
xor ( n18936 , n18932 , n18935 );
nor ( n18937 , n8737 , n3855 );
xor ( n18938 , n18936 , n18937 );
and ( n18939 , n18024 , n18025 );
and ( n18940 , n18026 , n18029 );
or ( n18941 , n18939 , n18940 );
xor ( n18942 , n18938 , n18941 );
nor ( n18943 , n9420 , n4153 );
xor ( n18944 , n18942 , n18943 );
and ( n18945 , n18030 , n18031 );
and ( n18946 , n18032 , n18035 );
or ( n18947 , n18945 , n18946 );
xor ( n18948 , n18944 , n18947 );
nor ( n18949 , n10312 , n4460 );
xor ( n18950 , n18948 , n18949 );
and ( n18951 , n18036 , n18037 );
and ( n18952 , n18038 , n18041 );
or ( n18953 , n18951 , n18952 );
xor ( n18954 , n18950 , n18953 );
nor ( n18955 , n11041 , n4788 );
xor ( n18956 , n18954 , n18955 );
and ( n18957 , n18042 , n18043 );
and ( n18958 , n18044 , n18047 );
or ( n18959 , n18957 , n18958 );
xor ( n18960 , n18956 , n18959 );
nor ( n18961 , n11790 , n5128 );
xor ( n18962 , n18960 , n18961 );
and ( n18963 , n18048 , n18049 );
and ( n18964 , n18050 , n18053 );
or ( n18965 , n18963 , n18964 );
xor ( n18966 , n18962 , n18965 );
nor ( n18967 , n12555 , n5479 );
xor ( n18968 , n18966 , n18967 );
and ( n18969 , n18054 , n18055 );
and ( n18970 , n18056 , n18059 );
or ( n18971 , n18969 , n18970 );
xor ( n18972 , n18968 , n18971 );
nor ( n18973 , n13340 , n5840 );
xor ( n18974 , n18972 , n18973 );
and ( n18975 , n18060 , n18061 );
and ( n18976 , n18062 , n18065 );
or ( n18977 , n18975 , n18976 );
xor ( n18978 , n18974 , n18977 );
nor ( n18979 , n14138 , n6214 );
xor ( n18980 , n18978 , n18979 );
and ( n18981 , n18066 , n18067 );
and ( n18982 , n18068 , n18071 );
or ( n18983 , n18981 , n18982 );
xor ( n18984 , n18980 , n18983 );
nor ( n18985 , n14959 , n6598 );
xor ( n18986 , n18984 , n18985 );
and ( n18987 , n18072 , n18073 );
and ( n18988 , n18074 , n18077 );
or ( n18989 , n18987 , n18988 );
xor ( n18990 , n18986 , n18989 );
nor ( n18991 , n15800 , n6999 );
xor ( n18992 , n18990 , n18991 );
and ( n18993 , n18078 , n18079 );
and ( n18994 , n18080 , n18083 );
or ( n18995 , n18993 , n18994 );
xor ( n18996 , n18992 , n18995 );
nor ( n18997 , n16660 , n7415 );
xor ( n18998 , n18996 , n18997 );
and ( n18999 , n18084 , n18085 );
and ( n19000 , n18086 , n18089 );
or ( n19001 , n18999 , n19000 );
xor ( n19002 , n18998 , n19001 );
nor ( n19003 , n17539 , n7843 );
xor ( n19004 , n19002 , n19003 );
and ( n19005 , n18090 , n18091 );
and ( n19006 , n18092 , n18095 );
or ( n19007 , n19005 , n19006 );
xor ( n19008 , n19004 , n19007 );
nor ( n19009 , n18439 , n8283 );
xor ( n19010 , n19008 , n19009 );
and ( n19011 , n18096 , n18097 );
and ( n19012 , n18098 , n18101 );
or ( n19013 , n19011 , n19012 );
xor ( n19014 , n19010 , n19013 );
and ( n19015 , n18420 , n18424 );
and ( n19016 , n18112 , n18418 );
and ( n19017 , n18418 , n18425 );
and ( n19018 , n18112 , n18425 );
or ( n19019 , n19016 , n19017 , n19018 );
xor ( n19020 , n19015 , n19019 );
and ( n19021 , n18116 , n18209 );
and ( n19022 , n18209 , n18417 );
and ( n19023 , n18116 , n18417 );
or ( n19024 , n19021 , n19022 , n19023 );
and ( n19025 , n18214 , n18292 );
and ( n19026 , n18292 , n18416 );
and ( n19027 , n18214 , n18416 );
or ( n19028 , n19025 , n19026 , n19027 );
and ( n19029 , n18297 , n18344 );
and ( n19030 , n18344 , n18415 );
and ( n19031 , n18297 , n18415 );
or ( n19032 , n19029 , n19030 , n19031 );
and ( n19033 , n18227 , n18264 );
and ( n19034 , n18264 , n18290 );
and ( n19035 , n18227 , n18290 );
or ( n19036 , n19033 , n19034 , n19035 );
and ( n19037 , n18301 , n18305 );
and ( n19038 , n18305 , n18343 );
and ( n19039 , n18301 , n18343 );
or ( n19040 , n19037 , n19038 , n19039 );
xor ( n19041 , n19036 , n19040 );
and ( n19042 , n18269 , n18273 );
and ( n19043 , n18273 , n18289 );
and ( n19044 , n18269 , n18289 );
or ( n19045 , n19042 , n19043 , n19044 );
and ( n19046 , n18251 , n18256 );
and ( n19047 , n18256 , n18262 );
and ( n19048 , n18251 , n18262 );
or ( n19049 , n19046 , n19047 , n19048 );
and ( n19050 , n18241 , n18242 );
and ( n19051 , n18242 , n18244 );
and ( n19052 , n18241 , n18244 );
or ( n19053 , n19050 , n19051 , n19052 );
and ( n19054 , n18252 , n18253 );
and ( n19055 , n18253 , n18255 );
and ( n19056 , n18252 , n18255 );
or ( n19057 , n19054 , n19055 , n19056 );
xor ( n19058 , n19053 , n19057 );
and ( n19059 , n7385 , n2100 );
and ( n19060 , n7808 , n1882 );
xor ( n19061 , n19059 , n19060 );
and ( n19062 , n8079 , n1738 );
xor ( n19063 , n19061 , n19062 );
xor ( n19064 , n19058 , n19063 );
xor ( n19065 , n19049 , n19064 );
and ( n19066 , n18258 , n18259 );
and ( n19067 , n18259 , n18261 );
and ( n19068 , n18258 , n18261 );
or ( n19069 , n19066 , n19067 , n19068 );
and ( n19070 , n6187 , n2739 );
and ( n19071 , n6569 , n2544 );
xor ( n19072 , n19070 , n19071 );
and ( n19073 , n6816 , n2298 );
xor ( n19074 , n19072 , n19073 );
xor ( n19075 , n19069 , n19074 );
and ( n19076 , n4959 , n3495 );
and ( n19077 , n5459 , n3271 );
xor ( n19078 , n19076 , n19077 );
and ( n19079 , n5819 , n2981 );
xor ( n19080 , n19078 , n19079 );
xor ( n19081 , n19075 , n19080 );
xor ( n19082 , n19065 , n19081 );
xor ( n19083 , n19045 , n19082 );
and ( n19084 , n18278 , n18282 );
and ( n19085 , n18282 , n18288 );
and ( n19086 , n18278 , n18288 );
or ( n19087 , n19084 , n19085 , n19086 );
and ( n19088 , n18314 , n18319 );
and ( n19089 , n18319 , n18325 );
and ( n19090 , n18314 , n18325 );
or ( n19091 , n19088 , n19089 , n19090 );
xor ( n19092 , n19087 , n19091 );
and ( n19093 , n18284 , n18285 );
and ( n19094 , n18285 , n18287 );
and ( n19095 , n18284 , n18287 );
or ( n19096 , n19093 , n19094 , n19095 );
and ( n19097 , n18315 , n18316 );
and ( n19098 , n18316 , n18318 );
and ( n19099 , n18315 , n18318 );
or ( n19100 , n19097 , n19098 , n19099 );
xor ( n19101 , n19096 , n19100 );
and ( n19102 , n4766 , n3749 );
buf ( n19103 , n19102 );
xor ( n19104 , n19101 , n19103 );
xor ( n19105 , n19092 , n19104 );
xor ( n19106 , n19083 , n19105 );
xor ( n19107 , n19041 , n19106 );
xor ( n19108 , n19032 , n19107 );
and ( n19109 , n18349 , n18375 );
and ( n19110 , n18375 , n18414 );
and ( n19111 , n18349 , n18414 );
or ( n19112 , n19109 , n19110 , n19111 );
and ( n19113 , n18310 , n18326 );
and ( n19114 , n18326 , n18342 );
and ( n19115 , n18310 , n18342 );
or ( n19116 , n19113 , n19114 , n19115 );
and ( n19117 , n18353 , n18357 );
and ( n19118 , n18357 , n18374 );
and ( n19119 , n18353 , n18374 );
or ( n19120 , n19117 , n19118 , n19119 );
xor ( n19121 , n19116 , n19120 );
and ( n19122 , n18331 , n18335 );
and ( n19123 , n18335 , n18341 );
and ( n19124 , n18331 , n18341 );
or ( n19125 , n19122 , n19123 , n19124 );
and ( n19126 , n18321 , n18322 );
and ( n19127 , n18322 , n18324 );
and ( n19128 , n18321 , n18324 );
or ( n19129 , n19126 , n19127 , n19128 );
and ( n19130 , n3182 , n5408 );
and ( n19131 , n3545 , n5103 );
xor ( n19132 , n19130 , n19131 );
and ( n19133 , n3801 , n4730 );
xor ( n19134 , n19132 , n19133 );
xor ( n19135 , n19129 , n19134 );
and ( n19136 , n2462 , n6504 );
and ( n19137 , n2779 , n6132 );
xor ( n19138 , n19136 , n19137 );
and ( n19139 , n3024 , n5765 );
xor ( n19140 , n19138 , n19139 );
xor ( n19141 , n19135 , n19140 );
xor ( n19142 , n19125 , n19141 );
and ( n19143 , n18337 , n18338 );
and ( n19144 , n18338 , n18340 );
and ( n19145 , n18337 , n18340 );
or ( n19146 , n19143 , n19144 , n19145 );
and ( n19147 , n18363 , n18364 );
and ( n19148 , n18364 , n18366 );
and ( n19149 , n18363 , n18366 );
or ( n19150 , n19147 , n19148 , n19149 );
xor ( n19151 , n19146 , n19150 );
and ( n19152 , n1933 , n7662 );
and ( n19153 , n2120 , n7310 );
xor ( n19154 , n19152 , n19153 );
and ( n19155 , n2324 , n6971 );
xor ( n19156 , n19154 , n19155 );
xor ( n19157 , n19151 , n19156 );
xor ( n19158 , n19142 , n19157 );
xor ( n19159 , n19121 , n19158 );
xor ( n19160 , n19112 , n19159 );
and ( n19161 , n18380 , n18395 );
and ( n19162 , n18395 , n18413 );
and ( n19163 , n18380 , n18413 );
or ( n19164 , n19161 , n19162 , n19163 );
and ( n19165 , n18362 , n18367 );
and ( n19166 , n18367 , n18373 );
and ( n19167 , n18362 , n18373 );
or ( n19168 , n19165 , n19166 , n19167 );
and ( n19169 , n18384 , n18388 );
and ( n19170 , n18388 , n18394 );
and ( n19171 , n18384 , n18394 );
or ( n19172 , n19169 , n19170 , n19171 );
xor ( n19173 , n19168 , n19172 );
and ( n19174 , n18369 , n18370 );
and ( n19175 , n18370 , n18372 );
and ( n19176 , n18369 , n18372 );
or ( n19177 , n19174 , n19175 , n19176 );
and ( n19178 , n1383 , n9348 );
and ( n19179 , n1580 , n8669 );
xor ( n19180 , n19178 , n19179 );
and ( n19181 , n1694 , n8243 );
xor ( n19182 , n19180 , n19181 );
xor ( n19183 , n19177 , n19182 );
and ( n19184 , n1047 , n11718 );
and ( n19185 , n1164 , n10977 );
xor ( n19186 , n19184 , n19185 );
and ( n19187 , n1287 , n10239 );
xor ( n19188 , n19186 , n19187 );
xor ( n19189 , n19183 , n19188 );
xor ( n19190 , n19173 , n19189 );
xor ( n19191 , n19164 , n19190 );
and ( n19192 , n18400 , n18405 );
and ( n19193 , n18405 , n18412 );
and ( n19194 , n18400 , n18412 );
or ( n19195 , n19192 , n19193 , n19194 );
and ( n19196 , n18390 , n18391 );
and ( n19197 , n18391 , n18393 );
and ( n19198 , n18390 , n18393 );
or ( n19199 , n19196 , n19197 , n19198 );
and ( n19200 , n18401 , n18402 );
and ( n19201 , n18402 , n18404 );
and ( n19202 , n18401 , n18404 );
or ( n19203 , n19200 , n19201 , n19202 );
xor ( n19204 , n19199 , n19203 );
and ( n19205 , n783 , n14044 );
and ( n19206 , n856 , n13256 );
xor ( n19207 , n19205 , n19206 );
and ( n19208 , n925 , n12531 );
xor ( n19209 , n19207 , n19208 );
xor ( n19210 , n19204 , n19209 );
xor ( n19211 , n19195 , n19210 );
and ( n19212 , n18408 , n18409 );
and ( n19213 , n18409 , n18411 );
and ( n19214 , n18408 , n18411 );
or ( n19215 , n19212 , n19213 , n19214 );
and ( n19216 , n632 , n16550 );
and ( n19217 , n671 , n15691 );
xor ( n19218 , n19216 , n19217 );
and ( n19219 , n715 , n14838 );
xor ( n19220 , n19218 , n19219 );
xor ( n19221 , n19215 , n19220 );
buf ( n19222 , n421 );
and ( n19223 , n599 , n19222 );
and ( n19224 , n608 , n18407 );
xor ( n19225 , n19223 , n19224 );
and ( n19226 , n611 , n17422 );
xor ( n19227 , n19225 , n19226 );
xor ( n19228 , n19221 , n19227 );
xor ( n19229 , n19211 , n19228 );
xor ( n19230 , n19191 , n19229 );
xor ( n19231 , n19160 , n19230 );
xor ( n19232 , n19108 , n19231 );
xor ( n19233 , n19028 , n19232 );
and ( n19234 , n18129 , n18170 );
and ( n19235 , n18170 , n18207 );
and ( n19236 , n18129 , n18207 );
or ( n19237 , n19234 , n19235 , n19236 );
and ( n19238 , n18218 , n18222 );
and ( n19239 , n18222 , n18291 );
and ( n19240 , n18218 , n18291 );
or ( n19241 , n19238 , n19239 , n19240 );
xor ( n19242 , n19237 , n19241 );
and ( n19243 , n18175 , n18179 );
and ( n19244 , n18179 , n18206 );
and ( n19245 , n18175 , n18206 );
or ( n19246 , n19243 , n19244 , n19245 );
and ( n19247 , n18184 , n18188 );
and ( n19248 , n18188 , n18205 );
and ( n19249 , n18184 , n18205 );
or ( n19250 , n19247 , n19248 , n19249 );
and ( n19251 , n18231 , n18246 );
and ( n19252 , n18246 , n18263 );
and ( n19253 , n18231 , n18263 );
or ( n19254 , n19251 , n19252 , n19253 );
xor ( n19255 , n19250 , n19254 );
and ( n19256 , n18193 , n18198 );
and ( n19257 , n18198 , n18204 );
and ( n19258 , n18193 , n18204 );
or ( n19259 , n19256 , n19257 , n19258 );
and ( n19260 , n18235 , n18239 );
and ( n19261 , n18239 , n18245 );
and ( n19262 , n18235 , n18245 );
or ( n19263 , n19260 , n19261 , n19262 );
xor ( n19264 , n19259 , n19263 );
and ( n19265 , n18200 , n18201 );
and ( n19266 , n18201 , n18203 );
and ( n19267 , n18200 , n18203 );
or ( n19268 , n19265 , n19266 , n19267 );
and ( n19269 , n11015 , n1134 );
and ( n19270 , n11769 , n1034 );
xor ( n19271 , n19269 , n19270 );
and ( n19272 , n12320 , n940 );
xor ( n19273 , n19271 , n19272 );
xor ( n19274 , n19268 , n19273 );
and ( n19275 , n8718 , n1551 );
and ( n19276 , n9400 , n1424 );
xor ( n19277 , n19275 , n19276 );
and ( n19278 , n10291 , n1254 );
xor ( n19279 , n19277 , n19278 );
xor ( n19280 , n19274 , n19279 );
xor ( n19281 , n19264 , n19280 );
xor ( n19282 , n19255 , n19281 );
xor ( n19283 , n19246 , n19282 );
and ( n19284 , n18143 , n18145 );
and ( n19285 , n18145 , n18151 );
and ( n19286 , n18143 , n18151 );
or ( n19287 , n19284 , n19285 , n19286 );
and ( n19288 , n18139 , n18152 );
and ( n19289 , n18152 , n18168 );
and ( n19290 , n18139 , n18168 );
or ( n19291 , n19288 , n19289 , n19290 );
xor ( n19292 , n19287 , n19291 );
and ( n19293 , n18157 , n18161 );
and ( n19294 , n18161 , n18167 );
and ( n19295 , n18157 , n18167 );
or ( n19296 , n19293 , n19294 , n19295 );
and ( n19297 , n18163 , n18164 );
and ( n19298 , n18164 , n18166 );
and ( n19299 , n18163 , n18166 );
or ( n19300 , n19297 , n19298 , n19299 );
and ( n19301 , n18194 , n18195 );
and ( n19302 , n18195 , n18197 );
and ( n19303 , n18194 , n18197 );
or ( n19304 , n19301 , n19302 , n19303 );
xor ( n19305 , n19300 , n19304 );
and ( n19306 , n13322 , n840 );
and ( n19307 , n14118 , n771 );
xor ( n19308 , n19306 , n19307 );
and ( n19309 , n14938 , n719 );
xor ( n19310 , n19308 , n19309 );
xor ( n19311 , n19305 , n19310 );
xor ( n19312 , n19296 , n19311 );
and ( n19313 , n18147 , n18148 );
and ( n19314 , n18148 , n18150 );
and ( n19315 , n18147 , n18150 );
or ( n19316 , n19313 , n19314 , n19315 );
and ( n19317 , n15758 , n663 );
and ( n19318 , n16637 , n635 );
xor ( n19319 , n19317 , n19318 );
and ( n19320 , n17512 , n606 );
xor ( n19321 , n19319 , n19320 );
xor ( n19322 , n19316 , n19321 );
and ( n19323 , n18144 , n615 );
buf ( n19324 , n421 );
and ( n19325 , n19324 , n612 );
xor ( n19326 , n19323 , n19325 );
xor ( n19327 , n19322 , n19326 );
xor ( n19328 , n19312 , n19327 );
xor ( n19329 , n19292 , n19328 );
xor ( n19330 , n19283 , n19329 );
xor ( n19331 , n19242 , n19330 );
xor ( n19332 , n19233 , n19331 );
xor ( n19333 , n19024 , n19332 );
and ( n19334 , n18130 , n18134 );
and ( n19335 , n18134 , n18169 );
and ( n19336 , n18130 , n18169 );
or ( n19337 , n19334 , n19335 , n19336 );
and ( n19338 , n18120 , n18124 );
and ( n19339 , n18124 , n18208 );
and ( n19340 , n18120 , n18208 );
or ( n19341 , n19338 , n19339 , n19340 );
xor ( n19342 , n19337 , n19341 );
xor ( n19343 , n19333 , n19342 );
xor ( n19344 , n19020 , n19343 );
and ( n19345 , n18103 , n18107 );
and ( n19346 , n18107 , n18426 );
and ( n19347 , n18103 , n18426 );
or ( n19348 , n19345 , n19346 , n19347 );
xor ( n19349 , n19344 , n19348 );
and ( n19350 , n18427 , n18431 );
and ( n19351 , n18432 , n18435 );
or ( n19352 , n19350 , n19351 );
xor ( n19353 , n19349 , n19352 );
buf ( n19354 , n19353 );
buf ( n19355 , n19354 );
not ( n19356 , n19355 );
nor ( n19357 , n19356 , n8739 );
xor ( n19358 , n19014 , n19357 );
and ( n19359 , n18102 , n18440 );
and ( n19360 , n18441 , n18444 );
or ( n19361 , n19359 , n19360 );
xor ( n19362 , n19358 , n19361 );
buf ( n19363 , n19362 );
buf ( n19364 , n19363 );
not ( n19365 , n19364 );
buf ( n19366 , n548 );
not ( n19367 , n19366 );
nor ( n19368 , n19365 , n19367 );
xor ( n19369 , n18732 , n19368 );
xor ( n19370 , n18456 , n18729 );
nor ( n19371 , n18448 , n19367 );
and ( n19372 , n19370 , n19371 );
xor ( n19373 , n19370 , n19371 );
xor ( n19374 , n18460 , n18727 );
nor ( n19375 , n17548 , n19367 );
and ( n19376 , n19374 , n19375 );
xor ( n19377 , n19374 , n19375 );
xor ( n19378 , n18464 , n18725 );
nor ( n19379 , n16669 , n19367 );
and ( n19380 , n19378 , n19379 );
xor ( n19381 , n19378 , n19379 );
xor ( n19382 , n18468 , n18723 );
nor ( n19383 , n15809 , n19367 );
and ( n19384 , n19382 , n19383 );
xor ( n19385 , n19382 , n19383 );
xor ( n19386 , n18472 , n18721 );
nor ( n19387 , n14968 , n19367 );
and ( n19388 , n19386 , n19387 );
xor ( n19389 , n19386 , n19387 );
xor ( n19390 , n18476 , n18719 );
nor ( n19391 , n14147 , n19367 );
and ( n19392 , n19390 , n19391 );
xor ( n19393 , n19390 , n19391 );
xor ( n19394 , n18480 , n18717 );
nor ( n19395 , n13349 , n19367 );
and ( n19396 , n19394 , n19395 );
xor ( n19397 , n19394 , n19395 );
xor ( n19398 , n18484 , n18715 );
nor ( n19399 , n12564 , n19367 );
and ( n19400 , n19398 , n19399 );
xor ( n19401 , n19398 , n19399 );
xor ( n19402 , n18488 , n18713 );
nor ( n19403 , n11799 , n19367 );
and ( n19404 , n19402 , n19403 );
xor ( n19405 , n19402 , n19403 );
xor ( n19406 , n18492 , n18711 );
nor ( n19407 , n11050 , n19367 );
and ( n19408 , n19406 , n19407 );
xor ( n19409 , n19406 , n19407 );
xor ( n19410 , n18496 , n18709 );
nor ( n19411 , n10321 , n19367 );
and ( n19412 , n19410 , n19411 );
xor ( n19413 , n19410 , n19411 );
xor ( n19414 , n18500 , n18707 );
nor ( n19415 , n9429 , n19367 );
and ( n19416 , n19414 , n19415 );
xor ( n19417 , n19414 , n19415 );
xor ( n19418 , n18504 , n18705 );
nor ( n19419 , n8949 , n19367 );
and ( n19420 , n19418 , n19419 );
xor ( n19421 , n19418 , n19419 );
xor ( n19422 , n18508 , n18703 );
nor ( n19423 , n9437 , n19367 );
and ( n19424 , n19422 , n19423 );
xor ( n19425 , n19422 , n19423 );
xor ( n19426 , n18512 , n18701 );
nor ( n19427 , n9446 , n19367 );
and ( n19428 , n19426 , n19427 );
xor ( n19429 , n19426 , n19427 );
xor ( n19430 , n18516 , n18699 );
nor ( n19431 , n9455 , n19367 );
and ( n19432 , n19430 , n19431 );
xor ( n19433 , n19430 , n19431 );
xor ( n19434 , n18520 , n18697 );
nor ( n19435 , n9464 , n19367 );
and ( n19436 , n19434 , n19435 );
xor ( n19437 , n19434 , n19435 );
xor ( n19438 , n18524 , n18695 );
nor ( n19439 , n9473 , n19367 );
and ( n19440 , n19438 , n19439 );
xor ( n19441 , n19438 , n19439 );
xor ( n19442 , n18528 , n18693 );
nor ( n19443 , n9482 , n19367 );
and ( n19444 , n19442 , n19443 );
xor ( n19445 , n19442 , n19443 );
xor ( n19446 , n18532 , n18691 );
nor ( n19447 , n9491 , n19367 );
and ( n19448 , n19446 , n19447 );
xor ( n19449 , n19446 , n19447 );
xor ( n19450 , n18536 , n18689 );
nor ( n19451 , n9500 , n19367 );
and ( n19452 , n19450 , n19451 );
xor ( n19453 , n19450 , n19451 );
xor ( n19454 , n18540 , n18687 );
nor ( n19455 , n9509 , n19367 );
and ( n19456 , n19454 , n19455 );
xor ( n19457 , n19454 , n19455 );
xor ( n19458 , n18544 , n18685 );
nor ( n19459 , n9518 , n19367 );
and ( n19460 , n19458 , n19459 );
xor ( n19461 , n19458 , n19459 );
xor ( n19462 , n18548 , n18683 );
nor ( n19463 , n9527 , n19367 );
and ( n19464 , n19462 , n19463 );
xor ( n19465 , n19462 , n19463 );
xor ( n19466 , n18552 , n18681 );
nor ( n19467 , n9536 , n19367 );
and ( n19468 , n19466 , n19467 );
xor ( n19469 , n19466 , n19467 );
xor ( n19470 , n18556 , n18679 );
nor ( n19471 , n9545 , n19367 );
and ( n19472 , n19470 , n19471 );
xor ( n19473 , n19470 , n19471 );
xor ( n19474 , n18560 , n18677 );
nor ( n19475 , n9554 , n19367 );
and ( n19476 , n19474 , n19475 );
xor ( n19477 , n19474 , n19475 );
xor ( n19478 , n18564 , n18675 );
nor ( n19479 , n9563 , n19367 );
and ( n19480 , n19478 , n19479 );
xor ( n19481 , n19478 , n19479 );
xor ( n19482 , n18568 , n18673 );
nor ( n19483 , n9572 , n19367 );
and ( n19484 , n19482 , n19483 );
xor ( n19485 , n19482 , n19483 );
xor ( n19486 , n18572 , n18671 );
nor ( n19487 , n9581 , n19367 );
and ( n19488 , n19486 , n19487 );
xor ( n19489 , n19486 , n19487 );
xor ( n19490 , n18576 , n18669 );
nor ( n19491 , n9590 , n19367 );
and ( n19492 , n19490 , n19491 );
xor ( n19493 , n19490 , n19491 );
xor ( n19494 , n18580 , n18667 );
nor ( n19495 , n9599 , n19367 );
and ( n19496 , n19494 , n19495 );
xor ( n19497 , n19494 , n19495 );
xor ( n19498 , n18584 , n18665 );
nor ( n19499 , n9608 , n19367 );
and ( n19500 , n19498 , n19499 );
xor ( n19501 , n19498 , n19499 );
xor ( n19502 , n18588 , n18663 );
nor ( n19503 , n9617 , n19367 );
and ( n19504 , n19502 , n19503 );
xor ( n19505 , n19502 , n19503 );
xor ( n19506 , n18592 , n18661 );
nor ( n19507 , n9626 , n19367 );
and ( n19508 , n19506 , n19507 );
xor ( n19509 , n19506 , n19507 );
xor ( n19510 , n18596 , n18659 );
nor ( n19511 , n9635 , n19367 );
and ( n19512 , n19510 , n19511 );
xor ( n19513 , n19510 , n19511 );
xor ( n19514 , n18600 , n18657 );
nor ( n19515 , n9644 , n19367 );
and ( n19516 , n19514 , n19515 );
xor ( n19517 , n19514 , n19515 );
xor ( n19518 , n18604 , n18655 );
nor ( n19519 , n9653 , n19367 );
and ( n19520 , n19518 , n19519 );
xor ( n19521 , n19518 , n19519 );
xor ( n19522 , n18608 , n18653 );
nor ( n19523 , n9662 , n19367 );
and ( n19524 , n19522 , n19523 );
xor ( n19525 , n19522 , n19523 );
xor ( n19526 , n18612 , n18651 );
nor ( n19527 , n9671 , n19367 );
and ( n19528 , n19526 , n19527 );
xor ( n19529 , n19526 , n19527 );
xor ( n19530 , n18616 , n18649 );
nor ( n19531 , n9680 , n19367 );
and ( n19532 , n19530 , n19531 );
xor ( n19533 , n19530 , n19531 );
xor ( n19534 , n18620 , n18647 );
nor ( n19535 , n9689 , n19367 );
and ( n19536 , n19534 , n19535 );
xor ( n19537 , n19534 , n19535 );
xor ( n19538 , n18624 , n18645 );
nor ( n19539 , n9698 , n19367 );
and ( n19540 , n19538 , n19539 );
xor ( n19541 , n19538 , n19539 );
xor ( n19542 , n18628 , n18643 );
nor ( n19543 , n9707 , n19367 );
and ( n19544 , n19542 , n19543 );
xor ( n19545 , n19542 , n19543 );
xor ( n19546 , n18632 , n18641 );
nor ( n19547 , n9716 , n19367 );
and ( n19548 , n19546 , n19547 );
xor ( n19549 , n19546 , n19547 );
xor ( n19550 , n18636 , n18639 );
nor ( n19551 , n9725 , n19367 );
and ( n19552 , n19550 , n19551 );
xor ( n19553 , n19550 , n19551 );
xor ( n19554 , n18637 , n18638 );
nor ( n19555 , n9734 , n19367 );
and ( n19556 , n19554 , n19555 );
xor ( n19557 , n19554 , n19555 );
nor ( n19558 , n9752 , n18450 );
nor ( n19559 , n9743 , n19367 );
and ( n19560 , n19558 , n19559 );
and ( n19561 , n19557 , n19560 );
or ( n19562 , n19556 , n19561 );
and ( n19563 , n19553 , n19562 );
or ( n19564 , n19552 , n19563 );
and ( n19565 , n19549 , n19564 );
or ( n19566 , n19548 , n19565 );
and ( n19567 , n19545 , n19566 );
or ( n19568 , n19544 , n19567 );
and ( n19569 , n19541 , n19568 );
or ( n19570 , n19540 , n19569 );
and ( n19571 , n19537 , n19570 );
or ( n19572 , n19536 , n19571 );
and ( n19573 , n19533 , n19572 );
or ( n19574 , n19532 , n19573 );
and ( n19575 , n19529 , n19574 );
or ( n19576 , n19528 , n19575 );
and ( n19577 , n19525 , n19576 );
or ( n19578 , n19524 , n19577 );
and ( n19579 , n19521 , n19578 );
or ( n19580 , n19520 , n19579 );
and ( n19581 , n19517 , n19580 );
or ( n19582 , n19516 , n19581 );
and ( n19583 , n19513 , n19582 );
or ( n19584 , n19512 , n19583 );
and ( n19585 , n19509 , n19584 );
or ( n19586 , n19508 , n19585 );
and ( n19587 , n19505 , n19586 );
or ( n19588 , n19504 , n19587 );
and ( n19589 , n19501 , n19588 );
or ( n19590 , n19500 , n19589 );
and ( n19591 , n19497 , n19590 );
or ( n19592 , n19496 , n19591 );
and ( n19593 , n19493 , n19592 );
or ( n19594 , n19492 , n19593 );
and ( n19595 , n19489 , n19594 );
or ( n19596 , n19488 , n19595 );
and ( n19597 , n19485 , n19596 );
or ( n19598 , n19484 , n19597 );
and ( n19599 , n19481 , n19598 );
or ( n19600 , n19480 , n19599 );
and ( n19601 , n19477 , n19600 );
or ( n19602 , n19476 , n19601 );
and ( n19603 , n19473 , n19602 );
or ( n19604 , n19472 , n19603 );
and ( n19605 , n19469 , n19604 );
or ( n19606 , n19468 , n19605 );
and ( n19607 , n19465 , n19606 );
or ( n19608 , n19464 , n19607 );
and ( n19609 , n19461 , n19608 );
or ( n19610 , n19460 , n19609 );
and ( n19611 , n19457 , n19610 );
or ( n19612 , n19456 , n19611 );
and ( n19613 , n19453 , n19612 );
or ( n19614 , n19452 , n19613 );
and ( n19615 , n19449 , n19614 );
or ( n19616 , n19448 , n19615 );
and ( n19617 , n19445 , n19616 );
or ( n19618 , n19444 , n19617 );
and ( n19619 , n19441 , n19618 );
or ( n19620 , n19440 , n19619 );
and ( n19621 , n19437 , n19620 );
or ( n19622 , n19436 , n19621 );
and ( n19623 , n19433 , n19622 );
or ( n19624 , n19432 , n19623 );
and ( n19625 , n19429 , n19624 );
or ( n19626 , n19428 , n19625 );
and ( n19627 , n19425 , n19626 );
or ( n19628 , n19424 , n19627 );
and ( n19629 , n19421 , n19628 );
or ( n19630 , n19420 , n19629 );
and ( n19631 , n19417 , n19630 );
or ( n19632 , n19416 , n19631 );
and ( n19633 , n19413 , n19632 );
or ( n19634 , n19412 , n19633 );
and ( n19635 , n19409 , n19634 );
or ( n19636 , n19408 , n19635 );
and ( n19637 , n19405 , n19636 );
or ( n19638 , n19404 , n19637 );
and ( n19639 , n19401 , n19638 );
or ( n19640 , n19400 , n19639 );
and ( n19641 , n19397 , n19640 );
or ( n19642 , n19396 , n19641 );
and ( n19643 , n19393 , n19642 );
or ( n19644 , n19392 , n19643 );
and ( n19645 , n19389 , n19644 );
or ( n19646 , n19388 , n19645 );
and ( n19647 , n19385 , n19646 );
or ( n19648 , n19384 , n19647 );
and ( n19649 , n19381 , n19648 );
or ( n19650 , n19380 , n19649 );
and ( n19651 , n19377 , n19650 );
or ( n19652 , n19376 , n19651 );
and ( n19653 , n19373 , n19652 );
or ( n19654 , n19372 , n19653 );
xor ( n19655 , n19369 , n19654 );
buf ( n19656 , n484 );
not ( n19657 , n19656 );
nor ( n19658 , n601 , n19657 );
buf ( n19659 , n19658 );
nor ( n19660 , n622 , n17828 );
xor ( n19661 , n19659 , n19660 );
buf ( n19662 , n19661 );
nor ( n19663 , n646 , n16943 );
xor ( n19664 , n19662 , n19663 );
and ( n19665 , n18736 , n18737 );
buf ( n19666 , n19665 );
xor ( n19667 , n19664 , n19666 );
nor ( n19668 , n684 , n16077 );
xor ( n19669 , n19667 , n19668 );
and ( n19670 , n18739 , n18740 );
and ( n19671 , n18741 , n18743 );
or ( n19672 , n19670 , n19671 );
xor ( n19673 , n19669 , n19672 );
nor ( n19674 , n733 , n15230 );
xor ( n19675 , n19673 , n19674 );
and ( n19676 , n18744 , n18745 );
and ( n19677 , n18746 , n18749 );
or ( n19678 , n19676 , n19677 );
xor ( n19679 , n19675 , n19678 );
nor ( n19680 , n796 , n14403 );
xor ( n19681 , n19679 , n19680 );
and ( n19682 , n18750 , n18751 );
and ( n19683 , n18752 , n18755 );
or ( n19684 , n19682 , n19683 );
xor ( n19685 , n19681 , n19684 );
nor ( n19686 , n868 , n13599 );
xor ( n19687 , n19685 , n19686 );
and ( n19688 , n18756 , n18757 );
and ( n19689 , n18758 , n18761 );
or ( n19690 , n19688 , n19689 );
xor ( n19691 , n19687 , n19690 );
nor ( n19692 , n958 , n12808 );
xor ( n19693 , n19691 , n19692 );
and ( n19694 , n18762 , n18763 );
and ( n19695 , n18764 , n18767 );
or ( n19696 , n19694 , n19695 );
xor ( n19697 , n19693 , n19696 );
nor ( n19698 , n1062 , n12037 );
xor ( n19699 , n19697 , n19698 );
and ( n19700 , n18768 , n18769 );
and ( n19701 , n18770 , n18773 );
or ( n19702 , n19700 , n19701 );
xor ( n19703 , n19699 , n19702 );
nor ( n19704 , n1176 , n11282 );
xor ( n19705 , n19703 , n19704 );
and ( n19706 , n18774 , n18775 );
and ( n19707 , n18776 , n18779 );
or ( n19708 , n19706 , n19707 );
xor ( n19709 , n19705 , n19708 );
nor ( n19710 , n1303 , n10547 );
xor ( n19711 , n19709 , n19710 );
and ( n19712 , n18780 , n18781 );
and ( n19713 , n18782 , n18785 );
or ( n19714 , n19712 , n19713 );
xor ( n19715 , n19711 , n19714 );
nor ( n19716 , n1445 , n9829 );
xor ( n19717 , n19715 , n19716 );
and ( n19718 , n18786 , n18787 );
and ( n19719 , n18788 , n18791 );
or ( n19720 , n19718 , n19719 );
xor ( n19721 , n19717 , n19720 );
nor ( n19722 , n1598 , n8955 );
xor ( n19723 , n19721 , n19722 );
and ( n19724 , n18792 , n18793 );
and ( n19725 , n18794 , n18797 );
or ( n19726 , n19724 , n19725 );
xor ( n19727 , n19723 , n19726 );
nor ( n19728 , n1766 , n603 );
xor ( n19729 , n19727 , n19728 );
and ( n19730 , n18798 , n18799 );
and ( n19731 , n18800 , n18803 );
or ( n19732 , n19730 , n19731 );
xor ( n19733 , n19729 , n19732 );
nor ( n19734 , n1945 , n652 );
xor ( n19735 , n19733 , n19734 );
and ( n19736 , n18804 , n18805 );
and ( n19737 , n18806 , n18809 );
or ( n19738 , n19736 , n19737 );
xor ( n19739 , n19735 , n19738 );
nor ( n19740 , n2137 , n624 );
xor ( n19741 , n19739 , n19740 );
and ( n19742 , n18810 , n18811 );
and ( n19743 , n18812 , n18815 );
or ( n19744 , n19742 , n19743 );
xor ( n19745 , n19741 , n19744 );
nor ( n19746 , n2343 , n648 );
xor ( n19747 , n19745 , n19746 );
and ( n19748 , n18816 , n18817 );
and ( n19749 , n18818 , n18821 );
or ( n19750 , n19748 , n19749 );
xor ( n19751 , n19747 , n19750 );
nor ( n19752 , n2566 , n686 );
xor ( n19753 , n19751 , n19752 );
and ( n19754 , n18822 , n18823 );
and ( n19755 , n18824 , n18827 );
or ( n19756 , n19754 , n19755 );
xor ( n19757 , n19753 , n19756 );
nor ( n19758 , n2797 , n735 );
xor ( n19759 , n19757 , n19758 );
and ( n19760 , n18828 , n18829 );
and ( n19761 , n18830 , n18833 );
or ( n19762 , n19760 , n19761 );
xor ( n19763 , n19759 , n19762 );
nor ( n19764 , n3043 , n798 );
xor ( n19765 , n19763 , n19764 );
and ( n19766 , n18834 , n18835 );
and ( n19767 , n18836 , n18839 );
or ( n19768 , n19766 , n19767 );
xor ( n19769 , n19765 , n19768 );
nor ( n19770 , n3300 , n870 );
xor ( n19771 , n19769 , n19770 );
and ( n19772 , n18840 , n18841 );
and ( n19773 , n18842 , n18845 );
or ( n19774 , n19772 , n19773 );
xor ( n19775 , n19771 , n19774 );
nor ( n19776 , n3570 , n960 );
xor ( n19777 , n19775 , n19776 );
and ( n19778 , n18846 , n18847 );
and ( n19779 , n18848 , n18851 );
or ( n19780 , n19778 , n19779 );
xor ( n19781 , n19777 , n19780 );
nor ( n19782 , n3853 , n1064 );
xor ( n19783 , n19781 , n19782 );
and ( n19784 , n18852 , n18853 );
and ( n19785 , n18854 , n18857 );
or ( n19786 , n19784 , n19785 );
xor ( n19787 , n19783 , n19786 );
nor ( n19788 , n4151 , n1178 );
xor ( n19789 , n19787 , n19788 );
and ( n19790 , n18858 , n18859 );
and ( n19791 , n18860 , n18863 );
or ( n19792 , n19790 , n19791 );
xor ( n19793 , n19789 , n19792 );
nor ( n19794 , n4458 , n1305 );
xor ( n19795 , n19793 , n19794 );
and ( n19796 , n18864 , n18865 );
and ( n19797 , n18866 , n18869 );
or ( n19798 , n19796 , n19797 );
xor ( n19799 , n19795 , n19798 );
nor ( n19800 , n4786 , n1447 );
xor ( n19801 , n19799 , n19800 );
and ( n19802 , n18870 , n18871 );
and ( n19803 , n18872 , n18875 );
or ( n19804 , n19802 , n19803 );
xor ( n19805 , n19801 , n19804 );
nor ( n19806 , n5126 , n1600 );
xor ( n19807 , n19805 , n19806 );
and ( n19808 , n18876 , n18877 );
and ( n19809 , n18878 , n18881 );
or ( n19810 , n19808 , n19809 );
xor ( n19811 , n19807 , n19810 );
nor ( n19812 , n5477 , n1768 );
xor ( n19813 , n19811 , n19812 );
and ( n19814 , n18882 , n18883 );
and ( n19815 , n18884 , n18887 );
or ( n19816 , n19814 , n19815 );
xor ( n19817 , n19813 , n19816 );
nor ( n19818 , n5838 , n1947 );
xor ( n19819 , n19817 , n19818 );
and ( n19820 , n18888 , n18889 );
and ( n19821 , n18890 , n18893 );
or ( n19822 , n19820 , n19821 );
xor ( n19823 , n19819 , n19822 );
nor ( n19824 , n6212 , n2139 );
xor ( n19825 , n19823 , n19824 );
and ( n19826 , n18894 , n18895 );
and ( n19827 , n18896 , n18899 );
or ( n19828 , n19826 , n19827 );
xor ( n19829 , n19825 , n19828 );
nor ( n19830 , n6596 , n2345 );
xor ( n19831 , n19829 , n19830 );
and ( n19832 , n18900 , n18901 );
and ( n19833 , n18902 , n18905 );
or ( n19834 , n19832 , n19833 );
xor ( n19835 , n19831 , n19834 );
nor ( n19836 , n6997 , n2568 );
xor ( n19837 , n19835 , n19836 );
and ( n19838 , n18906 , n18907 );
and ( n19839 , n18908 , n18911 );
or ( n19840 , n19838 , n19839 );
xor ( n19841 , n19837 , n19840 );
nor ( n19842 , n7413 , n2799 );
xor ( n19843 , n19841 , n19842 );
and ( n19844 , n18912 , n18913 );
and ( n19845 , n18914 , n18917 );
or ( n19846 , n19844 , n19845 );
xor ( n19847 , n19843 , n19846 );
nor ( n19848 , n7841 , n3045 );
xor ( n19849 , n19847 , n19848 );
and ( n19850 , n18918 , n18919 );
and ( n19851 , n18920 , n18923 );
or ( n19852 , n19850 , n19851 );
xor ( n19853 , n19849 , n19852 );
nor ( n19854 , n8281 , n3302 );
xor ( n19855 , n19853 , n19854 );
and ( n19856 , n18924 , n18925 );
and ( n19857 , n18926 , n18929 );
or ( n19858 , n19856 , n19857 );
xor ( n19859 , n19855 , n19858 );
nor ( n19860 , n8737 , n3572 );
xor ( n19861 , n19859 , n19860 );
and ( n19862 , n18930 , n18931 );
and ( n19863 , n18932 , n18935 );
or ( n19864 , n19862 , n19863 );
xor ( n19865 , n19861 , n19864 );
nor ( n19866 , n9420 , n3855 );
xor ( n19867 , n19865 , n19866 );
and ( n19868 , n18936 , n18937 );
and ( n19869 , n18938 , n18941 );
or ( n19870 , n19868 , n19869 );
xor ( n19871 , n19867 , n19870 );
nor ( n19872 , n10312 , n4153 );
xor ( n19873 , n19871 , n19872 );
and ( n19874 , n18942 , n18943 );
and ( n19875 , n18944 , n18947 );
or ( n19876 , n19874 , n19875 );
xor ( n19877 , n19873 , n19876 );
nor ( n19878 , n11041 , n4460 );
xor ( n19879 , n19877 , n19878 );
and ( n19880 , n18948 , n18949 );
and ( n19881 , n18950 , n18953 );
or ( n19882 , n19880 , n19881 );
xor ( n19883 , n19879 , n19882 );
nor ( n19884 , n11790 , n4788 );
xor ( n19885 , n19883 , n19884 );
and ( n19886 , n18954 , n18955 );
and ( n19887 , n18956 , n18959 );
or ( n19888 , n19886 , n19887 );
xor ( n19889 , n19885 , n19888 );
nor ( n19890 , n12555 , n5128 );
xor ( n19891 , n19889 , n19890 );
and ( n19892 , n18960 , n18961 );
and ( n19893 , n18962 , n18965 );
or ( n19894 , n19892 , n19893 );
xor ( n19895 , n19891 , n19894 );
nor ( n19896 , n13340 , n5479 );
xor ( n19897 , n19895 , n19896 );
and ( n19898 , n18966 , n18967 );
and ( n19899 , n18968 , n18971 );
or ( n19900 , n19898 , n19899 );
xor ( n19901 , n19897 , n19900 );
nor ( n19902 , n14138 , n5840 );
xor ( n19903 , n19901 , n19902 );
and ( n19904 , n18972 , n18973 );
and ( n19905 , n18974 , n18977 );
or ( n19906 , n19904 , n19905 );
xor ( n19907 , n19903 , n19906 );
nor ( n19908 , n14959 , n6214 );
xor ( n19909 , n19907 , n19908 );
and ( n19910 , n18978 , n18979 );
and ( n19911 , n18980 , n18983 );
or ( n19912 , n19910 , n19911 );
xor ( n19913 , n19909 , n19912 );
nor ( n19914 , n15800 , n6598 );
xor ( n19915 , n19913 , n19914 );
and ( n19916 , n18984 , n18985 );
and ( n19917 , n18986 , n18989 );
or ( n19918 , n19916 , n19917 );
xor ( n19919 , n19915 , n19918 );
nor ( n19920 , n16660 , n6999 );
xor ( n19921 , n19919 , n19920 );
and ( n19922 , n18990 , n18991 );
and ( n19923 , n18992 , n18995 );
or ( n19924 , n19922 , n19923 );
xor ( n19925 , n19921 , n19924 );
nor ( n19926 , n17539 , n7415 );
xor ( n19927 , n19925 , n19926 );
and ( n19928 , n18996 , n18997 );
and ( n19929 , n18998 , n19001 );
or ( n19930 , n19928 , n19929 );
xor ( n19931 , n19927 , n19930 );
nor ( n19932 , n18439 , n7843 );
xor ( n19933 , n19931 , n19932 );
and ( n19934 , n19002 , n19003 );
and ( n19935 , n19004 , n19007 );
or ( n19936 , n19934 , n19935 );
xor ( n19937 , n19933 , n19936 );
nor ( n19938 , n19356 , n8283 );
xor ( n19939 , n19937 , n19938 );
and ( n19940 , n19008 , n19009 );
and ( n19941 , n19010 , n19013 );
or ( n19942 , n19940 , n19941 );
xor ( n19943 , n19939 , n19942 );
and ( n19944 , n19337 , n19341 );
and ( n19945 , n19024 , n19332 );
and ( n19946 , n19332 , n19342 );
and ( n19947 , n19024 , n19342 );
or ( n19948 , n19945 , n19946 , n19947 );
xor ( n19949 , n19944 , n19948 );
and ( n19950 , n19028 , n19232 );
and ( n19951 , n19232 , n19331 );
and ( n19952 , n19028 , n19331 );
or ( n19953 , n19950 , n19951 , n19952 );
and ( n19954 , n19032 , n19107 );
and ( n19955 , n19107 , n19231 );
and ( n19956 , n19032 , n19231 );
or ( n19957 , n19954 , n19955 , n19956 );
and ( n19958 , n19112 , n19159 );
and ( n19959 , n19159 , n19230 );
and ( n19960 , n19112 , n19230 );
or ( n19961 , n19958 , n19959 , n19960 );
and ( n19962 , n19045 , n19082 );
and ( n19963 , n19082 , n19105 );
and ( n19964 , n19045 , n19105 );
or ( n19965 , n19962 , n19963 , n19964 );
and ( n19966 , n19116 , n19120 );
and ( n19967 , n19120 , n19158 );
and ( n19968 , n19116 , n19158 );
or ( n19969 , n19966 , n19967 , n19968 );
xor ( n19970 , n19965 , n19969 );
and ( n19971 , n19087 , n19091 );
and ( n19972 , n19091 , n19104 );
and ( n19973 , n19087 , n19104 );
or ( n19974 , n19971 , n19972 , n19973 );
and ( n19975 , n19069 , n19074 );
and ( n19976 , n19074 , n19080 );
and ( n19977 , n19069 , n19080 );
or ( n19978 , n19975 , n19976 , n19977 );
and ( n19979 , n19059 , n19060 );
and ( n19980 , n19060 , n19062 );
and ( n19981 , n19059 , n19062 );
or ( n19982 , n19979 , n19980 , n19981 );
and ( n19983 , n19070 , n19071 );
and ( n19984 , n19071 , n19073 );
and ( n19985 , n19070 , n19073 );
or ( n19986 , n19983 , n19984 , n19985 );
xor ( n19987 , n19982 , n19986 );
and ( n19988 , n7385 , n2298 );
and ( n19989 , n7808 , n2100 );
xor ( n19990 , n19988 , n19989 );
and ( n19991 , n8079 , n1882 );
xor ( n19992 , n19990 , n19991 );
xor ( n19993 , n19987 , n19992 );
xor ( n19994 , n19978 , n19993 );
and ( n19995 , n19076 , n19077 );
and ( n19996 , n19077 , n19079 );
and ( n19997 , n19076 , n19079 );
or ( n19998 , n19995 , n19996 , n19997 );
and ( n19999 , n6187 , n2981 );
and ( n20000 , n6569 , n2739 );
xor ( n20001 , n19999 , n20000 );
and ( n20002 , n6816 , n2544 );
xor ( n20003 , n20001 , n20002 );
xor ( n20004 , n19998 , n20003 );
and ( n20005 , n4959 , n3749 );
and ( n20006 , n5459 , n3495 );
xor ( n20007 , n20005 , n20006 );
and ( n20008 , n5819 , n3271 );
xor ( n20009 , n20007 , n20008 );
xor ( n20010 , n20004 , n20009 );
xor ( n20011 , n19994 , n20010 );
xor ( n20012 , n19974 , n20011 );
and ( n20013 , n19096 , n19100 );
and ( n20014 , n19100 , n19103 );
and ( n20015 , n19096 , n19103 );
or ( n20016 , n20013 , n20014 , n20015 );
and ( n20017 , n19129 , n19134 );
and ( n20018 , n19134 , n19140 );
and ( n20019 , n19129 , n19140 );
or ( n20020 , n20017 , n20018 , n20019 );
xor ( n20021 , n20016 , n20020 );
and ( n20022 , n4132 , n4403 );
and ( n20023 , n4438 , n4102 );
and ( n20024 , n20022 , n20023 );
and ( n20025 , n20023 , n19102 );
and ( n20026 , n20022 , n19102 );
or ( n20027 , n20024 , n20025 , n20026 );
and ( n20028 , n19130 , n19131 );
and ( n20029 , n19131 , n19133 );
and ( n20030 , n19130 , n19133 );
or ( n20031 , n20028 , n20029 , n20030 );
xor ( n20032 , n20027 , n20031 );
and ( n20033 , n4132 , n4730 );
buf ( n20034 , n4438 );
xor ( n20035 , n20033 , n20034 );
and ( n20036 , n4766 , n4102 );
xor ( n20037 , n20035 , n20036 );
xor ( n20038 , n20032 , n20037 );
xor ( n20039 , n20021 , n20038 );
xor ( n20040 , n20012 , n20039 );
xor ( n20041 , n19970 , n20040 );
xor ( n20042 , n19961 , n20041 );
and ( n20043 , n19164 , n19190 );
and ( n20044 , n19190 , n19229 );
and ( n20045 , n19164 , n19229 );
or ( n20046 , n20043 , n20044 , n20045 );
and ( n20047 , n19125 , n19141 );
and ( n20048 , n19141 , n19157 );
and ( n20049 , n19125 , n19157 );
or ( n20050 , n20047 , n20048 , n20049 );
and ( n20051 , n19168 , n19172 );
and ( n20052 , n19172 , n19189 );
and ( n20053 , n19168 , n19189 );
or ( n20054 , n20051 , n20052 , n20053 );
xor ( n20055 , n20050 , n20054 );
and ( n20056 , n19146 , n19150 );
and ( n20057 , n19150 , n19156 );
and ( n20058 , n19146 , n19156 );
or ( n20059 , n20056 , n20057 , n20058 );
and ( n20060 , n19136 , n19137 );
and ( n20061 , n19137 , n19139 );
and ( n20062 , n19136 , n19139 );
or ( n20063 , n20060 , n20061 , n20062 );
and ( n20064 , n3182 , n5765 );
and ( n20065 , n3545 , n5408 );
xor ( n20066 , n20064 , n20065 );
and ( n20067 , n3801 , n5103 );
xor ( n20068 , n20066 , n20067 );
xor ( n20069 , n20063 , n20068 );
and ( n20070 , n2462 , n6971 );
and ( n20071 , n2779 , n6504 );
xor ( n20072 , n20070 , n20071 );
and ( n20073 , n3024 , n6132 );
xor ( n20074 , n20072 , n20073 );
xor ( n20075 , n20069 , n20074 );
xor ( n20076 , n20059 , n20075 );
and ( n20077 , n19152 , n19153 );
and ( n20078 , n19153 , n19155 );
and ( n20079 , n19152 , n19155 );
or ( n20080 , n20077 , n20078 , n20079 );
and ( n20081 , n19178 , n19179 );
and ( n20082 , n19179 , n19181 );
and ( n20083 , n19178 , n19181 );
or ( n20084 , n20081 , n20082 , n20083 );
xor ( n20085 , n20080 , n20084 );
and ( n20086 , n1933 , n8243 );
and ( n20087 , n2120 , n7662 );
xor ( n20088 , n20086 , n20087 );
and ( n20089 , n2324 , n7310 );
xor ( n20090 , n20088 , n20089 );
xor ( n20091 , n20085 , n20090 );
xor ( n20092 , n20076 , n20091 );
xor ( n20093 , n20055 , n20092 );
xor ( n20094 , n20046 , n20093 );
and ( n20095 , n19195 , n19210 );
and ( n20096 , n19210 , n19228 );
and ( n20097 , n19195 , n19228 );
or ( n20098 , n20095 , n20096 , n20097 );
and ( n20099 , n19177 , n19182 );
and ( n20100 , n19182 , n19188 );
and ( n20101 , n19177 , n19188 );
or ( n20102 , n20099 , n20100 , n20101 );
and ( n20103 , n19199 , n19203 );
and ( n20104 , n19203 , n19209 );
and ( n20105 , n19199 , n19209 );
or ( n20106 , n20103 , n20104 , n20105 );
xor ( n20107 , n20102 , n20106 );
and ( n20108 , n19184 , n19185 );
and ( n20109 , n19185 , n19187 );
and ( n20110 , n19184 , n19187 );
or ( n20111 , n20108 , n20109 , n20110 );
and ( n20112 , n1383 , n10239 );
and ( n20113 , n1580 , n9348 );
xor ( n20114 , n20112 , n20113 );
and ( n20115 , n1694 , n8669 );
xor ( n20116 , n20114 , n20115 );
xor ( n20117 , n20111 , n20116 );
and ( n20118 , n1047 , n12531 );
and ( n20119 , n1164 , n11718 );
xor ( n20120 , n20118 , n20119 );
and ( n20121 , n1287 , n10977 );
xor ( n20122 , n20120 , n20121 );
xor ( n20123 , n20117 , n20122 );
xor ( n20124 , n20107 , n20123 );
xor ( n20125 , n20098 , n20124 );
and ( n20126 , n19215 , n19220 );
and ( n20127 , n19220 , n19227 );
and ( n20128 , n19215 , n19227 );
or ( n20129 , n20126 , n20127 , n20128 );
and ( n20130 , n19205 , n19206 );
and ( n20131 , n19206 , n19208 );
and ( n20132 , n19205 , n19208 );
or ( n20133 , n20130 , n20131 , n20132 );
and ( n20134 , n19216 , n19217 );
and ( n20135 , n19217 , n19219 );
and ( n20136 , n19216 , n19219 );
or ( n20137 , n20134 , n20135 , n20136 );
xor ( n20138 , n20133 , n20137 );
and ( n20139 , n783 , n14838 );
and ( n20140 , n856 , n14044 );
xor ( n20141 , n20139 , n20140 );
and ( n20142 , n925 , n13256 );
xor ( n20143 , n20141 , n20142 );
xor ( n20144 , n20138 , n20143 );
xor ( n20145 , n20129 , n20144 );
and ( n20146 , n19223 , n19224 );
and ( n20147 , n19224 , n19226 );
and ( n20148 , n19223 , n19226 );
or ( n20149 , n20146 , n20147 , n20148 );
and ( n20150 , n632 , n17422 );
and ( n20151 , n671 , n16550 );
xor ( n20152 , n20150 , n20151 );
and ( n20153 , n715 , n15691 );
xor ( n20154 , n20152 , n20153 );
xor ( n20155 , n20149 , n20154 );
buf ( n20156 , n420 );
and ( n20157 , n599 , n20156 );
and ( n20158 , n608 , n19222 );
xor ( n20159 , n20157 , n20158 );
and ( n20160 , n611 , n18407 );
xor ( n20161 , n20159 , n20160 );
xor ( n20162 , n20155 , n20161 );
xor ( n20163 , n20145 , n20162 );
xor ( n20164 , n20125 , n20163 );
xor ( n20165 , n20094 , n20164 );
xor ( n20166 , n20042 , n20165 );
xor ( n20167 , n19957 , n20166 );
and ( n20168 , n19036 , n19040 );
and ( n20169 , n19040 , n19106 );
and ( n20170 , n19036 , n19106 );
or ( n20171 , n20168 , n20169 , n20170 );
and ( n20172 , n19246 , n19282 );
and ( n20173 , n19282 , n19329 );
and ( n20174 , n19246 , n19329 );
or ( n20175 , n20172 , n20173 , n20174 );
xor ( n20176 , n20171 , n20175 );
and ( n20177 , n19250 , n19254 );
and ( n20178 , n19254 , n19281 );
and ( n20179 , n19250 , n19281 );
or ( n20180 , n20177 , n20178 , n20179 );
and ( n20181 , n19259 , n19263 );
and ( n20182 , n19263 , n19280 );
and ( n20183 , n19259 , n19280 );
or ( n20184 , n20181 , n20182 , n20183 );
and ( n20185 , n19049 , n19064 );
and ( n20186 , n19064 , n19081 );
and ( n20187 , n19049 , n19081 );
or ( n20188 , n20185 , n20186 , n20187 );
xor ( n20189 , n20184 , n20188 );
and ( n20190 , n19268 , n19273 );
and ( n20191 , n19273 , n19279 );
and ( n20192 , n19268 , n19279 );
or ( n20193 , n20190 , n20191 , n20192 );
and ( n20194 , n19053 , n19057 );
and ( n20195 , n19057 , n19063 );
and ( n20196 , n19053 , n19063 );
or ( n20197 , n20194 , n20195 , n20196 );
xor ( n20198 , n20193 , n20197 );
and ( n20199 , n19275 , n19276 );
and ( n20200 , n19276 , n19278 );
and ( n20201 , n19275 , n19278 );
or ( n20202 , n20199 , n20200 , n20201 );
and ( n20203 , n11015 , n1254 );
and ( n20204 , n11769 , n1134 );
xor ( n20205 , n20203 , n20204 );
and ( n20206 , n12320 , n1034 );
xor ( n20207 , n20205 , n20206 );
xor ( n20208 , n20202 , n20207 );
and ( n20209 , n8718 , n1738 );
and ( n20210 , n9400 , n1551 );
xor ( n20211 , n20209 , n20210 );
and ( n20212 , n10291 , n1424 );
xor ( n20213 , n20211 , n20212 );
xor ( n20214 , n20208 , n20213 );
xor ( n20215 , n20198 , n20214 );
xor ( n20216 , n20189 , n20215 );
xor ( n20217 , n20180 , n20216 );
and ( n20218 , n19296 , n19311 );
and ( n20219 , n19311 , n19327 );
and ( n20220 , n19296 , n19327 );
or ( n20221 , n20218 , n20219 , n20220 );
and ( n20222 , n19300 , n19304 );
and ( n20223 , n19304 , n19310 );
and ( n20224 , n19300 , n19310 );
or ( n20225 , n20222 , n20223 , n20224 );
and ( n20226 , n19317 , n19318 );
and ( n20227 , n19318 , n19320 );
and ( n20228 , n19317 , n19320 );
or ( n20229 , n20226 , n20227 , n20228 );
and ( n20230 , n18144 , n606 );
and ( n20231 , n19324 , n615 );
xor ( n20232 , n20230 , n20231 );
buf ( n20233 , n420 );
and ( n20234 , n20233 , n612 );
xor ( n20235 , n20232 , n20234 );
xor ( n20236 , n20229 , n20235 );
and ( n20237 , n15758 , n719 );
and ( n20238 , n16637 , n663 );
xor ( n20239 , n20237 , n20238 );
and ( n20240 , n17512 , n635 );
xor ( n20241 , n20239 , n20240 );
xor ( n20242 , n20236 , n20241 );
xor ( n20243 , n20225 , n20242 );
and ( n20244 , n19306 , n19307 );
and ( n20245 , n19307 , n19309 );
and ( n20246 , n19306 , n19309 );
or ( n20247 , n20244 , n20245 , n20246 );
and ( n20248 , n19269 , n19270 );
and ( n20249 , n19270 , n19272 );
and ( n20250 , n19269 , n19272 );
or ( n20251 , n20248 , n20249 , n20250 );
xor ( n20252 , n20247 , n20251 );
and ( n20253 , n13322 , n940 );
and ( n20254 , n14118 , n840 );
xor ( n20255 , n20253 , n20254 );
and ( n20256 , n14938 , n771 );
xor ( n20257 , n20255 , n20256 );
xor ( n20258 , n20252 , n20257 );
xor ( n20259 , n20243 , n20258 );
xor ( n20260 , n20221 , n20259 );
and ( n20261 , n19323 , n19325 );
and ( n20262 , n19316 , n19321 );
and ( n20263 , n19321 , n19326 );
and ( n20264 , n19316 , n19326 );
or ( n20265 , n20262 , n20263 , n20264 );
xor ( n20266 , n20261 , n20265 );
xor ( n20267 , n20260 , n20266 );
xor ( n20268 , n20217 , n20267 );
xor ( n20269 , n20176 , n20268 );
xor ( n20270 , n20167 , n20269 );
xor ( n20271 , n19953 , n20270 );
and ( n20272 , n19287 , n19291 );
and ( n20273 , n19291 , n19328 );
and ( n20274 , n19287 , n19328 );
or ( n20275 , n20272 , n20273 , n20274 );
and ( n20276 , n19237 , n19241 );
and ( n20277 , n19241 , n19330 );
and ( n20278 , n19237 , n19330 );
or ( n20279 , n20276 , n20277 , n20278 );
xor ( n20280 , n20275 , n20279 );
xor ( n20281 , n20271 , n20280 );
xor ( n20282 , n19949 , n20281 );
and ( n20283 , n19015 , n19019 );
and ( n20284 , n19019 , n19343 );
and ( n20285 , n19015 , n19343 );
or ( n20286 , n20283 , n20284 , n20285 );
xor ( n20287 , n20282 , n20286 );
and ( n20288 , n19344 , n19348 );
and ( n20289 , n19349 , n19352 );
or ( n20290 , n20288 , n20289 );
xor ( n20291 , n20287 , n20290 );
buf ( n20292 , n20291 );
buf ( n20293 , n20292 );
not ( n20294 , n20293 );
nor ( n20295 , n20294 , n8739 );
xor ( n20296 , n19943 , n20295 );
and ( n20297 , n19014 , n19357 );
and ( n20298 , n19358 , n19361 );
or ( n20299 , n20297 , n20298 );
xor ( n20300 , n20296 , n20299 );
buf ( n20301 , n20300 );
buf ( n20302 , n20301 );
not ( n20303 , n20302 );
buf ( n20304 , n549 );
not ( n20305 , n20304 );
nor ( n20306 , n20303 , n20305 );
xor ( n20307 , n19655 , n20306 );
xor ( n20308 , n19373 , n19652 );
nor ( n20309 , n19365 , n20305 );
and ( n20310 , n20308 , n20309 );
xor ( n20311 , n20308 , n20309 );
xor ( n20312 , n19377 , n19650 );
nor ( n20313 , n18448 , n20305 );
and ( n20314 , n20312 , n20313 );
xor ( n20315 , n20312 , n20313 );
xor ( n20316 , n19381 , n19648 );
nor ( n20317 , n17548 , n20305 );
and ( n20318 , n20316 , n20317 );
xor ( n20319 , n20316 , n20317 );
xor ( n20320 , n19385 , n19646 );
nor ( n20321 , n16669 , n20305 );
and ( n20322 , n20320 , n20321 );
xor ( n20323 , n20320 , n20321 );
xor ( n20324 , n19389 , n19644 );
nor ( n20325 , n15809 , n20305 );
and ( n20326 , n20324 , n20325 );
xor ( n20327 , n20324 , n20325 );
xor ( n20328 , n19393 , n19642 );
nor ( n20329 , n14968 , n20305 );
and ( n20330 , n20328 , n20329 );
xor ( n20331 , n20328 , n20329 );
xor ( n20332 , n19397 , n19640 );
nor ( n20333 , n14147 , n20305 );
and ( n20334 , n20332 , n20333 );
xor ( n20335 , n20332 , n20333 );
xor ( n20336 , n19401 , n19638 );
nor ( n20337 , n13349 , n20305 );
and ( n20338 , n20336 , n20337 );
xor ( n20339 , n20336 , n20337 );
xor ( n20340 , n19405 , n19636 );
nor ( n20341 , n12564 , n20305 );
and ( n20342 , n20340 , n20341 );
xor ( n20343 , n20340 , n20341 );
xor ( n20344 , n19409 , n19634 );
nor ( n20345 , n11799 , n20305 );
and ( n20346 , n20344 , n20345 );
xor ( n20347 , n20344 , n20345 );
xor ( n20348 , n19413 , n19632 );
nor ( n20349 , n11050 , n20305 );
and ( n20350 , n20348 , n20349 );
xor ( n20351 , n20348 , n20349 );
xor ( n20352 , n19417 , n19630 );
nor ( n20353 , n10321 , n20305 );
and ( n20354 , n20352 , n20353 );
xor ( n20355 , n20352 , n20353 );
xor ( n20356 , n19421 , n19628 );
nor ( n20357 , n9429 , n20305 );
and ( n20358 , n20356 , n20357 );
xor ( n20359 , n20356 , n20357 );
xor ( n20360 , n19425 , n19626 );
nor ( n20361 , n8949 , n20305 );
and ( n20362 , n20360 , n20361 );
xor ( n20363 , n20360 , n20361 );
xor ( n20364 , n19429 , n19624 );
nor ( n20365 , n9437 , n20305 );
and ( n20366 , n20364 , n20365 );
xor ( n20367 , n20364 , n20365 );
xor ( n20368 , n19433 , n19622 );
nor ( n20369 , n9446 , n20305 );
and ( n20370 , n20368 , n20369 );
xor ( n20371 , n20368 , n20369 );
xor ( n20372 , n19437 , n19620 );
nor ( n20373 , n9455 , n20305 );
and ( n20374 , n20372 , n20373 );
xor ( n20375 , n20372 , n20373 );
xor ( n20376 , n19441 , n19618 );
nor ( n20377 , n9464 , n20305 );
and ( n20378 , n20376 , n20377 );
xor ( n20379 , n20376 , n20377 );
xor ( n20380 , n19445 , n19616 );
nor ( n20381 , n9473 , n20305 );
and ( n20382 , n20380 , n20381 );
xor ( n20383 , n20380 , n20381 );
xor ( n20384 , n19449 , n19614 );
nor ( n20385 , n9482 , n20305 );
and ( n20386 , n20384 , n20385 );
xor ( n20387 , n20384 , n20385 );
xor ( n20388 , n19453 , n19612 );
nor ( n20389 , n9491 , n20305 );
and ( n20390 , n20388 , n20389 );
xor ( n20391 , n20388 , n20389 );
xor ( n20392 , n19457 , n19610 );
nor ( n20393 , n9500 , n20305 );
and ( n20394 , n20392 , n20393 );
xor ( n20395 , n20392 , n20393 );
xor ( n20396 , n19461 , n19608 );
nor ( n20397 , n9509 , n20305 );
and ( n20398 , n20396 , n20397 );
xor ( n20399 , n20396 , n20397 );
xor ( n20400 , n19465 , n19606 );
nor ( n20401 , n9518 , n20305 );
and ( n20402 , n20400 , n20401 );
xor ( n20403 , n20400 , n20401 );
xor ( n20404 , n19469 , n19604 );
nor ( n20405 , n9527 , n20305 );
and ( n20406 , n20404 , n20405 );
xor ( n20407 , n20404 , n20405 );
xor ( n20408 , n19473 , n19602 );
nor ( n20409 , n9536 , n20305 );
and ( n20410 , n20408 , n20409 );
xor ( n20411 , n20408 , n20409 );
xor ( n20412 , n19477 , n19600 );
nor ( n20413 , n9545 , n20305 );
and ( n20414 , n20412 , n20413 );
xor ( n20415 , n20412 , n20413 );
xor ( n20416 , n19481 , n19598 );
nor ( n20417 , n9554 , n20305 );
and ( n20418 , n20416 , n20417 );
xor ( n20419 , n20416 , n20417 );
xor ( n20420 , n19485 , n19596 );
nor ( n20421 , n9563 , n20305 );
and ( n20422 , n20420 , n20421 );
xor ( n20423 , n20420 , n20421 );
xor ( n20424 , n19489 , n19594 );
nor ( n20425 , n9572 , n20305 );
and ( n20426 , n20424 , n20425 );
xor ( n20427 , n20424 , n20425 );
xor ( n20428 , n19493 , n19592 );
nor ( n20429 , n9581 , n20305 );
and ( n20430 , n20428 , n20429 );
xor ( n20431 , n20428 , n20429 );
xor ( n20432 , n19497 , n19590 );
nor ( n20433 , n9590 , n20305 );
and ( n20434 , n20432 , n20433 );
xor ( n20435 , n20432 , n20433 );
xor ( n20436 , n19501 , n19588 );
nor ( n20437 , n9599 , n20305 );
and ( n20438 , n20436 , n20437 );
xor ( n20439 , n20436 , n20437 );
xor ( n20440 , n19505 , n19586 );
nor ( n20441 , n9608 , n20305 );
and ( n20442 , n20440 , n20441 );
xor ( n20443 , n20440 , n20441 );
xor ( n20444 , n19509 , n19584 );
nor ( n20445 , n9617 , n20305 );
and ( n20446 , n20444 , n20445 );
xor ( n20447 , n20444 , n20445 );
xor ( n20448 , n19513 , n19582 );
nor ( n20449 , n9626 , n20305 );
and ( n20450 , n20448 , n20449 );
xor ( n20451 , n20448 , n20449 );
xor ( n20452 , n19517 , n19580 );
nor ( n20453 , n9635 , n20305 );
and ( n20454 , n20452 , n20453 );
xor ( n20455 , n20452 , n20453 );
xor ( n20456 , n19521 , n19578 );
nor ( n20457 , n9644 , n20305 );
and ( n20458 , n20456 , n20457 );
xor ( n20459 , n20456 , n20457 );
xor ( n20460 , n19525 , n19576 );
nor ( n20461 , n9653 , n20305 );
and ( n20462 , n20460 , n20461 );
xor ( n20463 , n20460 , n20461 );
xor ( n20464 , n19529 , n19574 );
nor ( n20465 , n9662 , n20305 );
and ( n20466 , n20464 , n20465 );
xor ( n20467 , n20464 , n20465 );
xor ( n20468 , n19533 , n19572 );
nor ( n20469 , n9671 , n20305 );
and ( n20470 , n20468 , n20469 );
xor ( n20471 , n20468 , n20469 );
xor ( n20472 , n19537 , n19570 );
nor ( n20473 , n9680 , n20305 );
and ( n20474 , n20472 , n20473 );
xor ( n20475 , n20472 , n20473 );
xor ( n20476 , n19541 , n19568 );
nor ( n20477 , n9689 , n20305 );
and ( n20478 , n20476 , n20477 );
xor ( n20479 , n20476 , n20477 );
xor ( n20480 , n19545 , n19566 );
nor ( n20481 , n9698 , n20305 );
and ( n20482 , n20480 , n20481 );
xor ( n20483 , n20480 , n20481 );
xor ( n20484 , n19549 , n19564 );
nor ( n20485 , n9707 , n20305 );
and ( n20486 , n20484 , n20485 );
xor ( n20487 , n20484 , n20485 );
xor ( n20488 , n19553 , n19562 );
nor ( n20489 , n9716 , n20305 );
and ( n20490 , n20488 , n20489 );
xor ( n20491 , n20488 , n20489 );
xor ( n20492 , n19557 , n19560 );
nor ( n20493 , n9725 , n20305 );
and ( n20494 , n20492 , n20493 );
xor ( n20495 , n20492 , n20493 );
xor ( n20496 , n19558 , n19559 );
nor ( n20497 , n9734 , n20305 );
and ( n20498 , n20496 , n20497 );
xor ( n20499 , n20496 , n20497 );
nor ( n20500 , n9752 , n19367 );
nor ( n20501 , n9743 , n20305 );
and ( n20502 , n20500 , n20501 );
and ( n20503 , n20499 , n20502 );
or ( n20504 , n20498 , n20503 );
and ( n20505 , n20495 , n20504 );
or ( n20506 , n20494 , n20505 );
and ( n20507 , n20491 , n20506 );
or ( n20508 , n20490 , n20507 );
and ( n20509 , n20487 , n20508 );
or ( n20510 , n20486 , n20509 );
and ( n20511 , n20483 , n20510 );
or ( n20512 , n20482 , n20511 );
and ( n20513 , n20479 , n20512 );
or ( n20514 , n20478 , n20513 );
and ( n20515 , n20475 , n20514 );
or ( n20516 , n20474 , n20515 );
and ( n20517 , n20471 , n20516 );
or ( n20518 , n20470 , n20517 );
and ( n20519 , n20467 , n20518 );
or ( n20520 , n20466 , n20519 );
and ( n20521 , n20463 , n20520 );
or ( n20522 , n20462 , n20521 );
and ( n20523 , n20459 , n20522 );
or ( n20524 , n20458 , n20523 );
and ( n20525 , n20455 , n20524 );
or ( n20526 , n20454 , n20525 );
and ( n20527 , n20451 , n20526 );
or ( n20528 , n20450 , n20527 );
and ( n20529 , n20447 , n20528 );
or ( n20530 , n20446 , n20529 );
and ( n20531 , n20443 , n20530 );
or ( n20532 , n20442 , n20531 );
and ( n20533 , n20439 , n20532 );
or ( n20534 , n20438 , n20533 );
and ( n20535 , n20435 , n20534 );
or ( n20536 , n20434 , n20535 );
and ( n20537 , n20431 , n20536 );
or ( n20538 , n20430 , n20537 );
and ( n20539 , n20427 , n20538 );
or ( n20540 , n20426 , n20539 );
and ( n20541 , n20423 , n20540 );
or ( n20542 , n20422 , n20541 );
and ( n20543 , n20419 , n20542 );
or ( n20544 , n20418 , n20543 );
and ( n20545 , n20415 , n20544 );
or ( n20546 , n20414 , n20545 );
and ( n20547 , n20411 , n20546 );
or ( n20548 , n20410 , n20547 );
and ( n20549 , n20407 , n20548 );
or ( n20550 , n20406 , n20549 );
and ( n20551 , n20403 , n20550 );
or ( n20552 , n20402 , n20551 );
and ( n20553 , n20399 , n20552 );
or ( n20554 , n20398 , n20553 );
and ( n20555 , n20395 , n20554 );
or ( n20556 , n20394 , n20555 );
and ( n20557 , n20391 , n20556 );
or ( n20558 , n20390 , n20557 );
and ( n20559 , n20387 , n20558 );
or ( n20560 , n20386 , n20559 );
and ( n20561 , n20383 , n20560 );
or ( n20562 , n20382 , n20561 );
and ( n20563 , n20379 , n20562 );
or ( n20564 , n20378 , n20563 );
and ( n20565 , n20375 , n20564 );
or ( n20566 , n20374 , n20565 );
and ( n20567 , n20371 , n20566 );
or ( n20568 , n20370 , n20567 );
and ( n20569 , n20367 , n20568 );
or ( n20570 , n20366 , n20569 );
and ( n20571 , n20363 , n20570 );
or ( n20572 , n20362 , n20571 );
and ( n20573 , n20359 , n20572 );
or ( n20574 , n20358 , n20573 );
and ( n20575 , n20355 , n20574 );
or ( n20576 , n20354 , n20575 );
and ( n20577 , n20351 , n20576 );
or ( n20578 , n20350 , n20577 );
and ( n20579 , n20347 , n20578 );
or ( n20580 , n20346 , n20579 );
and ( n20581 , n20343 , n20580 );
or ( n20582 , n20342 , n20581 );
and ( n20583 , n20339 , n20582 );
or ( n20584 , n20338 , n20583 );
and ( n20585 , n20335 , n20584 );
or ( n20586 , n20334 , n20585 );
and ( n20587 , n20331 , n20586 );
or ( n20588 , n20330 , n20587 );
and ( n20589 , n20327 , n20588 );
or ( n20590 , n20326 , n20589 );
and ( n20591 , n20323 , n20590 );
or ( n20592 , n20322 , n20591 );
and ( n20593 , n20319 , n20592 );
or ( n20594 , n20318 , n20593 );
and ( n20595 , n20315 , n20594 );
or ( n20596 , n20314 , n20595 );
and ( n20597 , n20311 , n20596 );
or ( n20598 , n20310 , n20597 );
xor ( n20599 , n20307 , n20598 );
buf ( n20600 , n483 );
not ( n20601 , n20600 );
nor ( n20602 , n601 , n20601 );
buf ( n20603 , n20602 );
nor ( n20604 , n622 , n18734 );
xor ( n20605 , n20603 , n20604 );
buf ( n20606 , n20605 );
nor ( n20607 , n646 , n17828 );
xor ( n20608 , n20606 , n20607 );
and ( n20609 , n19659 , n19660 );
buf ( n20610 , n20609 );
xor ( n20611 , n20608 , n20610 );
nor ( n20612 , n684 , n16943 );
xor ( n20613 , n20611 , n20612 );
and ( n20614 , n19662 , n19663 );
and ( n20615 , n19664 , n19666 );
or ( n20616 , n20614 , n20615 );
xor ( n20617 , n20613 , n20616 );
nor ( n20618 , n733 , n16077 );
xor ( n20619 , n20617 , n20618 );
and ( n20620 , n19667 , n19668 );
and ( n20621 , n19669 , n19672 );
or ( n20622 , n20620 , n20621 );
xor ( n20623 , n20619 , n20622 );
nor ( n20624 , n796 , n15230 );
xor ( n20625 , n20623 , n20624 );
and ( n20626 , n19673 , n19674 );
and ( n20627 , n19675 , n19678 );
or ( n20628 , n20626 , n20627 );
xor ( n20629 , n20625 , n20628 );
nor ( n20630 , n868 , n14403 );
xor ( n20631 , n20629 , n20630 );
and ( n20632 , n19679 , n19680 );
and ( n20633 , n19681 , n19684 );
or ( n20634 , n20632 , n20633 );
xor ( n20635 , n20631 , n20634 );
nor ( n20636 , n958 , n13599 );
xor ( n20637 , n20635 , n20636 );
and ( n20638 , n19685 , n19686 );
and ( n20639 , n19687 , n19690 );
or ( n20640 , n20638 , n20639 );
xor ( n20641 , n20637 , n20640 );
nor ( n20642 , n1062 , n12808 );
xor ( n20643 , n20641 , n20642 );
and ( n20644 , n19691 , n19692 );
and ( n20645 , n19693 , n19696 );
or ( n20646 , n20644 , n20645 );
xor ( n20647 , n20643 , n20646 );
nor ( n20648 , n1176 , n12037 );
xor ( n20649 , n20647 , n20648 );
and ( n20650 , n19697 , n19698 );
and ( n20651 , n19699 , n19702 );
or ( n20652 , n20650 , n20651 );
xor ( n20653 , n20649 , n20652 );
nor ( n20654 , n1303 , n11282 );
xor ( n20655 , n20653 , n20654 );
and ( n20656 , n19703 , n19704 );
and ( n20657 , n19705 , n19708 );
or ( n20658 , n20656 , n20657 );
xor ( n20659 , n20655 , n20658 );
nor ( n20660 , n1445 , n10547 );
xor ( n20661 , n20659 , n20660 );
and ( n20662 , n19709 , n19710 );
and ( n20663 , n19711 , n19714 );
or ( n20664 , n20662 , n20663 );
xor ( n20665 , n20661 , n20664 );
nor ( n20666 , n1598 , n9829 );
xor ( n20667 , n20665 , n20666 );
and ( n20668 , n19715 , n19716 );
and ( n20669 , n19717 , n19720 );
or ( n20670 , n20668 , n20669 );
xor ( n20671 , n20667 , n20670 );
nor ( n20672 , n1766 , n8955 );
xor ( n20673 , n20671 , n20672 );
and ( n20674 , n19721 , n19722 );
and ( n20675 , n19723 , n19726 );
or ( n20676 , n20674 , n20675 );
xor ( n20677 , n20673 , n20676 );
nor ( n20678 , n1945 , n603 );
xor ( n20679 , n20677 , n20678 );
and ( n20680 , n19727 , n19728 );
and ( n20681 , n19729 , n19732 );
or ( n20682 , n20680 , n20681 );
xor ( n20683 , n20679 , n20682 );
nor ( n20684 , n2137 , n652 );
xor ( n20685 , n20683 , n20684 );
and ( n20686 , n19733 , n19734 );
and ( n20687 , n19735 , n19738 );
or ( n20688 , n20686 , n20687 );
xor ( n20689 , n20685 , n20688 );
nor ( n20690 , n2343 , n624 );
xor ( n20691 , n20689 , n20690 );
and ( n20692 , n19739 , n19740 );
and ( n20693 , n19741 , n19744 );
or ( n20694 , n20692 , n20693 );
xor ( n20695 , n20691 , n20694 );
nor ( n20696 , n2566 , n648 );
xor ( n20697 , n20695 , n20696 );
and ( n20698 , n19745 , n19746 );
and ( n20699 , n19747 , n19750 );
or ( n20700 , n20698 , n20699 );
xor ( n20701 , n20697 , n20700 );
nor ( n20702 , n2797 , n686 );
xor ( n20703 , n20701 , n20702 );
and ( n20704 , n19751 , n19752 );
and ( n20705 , n19753 , n19756 );
or ( n20706 , n20704 , n20705 );
xor ( n20707 , n20703 , n20706 );
nor ( n20708 , n3043 , n735 );
xor ( n20709 , n20707 , n20708 );
and ( n20710 , n19757 , n19758 );
and ( n20711 , n19759 , n19762 );
or ( n20712 , n20710 , n20711 );
xor ( n20713 , n20709 , n20712 );
nor ( n20714 , n3300 , n798 );
xor ( n20715 , n20713 , n20714 );
and ( n20716 , n19763 , n19764 );
and ( n20717 , n19765 , n19768 );
or ( n20718 , n20716 , n20717 );
xor ( n20719 , n20715 , n20718 );
nor ( n20720 , n3570 , n870 );
xor ( n20721 , n20719 , n20720 );
and ( n20722 , n19769 , n19770 );
and ( n20723 , n19771 , n19774 );
or ( n20724 , n20722 , n20723 );
xor ( n20725 , n20721 , n20724 );
nor ( n20726 , n3853 , n960 );
xor ( n20727 , n20725 , n20726 );
and ( n20728 , n19775 , n19776 );
and ( n20729 , n19777 , n19780 );
or ( n20730 , n20728 , n20729 );
xor ( n20731 , n20727 , n20730 );
nor ( n20732 , n4151 , n1064 );
xor ( n20733 , n20731 , n20732 );
and ( n20734 , n19781 , n19782 );
and ( n20735 , n19783 , n19786 );
or ( n20736 , n20734 , n20735 );
xor ( n20737 , n20733 , n20736 );
nor ( n20738 , n4458 , n1178 );
xor ( n20739 , n20737 , n20738 );
and ( n20740 , n19787 , n19788 );
and ( n20741 , n19789 , n19792 );
or ( n20742 , n20740 , n20741 );
xor ( n20743 , n20739 , n20742 );
nor ( n20744 , n4786 , n1305 );
xor ( n20745 , n20743 , n20744 );
and ( n20746 , n19793 , n19794 );
and ( n20747 , n19795 , n19798 );
or ( n20748 , n20746 , n20747 );
xor ( n20749 , n20745 , n20748 );
nor ( n20750 , n5126 , n1447 );
xor ( n20751 , n20749 , n20750 );
and ( n20752 , n19799 , n19800 );
and ( n20753 , n19801 , n19804 );
or ( n20754 , n20752 , n20753 );
xor ( n20755 , n20751 , n20754 );
nor ( n20756 , n5477 , n1600 );
xor ( n20757 , n20755 , n20756 );
and ( n20758 , n19805 , n19806 );
and ( n20759 , n19807 , n19810 );
or ( n20760 , n20758 , n20759 );
xor ( n20761 , n20757 , n20760 );
nor ( n20762 , n5838 , n1768 );
xor ( n20763 , n20761 , n20762 );
and ( n20764 , n19811 , n19812 );
and ( n20765 , n19813 , n19816 );
or ( n20766 , n20764 , n20765 );
xor ( n20767 , n20763 , n20766 );
nor ( n20768 , n6212 , n1947 );
xor ( n20769 , n20767 , n20768 );
and ( n20770 , n19817 , n19818 );
and ( n20771 , n19819 , n19822 );
or ( n20772 , n20770 , n20771 );
xor ( n20773 , n20769 , n20772 );
nor ( n20774 , n6596 , n2139 );
xor ( n20775 , n20773 , n20774 );
and ( n20776 , n19823 , n19824 );
and ( n20777 , n19825 , n19828 );
or ( n20778 , n20776 , n20777 );
xor ( n20779 , n20775 , n20778 );
nor ( n20780 , n6997 , n2345 );
xor ( n20781 , n20779 , n20780 );
and ( n20782 , n19829 , n19830 );
and ( n20783 , n19831 , n19834 );
or ( n20784 , n20782 , n20783 );
xor ( n20785 , n20781 , n20784 );
nor ( n20786 , n7413 , n2568 );
xor ( n20787 , n20785 , n20786 );
and ( n20788 , n19835 , n19836 );
and ( n20789 , n19837 , n19840 );
or ( n20790 , n20788 , n20789 );
xor ( n20791 , n20787 , n20790 );
nor ( n20792 , n7841 , n2799 );
xor ( n20793 , n20791 , n20792 );
and ( n20794 , n19841 , n19842 );
and ( n20795 , n19843 , n19846 );
or ( n20796 , n20794 , n20795 );
xor ( n20797 , n20793 , n20796 );
nor ( n20798 , n8281 , n3045 );
xor ( n20799 , n20797 , n20798 );
and ( n20800 , n19847 , n19848 );
and ( n20801 , n19849 , n19852 );
or ( n20802 , n20800 , n20801 );
xor ( n20803 , n20799 , n20802 );
nor ( n20804 , n8737 , n3302 );
xor ( n20805 , n20803 , n20804 );
and ( n20806 , n19853 , n19854 );
and ( n20807 , n19855 , n19858 );
or ( n20808 , n20806 , n20807 );
xor ( n20809 , n20805 , n20808 );
nor ( n20810 , n9420 , n3572 );
xor ( n20811 , n20809 , n20810 );
and ( n20812 , n19859 , n19860 );
and ( n20813 , n19861 , n19864 );
or ( n20814 , n20812 , n20813 );
xor ( n20815 , n20811 , n20814 );
nor ( n20816 , n10312 , n3855 );
xor ( n20817 , n20815 , n20816 );
and ( n20818 , n19865 , n19866 );
and ( n20819 , n19867 , n19870 );
or ( n20820 , n20818 , n20819 );
xor ( n20821 , n20817 , n20820 );
nor ( n20822 , n11041 , n4153 );
xor ( n20823 , n20821 , n20822 );
and ( n20824 , n19871 , n19872 );
and ( n20825 , n19873 , n19876 );
or ( n20826 , n20824 , n20825 );
xor ( n20827 , n20823 , n20826 );
nor ( n20828 , n11790 , n4460 );
xor ( n20829 , n20827 , n20828 );
and ( n20830 , n19877 , n19878 );
and ( n20831 , n19879 , n19882 );
or ( n20832 , n20830 , n20831 );
xor ( n20833 , n20829 , n20832 );
nor ( n20834 , n12555 , n4788 );
xor ( n20835 , n20833 , n20834 );
and ( n20836 , n19883 , n19884 );
and ( n20837 , n19885 , n19888 );
or ( n20838 , n20836 , n20837 );
xor ( n20839 , n20835 , n20838 );
nor ( n20840 , n13340 , n5128 );
xor ( n20841 , n20839 , n20840 );
and ( n20842 , n19889 , n19890 );
and ( n20843 , n19891 , n19894 );
or ( n20844 , n20842 , n20843 );
xor ( n20845 , n20841 , n20844 );
nor ( n20846 , n14138 , n5479 );
xor ( n20847 , n20845 , n20846 );
and ( n20848 , n19895 , n19896 );
and ( n20849 , n19897 , n19900 );
or ( n20850 , n20848 , n20849 );
xor ( n20851 , n20847 , n20850 );
nor ( n20852 , n14959 , n5840 );
xor ( n20853 , n20851 , n20852 );
and ( n20854 , n19901 , n19902 );
and ( n20855 , n19903 , n19906 );
or ( n20856 , n20854 , n20855 );
xor ( n20857 , n20853 , n20856 );
nor ( n20858 , n15800 , n6214 );
xor ( n20859 , n20857 , n20858 );
and ( n20860 , n19907 , n19908 );
and ( n20861 , n19909 , n19912 );
or ( n20862 , n20860 , n20861 );
xor ( n20863 , n20859 , n20862 );
nor ( n20864 , n16660 , n6598 );
xor ( n20865 , n20863 , n20864 );
and ( n20866 , n19913 , n19914 );
and ( n20867 , n19915 , n19918 );
or ( n20868 , n20866 , n20867 );
xor ( n20869 , n20865 , n20868 );
nor ( n20870 , n17539 , n6999 );
xor ( n20871 , n20869 , n20870 );
and ( n20872 , n19919 , n19920 );
and ( n20873 , n19921 , n19924 );
or ( n20874 , n20872 , n20873 );
xor ( n20875 , n20871 , n20874 );
nor ( n20876 , n18439 , n7415 );
xor ( n20877 , n20875 , n20876 );
and ( n20878 , n19925 , n19926 );
and ( n20879 , n19927 , n19930 );
or ( n20880 , n20878 , n20879 );
xor ( n20881 , n20877 , n20880 );
nor ( n20882 , n19356 , n7843 );
xor ( n20883 , n20881 , n20882 );
and ( n20884 , n19931 , n19932 );
and ( n20885 , n19933 , n19936 );
or ( n20886 , n20884 , n20885 );
xor ( n20887 , n20883 , n20886 );
nor ( n20888 , n20294 , n8283 );
xor ( n20889 , n20887 , n20888 );
and ( n20890 , n19937 , n19938 );
and ( n20891 , n19939 , n19942 );
or ( n20892 , n20890 , n20891 );
xor ( n20893 , n20889 , n20892 );
and ( n20894 , n20275 , n20279 );
and ( n20895 , n19953 , n20270 );
and ( n20896 , n20270 , n20280 );
and ( n20897 , n19953 , n20280 );
or ( n20898 , n20895 , n20896 , n20897 );
xor ( n20899 , n20894 , n20898 );
and ( n20900 , n19957 , n20166 );
and ( n20901 , n20166 , n20269 );
and ( n20902 , n19957 , n20269 );
or ( n20903 , n20900 , n20901 , n20902 );
and ( n20904 , n19961 , n20041 );
and ( n20905 , n20041 , n20165 );
and ( n20906 , n19961 , n20165 );
or ( n20907 , n20904 , n20905 , n20906 );
and ( n20908 , n20046 , n20093 );
and ( n20909 , n20093 , n20164 );
and ( n20910 , n20046 , n20164 );
or ( n20911 , n20908 , n20909 , n20910 );
and ( n20912 , n20098 , n20124 );
and ( n20913 , n20124 , n20163 );
and ( n20914 , n20098 , n20163 );
or ( n20915 , n20912 , n20913 , n20914 );
and ( n20916 , n20059 , n20075 );
and ( n20917 , n20075 , n20091 );
and ( n20918 , n20059 , n20091 );
or ( n20919 , n20916 , n20917 , n20918 );
and ( n20920 , n20102 , n20106 );
and ( n20921 , n20106 , n20123 );
and ( n20922 , n20102 , n20123 );
or ( n20923 , n20920 , n20921 , n20922 );
xor ( n20924 , n20919 , n20923 );
and ( n20925 , n20080 , n20084 );
and ( n20926 , n20084 , n20090 );
and ( n20927 , n20080 , n20090 );
or ( n20928 , n20925 , n20926 , n20927 );
and ( n20929 , n20070 , n20071 );
and ( n20930 , n20071 , n20073 );
and ( n20931 , n20070 , n20073 );
or ( n20932 , n20929 , n20930 , n20931 );
and ( n20933 , n3182 , n6132 );
and ( n20934 , n3545 , n5765 );
xor ( n20935 , n20933 , n20934 );
and ( n20936 , n3801 , n5408 );
xor ( n20937 , n20935 , n20936 );
xor ( n20938 , n20932 , n20937 );
and ( n20939 , n2462 , n7310 );
and ( n20940 , n2779 , n6971 );
xor ( n20941 , n20939 , n20940 );
and ( n20942 , n3024 , n6504 );
xor ( n20943 , n20941 , n20942 );
xor ( n20944 , n20938 , n20943 );
xor ( n20945 , n20928 , n20944 );
and ( n20946 , n20086 , n20087 );
and ( n20947 , n20087 , n20089 );
and ( n20948 , n20086 , n20089 );
or ( n20949 , n20946 , n20947 , n20948 );
and ( n20950 , n20112 , n20113 );
and ( n20951 , n20113 , n20115 );
and ( n20952 , n20112 , n20115 );
or ( n20953 , n20950 , n20951 , n20952 );
xor ( n20954 , n20949 , n20953 );
and ( n20955 , n1933 , n8669 );
and ( n20956 , n2120 , n8243 );
xor ( n20957 , n20955 , n20956 );
and ( n20958 , n2324 , n7662 );
xor ( n20959 , n20957 , n20958 );
xor ( n20960 , n20954 , n20959 );
xor ( n20961 , n20945 , n20960 );
xor ( n20962 , n20924 , n20961 );
xor ( n20963 , n20915 , n20962 );
and ( n20964 , n20129 , n20144 );
and ( n20965 , n20144 , n20162 );
and ( n20966 , n20129 , n20162 );
or ( n20967 , n20964 , n20965 , n20966 );
and ( n20968 , n20149 , n20154 );
and ( n20969 , n20154 , n20161 );
and ( n20970 , n20149 , n20161 );
or ( n20971 , n20968 , n20969 , n20970 );
and ( n20972 , n20157 , n20158 );
and ( n20973 , n20158 , n20160 );
and ( n20974 , n20157 , n20160 );
or ( n20975 , n20972 , n20973 , n20974 );
buf ( n20976 , n419 );
and ( n20977 , n599 , n20976 );
and ( n20978 , n608 , n20156 );
xor ( n20979 , n20977 , n20978 );
and ( n20980 , n611 , n19222 );
xor ( n20981 , n20979 , n20980 );
xor ( n20982 , n20975 , n20981 );
and ( n20983 , n632 , n18407 );
and ( n20984 , n671 , n17422 );
xor ( n20985 , n20983 , n20984 );
and ( n20986 , n715 , n16550 );
xor ( n20987 , n20985 , n20986 );
xor ( n20988 , n20982 , n20987 );
xor ( n20989 , n20971 , n20988 );
and ( n20990 , n20139 , n20140 );
and ( n20991 , n20140 , n20142 );
and ( n20992 , n20139 , n20142 );
or ( n20993 , n20990 , n20991 , n20992 );
and ( n20994 , n20150 , n20151 );
and ( n20995 , n20151 , n20153 );
and ( n20996 , n20150 , n20153 );
or ( n20997 , n20994 , n20995 , n20996 );
xor ( n20998 , n20993 , n20997 );
and ( n20999 , n783 , n15691 );
and ( n21000 , n856 , n14838 );
xor ( n21001 , n20999 , n21000 );
and ( n21002 , n925 , n14044 );
xor ( n21003 , n21001 , n21002 );
xor ( n21004 , n20998 , n21003 );
xor ( n21005 , n20989 , n21004 );
xor ( n21006 , n20967 , n21005 );
and ( n21007 , n20111 , n20116 );
and ( n21008 , n20116 , n20122 );
and ( n21009 , n20111 , n20122 );
or ( n21010 , n21007 , n21008 , n21009 );
and ( n21011 , n20133 , n20137 );
and ( n21012 , n20137 , n20143 );
and ( n21013 , n20133 , n20143 );
or ( n21014 , n21011 , n21012 , n21013 );
xor ( n21015 , n21010 , n21014 );
and ( n21016 , n20118 , n20119 );
and ( n21017 , n20119 , n20121 );
and ( n21018 , n20118 , n20121 );
or ( n21019 , n21016 , n21017 , n21018 );
and ( n21020 , n1047 , n13256 );
and ( n21021 , n1164 , n12531 );
xor ( n21022 , n21020 , n21021 );
and ( n21023 , n1287 , n11718 );
xor ( n21024 , n21022 , n21023 );
xor ( n21025 , n21019 , n21024 );
and ( n21026 , n1383 , n10977 );
and ( n21027 , n1580 , n10239 );
xor ( n21028 , n21026 , n21027 );
and ( n21029 , n1694 , n9348 );
xor ( n21030 , n21028 , n21029 );
xor ( n21031 , n21025 , n21030 );
xor ( n21032 , n21015 , n21031 );
xor ( n21033 , n21006 , n21032 );
xor ( n21034 , n20963 , n21033 );
xor ( n21035 , n20911 , n21034 );
and ( n21036 , n19974 , n20011 );
and ( n21037 , n20011 , n20039 );
and ( n21038 , n19974 , n20039 );
or ( n21039 , n21036 , n21037 , n21038 );
and ( n21040 , n20050 , n20054 );
and ( n21041 , n20054 , n20092 );
and ( n21042 , n20050 , n20092 );
or ( n21043 , n21040 , n21041 , n21042 );
xor ( n21044 , n21039 , n21043 );
and ( n21045 , n20016 , n20020 );
and ( n21046 , n20020 , n20038 );
and ( n21047 , n20016 , n20038 );
or ( n21048 , n21045 , n21046 , n21047 );
and ( n21049 , n19998 , n20003 );
and ( n21050 , n20003 , n20009 );
and ( n21051 , n19998 , n20009 );
or ( n21052 , n21049 , n21050 , n21051 );
and ( n21053 , n19988 , n19989 );
and ( n21054 , n19989 , n19991 );
and ( n21055 , n19988 , n19991 );
or ( n21056 , n21053 , n21054 , n21055 );
and ( n21057 , n19999 , n20000 );
and ( n21058 , n20000 , n20002 );
and ( n21059 , n19999 , n20002 );
or ( n21060 , n21057 , n21058 , n21059 );
xor ( n21061 , n21056 , n21060 );
and ( n21062 , n7385 , n2544 );
and ( n21063 , n7808 , n2298 );
xor ( n21064 , n21062 , n21063 );
and ( n21065 , n8079 , n2100 );
xor ( n21066 , n21064 , n21065 );
xor ( n21067 , n21061 , n21066 );
xor ( n21068 , n21052 , n21067 );
and ( n21069 , n20005 , n20006 );
and ( n21070 , n20006 , n20008 );
and ( n21071 , n20005 , n20008 );
or ( n21072 , n21069 , n21070 , n21071 );
and ( n21073 , n6187 , n3271 );
and ( n21074 , n6569 , n2981 );
xor ( n21075 , n21073 , n21074 );
and ( n21076 , n6816 , n2739 );
xor ( n21077 , n21075 , n21076 );
xor ( n21078 , n21072 , n21077 );
and ( n21079 , n4959 , n4102 );
and ( n21080 , n5459 , n3749 );
xor ( n21081 , n21079 , n21080 );
and ( n21082 , n5819 , n3495 );
xor ( n21083 , n21081 , n21082 );
xor ( n21084 , n21078 , n21083 );
xor ( n21085 , n21068 , n21084 );
xor ( n21086 , n21048 , n21085 );
and ( n21087 , n20027 , n20031 );
and ( n21088 , n20031 , n20037 );
and ( n21089 , n20027 , n20037 );
or ( n21090 , n21087 , n21088 , n21089 );
and ( n21091 , n20063 , n20068 );
and ( n21092 , n20068 , n20074 );
and ( n21093 , n20063 , n20074 );
or ( n21094 , n21091 , n21092 , n21093 );
xor ( n21095 , n21090 , n21094 );
and ( n21096 , n20033 , n20034 );
and ( n21097 , n20034 , n20036 );
and ( n21098 , n20033 , n20036 );
or ( n21099 , n21096 , n21097 , n21098 );
and ( n21100 , n20064 , n20065 );
and ( n21101 , n20065 , n20067 );
and ( n21102 , n20064 , n20067 );
or ( n21103 , n21100 , n21101 , n21102 );
xor ( n21104 , n21099 , n21103 );
and ( n21105 , n4132 , n5103 );
and ( n21106 , n4438 , n4730 );
xor ( n21107 , n21105 , n21106 );
and ( n21108 , n4766 , n4403 );
xor ( n21109 , n21107 , n21108 );
xor ( n21110 , n21104 , n21109 );
xor ( n21111 , n21095 , n21110 );
xor ( n21112 , n21086 , n21111 );
xor ( n21113 , n21044 , n21112 );
xor ( n21114 , n21035 , n21113 );
xor ( n21115 , n20907 , n21114 );
and ( n21116 , n19965 , n19969 );
and ( n21117 , n19969 , n20040 );
and ( n21118 , n19965 , n20040 );
or ( n21119 , n21116 , n21117 , n21118 );
and ( n21120 , n20180 , n20216 );
and ( n21121 , n20216 , n20267 );
and ( n21122 , n20180 , n20267 );
or ( n21123 , n21120 , n21121 , n21122 );
xor ( n21124 , n21119 , n21123 );
and ( n21125 , n20184 , n20188 );
and ( n21126 , n20188 , n20215 );
and ( n21127 , n20184 , n20215 );
or ( n21128 , n21125 , n21126 , n21127 );
and ( n21129 , n20193 , n20197 );
and ( n21130 , n20197 , n20214 );
and ( n21131 , n20193 , n20214 );
or ( n21132 , n21129 , n21130 , n21131 );
and ( n21133 , n19978 , n19993 );
and ( n21134 , n19993 , n20010 );
and ( n21135 , n19978 , n20010 );
or ( n21136 , n21133 , n21134 , n21135 );
xor ( n21137 , n21132 , n21136 );
and ( n21138 , n20202 , n20207 );
and ( n21139 , n20207 , n20213 );
and ( n21140 , n20202 , n20213 );
or ( n21141 , n21138 , n21139 , n21140 );
and ( n21142 , n19982 , n19986 );
and ( n21143 , n19986 , n19992 );
and ( n21144 , n19982 , n19992 );
or ( n21145 , n21142 , n21143 , n21144 );
xor ( n21146 , n21141 , n21145 );
and ( n21147 , n20209 , n20210 );
and ( n21148 , n20210 , n20212 );
and ( n21149 , n20209 , n20212 );
or ( n21150 , n21147 , n21148 , n21149 );
and ( n21151 , n11015 , n1424 );
and ( n21152 , n11769 , n1254 );
xor ( n21153 , n21151 , n21152 );
and ( n21154 , n12320 , n1134 );
xor ( n21155 , n21153 , n21154 );
xor ( n21156 , n21150 , n21155 );
and ( n21157 , n8718 , n1882 );
and ( n21158 , n9400 , n1738 );
xor ( n21159 , n21157 , n21158 );
and ( n21160 , n10291 , n1551 );
xor ( n21161 , n21159 , n21160 );
xor ( n21162 , n21156 , n21161 );
xor ( n21163 , n21146 , n21162 );
xor ( n21164 , n21137 , n21163 );
xor ( n21165 , n21128 , n21164 );
and ( n21166 , n20225 , n20242 );
and ( n21167 , n20242 , n20258 );
and ( n21168 , n20225 , n20258 );
or ( n21169 , n21166 , n21167 , n21168 );
and ( n21170 , n20247 , n20251 );
and ( n21171 , n20251 , n20257 );
and ( n21172 , n20247 , n20257 );
or ( n21173 , n21170 , n21171 , n21172 );
and ( n21174 , n20237 , n20238 );
and ( n21175 , n20238 , n20240 );
and ( n21176 , n20237 , n20240 );
or ( n21177 , n21174 , n21175 , n21176 );
and ( n21178 , n18144 , n635 );
and ( n21179 , n19324 , n606 );
xor ( n21180 , n21178 , n21179 );
and ( n21181 , n20233 , n615 );
xor ( n21182 , n21180 , n21181 );
xor ( n21183 , n21177 , n21182 );
and ( n21184 , n15758 , n771 );
and ( n21185 , n16637 , n719 );
xor ( n21186 , n21184 , n21185 );
and ( n21187 , n17512 , n663 );
xor ( n21188 , n21186 , n21187 );
xor ( n21189 , n21183 , n21188 );
xor ( n21190 , n21173 , n21189 );
and ( n21191 , n20253 , n20254 );
and ( n21192 , n20254 , n20256 );
and ( n21193 , n20253 , n20256 );
or ( n21194 , n21191 , n21192 , n21193 );
and ( n21195 , n20203 , n20204 );
and ( n21196 , n20204 , n20206 );
and ( n21197 , n20203 , n20206 );
or ( n21198 , n21195 , n21196 , n21197 );
xor ( n21199 , n21194 , n21198 );
and ( n21200 , n13322 , n1034 );
and ( n21201 , n14118 , n940 );
xor ( n21202 , n21200 , n21201 );
and ( n21203 , n14938 , n840 );
xor ( n21204 , n21202 , n21203 );
xor ( n21205 , n21199 , n21204 );
xor ( n21206 , n21190 , n21205 );
xor ( n21207 , n21169 , n21206 );
and ( n21208 , n20229 , n20235 );
and ( n21209 , n20235 , n20241 );
and ( n21210 , n20229 , n20241 );
or ( n21211 , n21208 , n21209 , n21210 );
and ( n21212 , n20230 , n20231 );
and ( n21213 , n20231 , n20234 );
and ( n21214 , n20230 , n20234 );
or ( n21215 , n21212 , n21213 , n21214 );
buf ( n21216 , n419 );
and ( n21217 , n21216 , n612 );
xor ( n21218 , n21215 , n21217 );
xor ( n21219 , n21211 , n21218 );
xor ( n21220 , n21207 , n21219 );
xor ( n21221 , n21165 , n21220 );
xor ( n21222 , n21124 , n21221 );
xor ( n21223 , n21115 , n21222 );
xor ( n21224 , n20903 , n21223 );
and ( n21225 , n20171 , n20175 );
and ( n21226 , n20175 , n20268 );
and ( n21227 , n20171 , n20268 );
or ( n21228 , n21225 , n21226 , n21227 );
and ( n21229 , n20261 , n20265 );
and ( n21230 , n20221 , n20259 );
and ( n21231 , n20259 , n20266 );
and ( n21232 , n20221 , n20266 );
or ( n21233 , n21230 , n21231 , n21232 );
xor ( n21234 , n21229 , n21233 );
xor ( n21235 , n21228 , n21234 );
xor ( n21236 , n21224 , n21235 );
xor ( n21237 , n20899 , n21236 );
and ( n21238 , n19944 , n19948 );
and ( n21239 , n19948 , n20281 );
and ( n21240 , n19944 , n20281 );
or ( n21241 , n21238 , n21239 , n21240 );
xor ( n21242 , n21237 , n21241 );
and ( n21243 , n20282 , n20286 );
and ( n21244 , n20287 , n20290 );
or ( n21245 , n21243 , n21244 );
xor ( n21246 , n21242 , n21245 );
buf ( n21247 , n21246 );
buf ( n21248 , n21247 );
not ( n21249 , n21248 );
nor ( n21250 , n21249 , n8739 );
xor ( n21251 , n20893 , n21250 );
and ( n21252 , n19943 , n20295 );
and ( n21253 , n20296 , n20299 );
or ( n21254 , n21252 , n21253 );
xor ( n21255 , n21251 , n21254 );
buf ( n21256 , n21255 );
buf ( n21257 , n21256 );
not ( n21258 , n21257 );
buf ( n21259 , n550 );
not ( n21260 , n21259 );
nor ( n21261 , n21258 , n21260 );
xor ( n21262 , n20599 , n21261 );
xor ( n21263 , n20311 , n20596 );
nor ( n21264 , n20303 , n21260 );
and ( n21265 , n21263 , n21264 );
xor ( n21266 , n21263 , n21264 );
xor ( n21267 , n20315 , n20594 );
nor ( n21268 , n19365 , n21260 );
and ( n21269 , n21267 , n21268 );
xor ( n21270 , n21267 , n21268 );
xor ( n21271 , n20319 , n20592 );
nor ( n21272 , n18448 , n21260 );
and ( n21273 , n21271 , n21272 );
xor ( n21274 , n21271 , n21272 );
xor ( n21275 , n20323 , n20590 );
nor ( n21276 , n17548 , n21260 );
and ( n21277 , n21275 , n21276 );
xor ( n21278 , n21275 , n21276 );
xor ( n21279 , n20327 , n20588 );
nor ( n21280 , n16669 , n21260 );
and ( n21281 , n21279 , n21280 );
xor ( n21282 , n21279 , n21280 );
xor ( n21283 , n20331 , n20586 );
nor ( n21284 , n15809 , n21260 );
and ( n21285 , n21283 , n21284 );
xor ( n21286 , n21283 , n21284 );
xor ( n21287 , n20335 , n20584 );
nor ( n21288 , n14968 , n21260 );
and ( n21289 , n21287 , n21288 );
xor ( n21290 , n21287 , n21288 );
xor ( n21291 , n20339 , n20582 );
nor ( n21292 , n14147 , n21260 );
and ( n21293 , n21291 , n21292 );
xor ( n21294 , n21291 , n21292 );
xor ( n21295 , n20343 , n20580 );
nor ( n21296 , n13349 , n21260 );
and ( n21297 , n21295 , n21296 );
xor ( n21298 , n21295 , n21296 );
xor ( n21299 , n20347 , n20578 );
nor ( n21300 , n12564 , n21260 );
and ( n21301 , n21299 , n21300 );
xor ( n21302 , n21299 , n21300 );
xor ( n21303 , n20351 , n20576 );
nor ( n21304 , n11799 , n21260 );
and ( n21305 , n21303 , n21304 );
xor ( n21306 , n21303 , n21304 );
xor ( n21307 , n20355 , n20574 );
nor ( n21308 , n11050 , n21260 );
and ( n21309 , n21307 , n21308 );
xor ( n21310 , n21307 , n21308 );
xor ( n21311 , n20359 , n20572 );
nor ( n21312 , n10321 , n21260 );
and ( n21313 , n21311 , n21312 );
xor ( n21314 , n21311 , n21312 );
xor ( n21315 , n20363 , n20570 );
nor ( n21316 , n9429 , n21260 );
and ( n21317 , n21315 , n21316 );
xor ( n21318 , n21315 , n21316 );
xor ( n21319 , n20367 , n20568 );
nor ( n21320 , n8949 , n21260 );
and ( n21321 , n21319 , n21320 );
xor ( n21322 , n21319 , n21320 );
xor ( n21323 , n20371 , n20566 );
nor ( n21324 , n9437 , n21260 );
and ( n21325 , n21323 , n21324 );
xor ( n21326 , n21323 , n21324 );
xor ( n21327 , n20375 , n20564 );
nor ( n21328 , n9446 , n21260 );
and ( n21329 , n21327 , n21328 );
xor ( n21330 , n21327 , n21328 );
xor ( n21331 , n20379 , n20562 );
nor ( n21332 , n9455 , n21260 );
and ( n21333 , n21331 , n21332 );
xor ( n21334 , n21331 , n21332 );
xor ( n21335 , n20383 , n20560 );
nor ( n21336 , n9464 , n21260 );
and ( n21337 , n21335 , n21336 );
xor ( n21338 , n21335 , n21336 );
xor ( n21339 , n20387 , n20558 );
nor ( n21340 , n9473 , n21260 );
and ( n21341 , n21339 , n21340 );
xor ( n21342 , n21339 , n21340 );
xor ( n21343 , n20391 , n20556 );
nor ( n21344 , n9482 , n21260 );
and ( n21345 , n21343 , n21344 );
xor ( n21346 , n21343 , n21344 );
xor ( n21347 , n20395 , n20554 );
nor ( n21348 , n9491 , n21260 );
and ( n21349 , n21347 , n21348 );
xor ( n21350 , n21347 , n21348 );
xor ( n21351 , n20399 , n20552 );
nor ( n21352 , n9500 , n21260 );
and ( n21353 , n21351 , n21352 );
xor ( n21354 , n21351 , n21352 );
xor ( n21355 , n20403 , n20550 );
nor ( n21356 , n9509 , n21260 );
and ( n21357 , n21355 , n21356 );
xor ( n21358 , n21355 , n21356 );
xor ( n21359 , n20407 , n20548 );
nor ( n21360 , n9518 , n21260 );
and ( n21361 , n21359 , n21360 );
xor ( n21362 , n21359 , n21360 );
xor ( n21363 , n20411 , n20546 );
nor ( n21364 , n9527 , n21260 );
and ( n21365 , n21363 , n21364 );
xor ( n21366 , n21363 , n21364 );
xor ( n21367 , n20415 , n20544 );
nor ( n21368 , n9536 , n21260 );
and ( n21369 , n21367 , n21368 );
xor ( n21370 , n21367 , n21368 );
xor ( n21371 , n20419 , n20542 );
nor ( n21372 , n9545 , n21260 );
and ( n21373 , n21371 , n21372 );
xor ( n21374 , n21371 , n21372 );
xor ( n21375 , n20423 , n20540 );
nor ( n21376 , n9554 , n21260 );
and ( n21377 , n21375 , n21376 );
xor ( n21378 , n21375 , n21376 );
xor ( n21379 , n20427 , n20538 );
nor ( n21380 , n9563 , n21260 );
and ( n21381 , n21379 , n21380 );
xor ( n21382 , n21379 , n21380 );
xor ( n21383 , n20431 , n20536 );
nor ( n21384 , n9572 , n21260 );
and ( n21385 , n21383 , n21384 );
xor ( n21386 , n21383 , n21384 );
xor ( n21387 , n20435 , n20534 );
nor ( n21388 , n9581 , n21260 );
and ( n21389 , n21387 , n21388 );
xor ( n21390 , n21387 , n21388 );
xor ( n21391 , n20439 , n20532 );
nor ( n21392 , n9590 , n21260 );
and ( n21393 , n21391 , n21392 );
xor ( n21394 , n21391 , n21392 );
xor ( n21395 , n20443 , n20530 );
nor ( n21396 , n9599 , n21260 );
and ( n21397 , n21395 , n21396 );
xor ( n21398 , n21395 , n21396 );
xor ( n21399 , n20447 , n20528 );
nor ( n21400 , n9608 , n21260 );
and ( n21401 , n21399 , n21400 );
xor ( n21402 , n21399 , n21400 );
xor ( n21403 , n20451 , n20526 );
nor ( n21404 , n9617 , n21260 );
and ( n21405 , n21403 , n21404 );
xor ( n21406 , n21403 , n21404 );
xor ( n21407 , n20455 , n20524 );
nor ( n21408 , n9626 , n21260 );
and ( n21409 , n21407 , n21408 );
xor ( n21410 , n21407 , n21408 );
xor ( n21411 , n20459 , n20522 );
nor ( n21412 , n9635 , n21260 );
and ( n21413 , n21411 , n21412 );
xor ( n21414 , n21411 , n21412 );
xor ( n21415 , n20463 , n20520 );
nor ( n21416 , n9644 , n21260 );
and ( n21417 , n21415 , n21416 );
xor ( n21418 , n21415 , n21416 );
xor ( n21419 , n20467 , n20518 );
nor ( n21420 , n9653 , n21260 );
and ( n21421 , n21419 , n21420 );
xor ( n21422 , n21419 , n21420 );
xor ( n21423 , n20471 , n20516 );
nor ( n21424 , n9662 , n21260 );
and ( n21425 , n21423 , n21424 );
xor ( n21426 , n21423 , n21424 );
xor ( n21427 , n20475 , n20514 );
nor ( n21428 , n9671 , n21260 );
and ( n21429 , n21427 , n21428 );
xor ( n21430 , n21427 , n21428 );
xor ( n21431 , n20479 , n20512 );
nor ( n21432 , n9680 , n21260 );
and ( n21433 , n21431 , n21432 );
xor ( n21434 , n21431 , n21432 );
xor ( n21435 , n20483 , n20510 );
nor ( n21436 , n9689 , n21260 );
and ( n21437 , n21435 , n21436 );
xor ( n21438 , n21435 , n21436 );
xor ( n21439 , n20487 , n20508 );
nor ( n21440 , n9698 , n21260 );
and ( n21441 , n21439 , n21440 );
xor ( n21442 , n21439 , n21440 );
xor ( n21443 , n20491 , n20506 );
nor ( n21444 , n9707 , n21260 );
and ( n21445 , n21443 , n21444 );
xor ( n21446 , n21443 , n21444 );
xor ( n21447 , n20495 , n20504 );
nor ( n21448 , n9716 , n21260 );
and ( n21449 , n21447 , n21448 );
xor ( n21450 , n21447 , n21448 );
xor ( n21451 , n20499 , n20502 );
nor ( n21452 , n9725 , n21260 );
and ( n21453 , n21451 , n21452 );
xor ( n21454 , n21451 , n21452 );
xor ( n21455 , n20500 , n20501 );
nor ( n21456 , n9734 , n21260 );
and ( n21457 , n21455 , n21456 );
xor ( n21458 , n21455 , n21456 );
nor ( n21459 , n9752 , n20305 );
nor ( n21460 , n9743 , n21260 );
and ( n21461 , n21459 , n21460 );
and ( n21462 , n21458 , n21461 );
or ( n21463 , n21457 , n21462 );
and ( n21464 , n21454 , n21463 );
or ( n21465 , n21453 , n21464 );
and ( n21466 , n21450 , n21465 );
or ( n21467 , n21449 , n21466 );
and ( n21468 , n21446 , n21467 );
or ( n21469 , n21445 , n21468 );
and ( n21470 , n21442 , n21469 );
or ( n21471 , n21441 , n21470 );
and ( n21472 , n21438 , n21471 );
or ( n21473 , n21437 , n21472 );
and ( n21474 , n21434 , n21473 );
or ( n21475 , n21433 , n21474 );
and ( n21476 , n21430 , n21475 );
or ( n21477 , n21429 , n21476 );
and ( n21478 , n21426 , n21477 );
or ( n21479 , n21425 , n21478 );
and ( n21480 , n21422 , n21479 );
or ( n21481 , n21421 , n21480 );
and ( n21482 , n21418 , n21481 );
or ( n21483 , n21417 , n21482 );
and ( n21484 , n21414 , n21483 );
or ( n21485 , n21413 , n21484 );
and ( n21486 , n21410 , n21485 );
or ( n21487 , n21409 , n21486 );
and ( n21488 , n21406 , n21487 );
or ( n21489 , n21405 , n21488 );
and ( n21490 , n21402 , n21489 );
or ( n21491 , n21401 , n21490 );
and ( n21492 , n21398 , n21491 );
or ( n21493 , n21397 , n21492 );
and ( n21494 , n21394 , n21493 );
or ( n21495 , n21393 , n21494 );
and ( n21496 , n21390 , n21495 );
or ( n21497 , n21389 , n21496 );
and ( n21498 , n21386 , n21497 );
or ( n21499 , n21385 , n21498 );
and ( n21500 , n21382 , n21499 );
or ( n21501 , n21381 , n21500 );
and ( n21502 , n21378 , n21501 );
or ( n21503 , n21377 , n21502 );
and ( n21504 , n21374 , n21503 );
or ( n21505 , n21373 , n21504 );
and ( n21506 , n21370 , n21505 );
or ( n21507 , n21369 , n21506 );
and ( n21508 , n21366 , n21507 );
or ( n21509 , n21365 , n21508 );
and ( n21510 , n21362 , n21509 );
or ( n21511 , n21361 , n21510 );
and ( n21512 , n21358 , n21511 );
or ( n21513 , n21357 , n21512 );
and ( n21514 , n21354 , n21513 );
or ( n21515 , n21353 , n21514 );
and ( n21516 , n21350 , n21515 );
or ( n21517 , n21349 , n21516 );
and ( n21518 , n21346 , n21517 );
or ( n21519 , n21345 , n21518 );
and ( n21520 , n21342 , n21519 );
or ( n21521 , n21341 , n21520 );
and ( n21522 , n21338 , n21521 );
or ( n21523 , n21337 , n21522 );
and ( n21524 , n21334 , n21523 );
or ( n21525 , n21333 , n21524 );
and ( n21526 , n21330 , n21525 );
or ( n21527 , n21329 , n21526 );
and ( n21528 , n21326 , n21527 );
or ( n21529 , n21325 , n21528 );
and ( n21530 , n21322 , n21529 );
or ( n21531 , n21321 , n21530 );
and ( n21532 , n21318 , n21531 );
or ( n21533 , n21317 , n21532 );
and ( n21534 , n21314 , n21533 );
or ( n21535 , n21313 , n21534 );
and ( n21536 , n21310 , n21535 );
or ( n21537 , n21309 , n21536 );
and ( n21538 , n21306 , n21537 );
or ( n21539 , n21305 , n21538 );
and ( n21540 , n21302 , n21539 );
or ( n21541 , n21301 , n21540 );
and ( n21542 , n21298 , n21541 );
or ( n21543 , n21297 , n21542 );
and ( n21544 , n21294 , n21543 );
or ( n21545 , n21293 , n21544 );
and ( n21546 , n21290 , n21545 );
or ( n21547 , n21289 , n21546 );
and ( n21548 , n21286 , n21547 );
or ( n21549 , n21285 , n21548 );
and ( n21550 , n21282 , n21549 );
or ( n21551 , n21281 , n21550 );
and ( n21552 , n21278 , n21551 );
or ( n21553 , n21277 , n21552 );
and ( n21554 , n21274 , n21553 );
or ( n21555 , n21273 , n21554 );
and ( n21556 , n21270 , n21555 );
or ( n21557 , n21269 , n21556 );
and ( n21558 , n21266 , n21557 );
or ( n21559 , n21265 , n21558 );
xor ( n21560 , n21262 , n21559 );
buf ( n21561 , n482 );
not ( n21562 , n21561 );
nor ( n21563 , n601 , n21562 );
buf ( n21564 , n21563 );
nor ( n21565 , n622 , n19657 );
xor ( n21566 , n21564 , n21565 );
buf ( n21567 , n21566 );
nor ( n21568 , n646 , n18734 );
xor ( n21569 , n21567 , n21568 );
and ( n21570 , n20603 , n20604 );
buf ( n21571 , n21570 );
xor ( n21572 , n21569 , n21571 );
nor ( n21573 , n684 , n17828 );
xor ( n21574 , n21572 , n21573 );
and ( n21575 , n20606 , n20607 );
and ( n21576 , n20608 , n20610 );
or ( n21577 , n21575 , n21576 );
xor ( n21578 , n21574 , n21577 );
nor ( n21579 , n733 , n16943 );
xor ( n21580 , n21578 , n21579 );
and ( n21581 , n20611 , n20612 );
and ( n21582 , n20613 , n20616 );
or ( n21583 , n21581 , n21582 );
xor ( n21584 , n21580 , n21583 );
nor ( n21585 , n796 , n16077 );
xor ( n21586 , n21584 , n21585 );
and ( n21587 , n20617 , n20618 );
and ( n21588 , n20619 , n20622 );
or ( n21589 , n21587 , n21588 );
xor ( n21590 , n21586 , n21589 );
nor ( n21591 , n868 , n15230 );
xor ( n21592 , n21590 , n21591 );
and ( n21593 , n20623 , n20624 );
and ( n21594 , n20625 , n20628 );
or ( n21595 , n21593 , n21594 );
xor ( n21596 , n21592 , n21595 );
nor ( n21597 , n958 , n14403 );
xor ( n21598 , n21596 , n21597 );
and ( n21599 , n20629 , n20630 );
and ( n21600 , n20631 , n20634 );
or ( n21601 , n21599 , n21600 );
xor ( n21602 , n21598 , n21601 );
nor ( n21603 , n1062 , n13599 );
xor ( n21604 , n21602 , n21603 );
and ( n21605 , n20635 , n20636 );
and ( n21606 , n20637 , n20640 );
or ( n21607 , n21605 , n21606 );
xor ( n21608 , n21604 , n21607 );
nor ( n21609 , n1176 , n12808 );
xor ( n21610 , n21608 , n21609 );
and ( n21611 , n20641 , n20642 );
and ( n21612 , n20643 , n20646 );
or ( n21613 , n21611 , n21612 );
xor ( n21614 , n21610 , n21613 );
nor ( n21615 , n1303 , n12037 );
xor ( n21616 , n21614 , n21615 );
and ( n21617 , n20647 , n20648 );
and ( n21618 , n20649 , n20652 );
or ( n21619 , n21617 , n21618 );
xor ( n21620 , n21616 , n21619 );
nor ( n21621 , n1445 , n11282 );
xor ( n21622 , n21620 , n21621 );
and ( n21623 , n20653 , n20654 );
and ( n21624 , n20655 , n20658 );
or ( n21625 , n21623 , n21624 );
xor ( n21626 , n21622 , n21625 );
nor ( n21627 , n1598 , n10547 );
xor ( n21628 , n21626 , n21627 );
and ( n21629 , n20659 , n20660 );
and ( n21630 , n20661 , n20664 );
or ( n21631 , n21629 , n21630 );
xor ( n21632 , n21628 , n21631 );
nor ( n21633 , n1766 , n9829 );
xor ( n21634 , n21632 , n21633 );
and ( n21635 , n20665 , n20666 );
and ( n21636 , n20667 , n20670 );
or ( n21637 , n21635 , n21636 );
xor ( n21638 , n21634 , n21637 );
nor ( n21639 , n1945 , n8955 );
xor ( n21640 , n21638 , n21639 );
and ( n21641 , n20671 , n20672 );
and ( n21642 , n20673 , n20676 );
or ( n21643 , n21641 , n21642 );
xor ( n21644 , n21640 , n21643 );
nor ( n21645 , n2137 , n603 );
xor ( n21646 , n21644 , n21645 );
and ( n21647 , n20677 , n20678 );
and ( n21648 , n20679 , n20682 );
or ( n21649 , n21647 , n21648 );
xor ( n21650 , n21646 , n21649 );
nor ( n21651 , n2343 , n652 );
xor ( n21652 , n21650 , n21651 );
and ( n21653 , n20683 , n20684 );
and ( n21654 , n20685 , n20688 );
or ( n21655 , n21653 , n21654 );
xor ( n21656 , n21652 , n21655 );
nor ( n21657 , n2566 , n624 );
xor ( n21658 , n21656 , n21657 );
and ( n21659 , n20689 , n20690 );
and ( n21660 , n20691 , n20694 );
or ( n21661 , n21659 , n21660 );
xor ( n21662 , n21658 , n21661 );
nor ( n21663 , n2797 , n648 );
xor ( n21664 , n21662 , n21663 );
and ( n21665 , n20695 , n20696 );
and ( n21666 , n20697 , n20700 );
or ( n21667 , n21665 , n21666 );
xor ( n21668 , n21664 , n21667 );
nor ( n21669 , n3043 , n686 );
xor ( n21670 , n21668 , n21669 );
and ( n21671 , n20701 , n20702 );
and ( n21672 , n20703 , n20706 );
or ( n21673 , n21671 , n21672 );
xor ( n21674 , n21670 , n21673 );
nor ( n21675 , n3300 , n735 );
xor ( n21676 , n21674 , n21675 );
and ( n21677 , n20707 , n20708 );
and ( n21678 , n20709 , n20712 );
or ( n21679 , n21677 , n21678 );
xor ( n21680 , n21676 , n21679 );
nor ( n21681 , n3570 , n798 );
xor ( n21682 , n21680 , n21681 );
and ( n21683 , n20713 , n20714 );
and ( n21684 , n20715 , n20718 );
or ( n21685 , n21683 , n21684 );
xor ( n21686 , n21682 , n21685 );
nor ( n21687 , n3853 , n870 );
xor ( n21688 , n21686 , n21687 );
and ( n21689 , n20719 , n20720 );
and ( n21690 , n20721 , n20724 );
or ( n21691 , n21689 , n21690 );
xor ( n21692 , n21688 , n21691 );
nor ( n21693 , n4151 , n960 );
xor ( n21694 , n21692 , n21693 );
and ( n21695 , n20725 , n20726 );
and ( n21696 , n20727 , n20730 );
or ( n21697 , n21695 , n21696 );
xor ( n21698 , n21694 , n21697 );
nor ( n21699 , n4458 , n1064 );
xor ( n21700 , n21698 , n21699 );
and ( n21701 , n20731 , n20732 );
and ( n21702 , n20733 , n20736 );
or ( n21703 , n21701 , n21702 );
xor ( n21704 , n21700 , n21703 );
nor ( n21705 , n4786 , n1178 );
xor ( n21706 , n21704 , n21705 );
and ( n21707 , n20737 , n20738 );
and ( n21708 , n20739 , n20742 );
or ( n21709 , n21707 , n21708 );
xor ( n21710 , n21706 , n21709 );
nor ( n21711 , n5126 , n1305 );
xor ( n21712 , n21710 , n21711 );
and ( n21713 , n20743 , n20744 );
and ( n21714 , n20745 , n20748 );
or ( n21715 , n21713 , n21714 );
xor ( n21716 , n21712 , n21715 );
nor ( n21717 , n5477 , n1447 );
xor ( n21718 , n21716 , n21717 );
and ( n21719 , n20749 , n20750 );
and ( n21720 , n20751 , n20754 );
or ( n21721 , n21719 , n21720 );
xor ( n21722 , n21718 , n21721 );
nor ( n21723 , n5838 , n1600 );
xor ( n21724 , n21722 , n21723 );
and ( n21725 , n20755 , n20756 );
and ( n21726 , n20757 , n20760 );
or ( n21727 , n21725 , n21726 );
xor ( n21728 , n21724 , n21727 );
nor ( n21729 , n6212 , n1768 );
xor ( n21730 , n21728 , n21729 );
and ( n21731 , n20761 , n20762 );
and ( n21732 , n20763 , n20766 );
or ( n21733 , n21731 , n21732 );
xor ( n21734 , n21730 , n21733 );
nor ( n21735 , n6596 , n1947 );
xor ( n21736 , n21734 , n21735 );
and ( n21737 , n20767 , n20768 );
and ( n21738 , n20769 , n20772 );
or ( n21739 , n21737 , n21738 );
xor ( n21740 , n21736 , n21739 );
nor ( n21741 , n6997 , n2139 );
xor ( n21742 , n21740 , n21741 );
and ( n21743 , n20773 , n20774 );
and ( n21744 , n20775 , n20778 );
or ( n21745 , n21743 , n21744 );
xor ( n21746 , n21742 , n21745 );
nor ( n21747 , n7413 , n2345 );
xor ( n21748 , n21746 , n21747 );
and ( n21749 , n20779 , n20780 );
and ( n21750 , n20781 , n20784 );
or ( n21751 , n21749 , n21750 );
xor ( n21752 , n21748 , n21751 );
nor ( n21753 , n7841 , n2568 );
xor ( n21754 , n21752 , n21753 );
and ( n21755 , n20785 , n20786 );
and ( n21756 , n20787 , n20790 );
or ( n21757 , n21755 , n21756 );
xor ( n21758 , n21754 , n21757 );
nor ( n21759 , n8281 , n2799 );
xor ( n21760 , n21758 , n21759 );
and ( n21761 , n20791 , n20792 );
and ( n21762 , n20793 , n20796 );
or ( n21763 , n21761 , n21762 );
xor ( n21764 , n21760 , n21763 );
nor ( n21765 , n8737 , n3045 );
xor ( n21766 , n21764 , n21765 );
and ( n21767 , n20797 , n20798 );
and ( n21768 , n20799 , n20802 );
or ( n21769 , n21767 , n21768 );
xor ( n21770 , n21766 , n21769 );
nor ( n21771 , n9420 , n3302 );
xor ( n21772 , n21770 , n21771 );
and ( n21773 , n20803 , n20804 );
and ( n21774 , n20805 , n20808 );
or ( n21775 , n21773 , n21774 );
xor ( n21776 , n21772 , n21775 );
nor ( n21777 , n10312 , n3572 );
xor ( n21778 , n21776 , n21777 );
and ( n21779 , n20809 , n20810 );
and ( n21780 , n20811 , n20814 );
or ( n21781 , n21779 , n21780 );
xor ( n21782 , n21778 , n21781 );
nor ( n21783 , n11041 , n3855 );
xor ( n21784 , n21782 , n21783 );
and ( n21785 , n20815 , n20816 );
and ( n21786 , n20817 , n20820 );
or ( n21787 , n21785 , n21786 );
xor ( n21788 , n21784 , n21787 );
nor ( n21789 , n11790 , n4153 );
xor ( n21790 , n21788 , n21789 );
and ( n21791 , n20821 , n20822 );
and ( n21792 , n20823 , n20826 );
or ( n21793 , n21791 , n21792 );
xor ( n21794 , n21790 , n21793 );
nor ( n21795 , n12555 , n4460 );
xor ( n21796 , n21794 , n21795 );
and ( n21797 , n20827 , n20828 );
and ( n21798 , n20829 , n20832 );
or ( n21799 , n21797 , n21798 );
xor ( n21800 , n21796 , n21799 );
nor ( n21801 , n13340 , n4788 );
xor ( n21802 , n21800 , n21801 );
and ( n21803 , n20833 , n20834 );
and ( n21804 , n20835 , n20838 );
or ( n21805 , n21803 , n21804 );
xor ( n21806 , n21802 , n21805 );
nor ( n21807 , n14138 , n5128 );
xor ( n21808 , n21806 , n21807 );
and ( n21809 , n20839 , n20840 );
and ( n21810 , n20841 , n20844 );
or ( n21811 , n21809 , n21810 );
xor ( n21812 , n21808 , n21811 );
nor ( n21813 , n14959 , n5479 );
xor ( n21814 , n21812 , n21813 );
and ( n21815 , n20845 , n20846 );
and ( n21816 , n20847 , n20850 );
or ( n21817 , n21815 , n21816 );
xor ( n21818 , n21814 , n21817 );
nor ( n21819 , n15800 , n5840 );
xor ( n21820 , n21818 , n21819 );
and ( n21821 , n20851 , n20852 );
and ( n21822 , n20853 , n20856 );
or ( n21823 , n21821 , n21822 );
xor ( n21824 , n21820 , n21823 );
nor ( n21825 , n16660 , n6214 );
xor ( n21826 , n21824 , n21825 );
and ( n21827 , n20857 , n20858 );
and ( n21828 , n20859 , n20862 );
or ( n21829 , n21827 , n21828 );
xor ( n21830 , n21826 , n21829 );
nor ( n21831 , n17539 , n6598 );
xor ( n21832 , n21830 , n21831 );
and ( n21833 , n20863 , n20864 );
and ( n21834 , n20865 , n20868 );
or ( n21835 , n21833 , n21834 );
xor ( n21836 , n21832 , n21835 );
nor ( n21837 , n18439 , n6999 );
xor ( n21838 , n21836 , n21837 );
and ( n21839 , n20869 , n20870 );
and ( n21840 , n20871 , n20874 );
or ( n21841 , n21839 , n21840 );
xor ( n21842 , n21838 , n21841 );
nor ( n21843 , n19356 , n7415 );
xor ( n21844 , n21842 , n21843 );
and ( n21845 , n20875 , n20876 );
and ( n21846 , n20877 , n20880 );
or ( n21847 , n21845 , n21846 );
xor ( n21848 , n21844 , n21847 );
nor ( n21849 , n20294 , n7843 );
xor ( n21850 , n21848 , n21849 );
and ( n21851 , n20881 , n20882 );
and ( n21852 , n20883 , n20886 );
or ( n21853 , n21851 , n21852 );
xor ( n21854 , n21850 , n21853 );
nor ( n21855 , n21249 , n8283 );
xor ( n21856 , n21854 , n21855 );
and ( n21857 , n20887 , n20888 );
and ( n21858 , n20889 , n20892 );
or ( n21859 , n21857 , n21858 );
xor ( n21860 , n21856 , n21859 );
and ( n21861 , n21228 , n21234 );
and ( n21862 , n20903 , n21223 );
and ( n21863 , n21223 , n21235 );
and ( n21864 , n20903 , n21235 );
or ( n21865 , n21862 , n21863 , n21864 );
xor ( n21866 , n21861 , n21865 );
and ( n21867 , n20907 , n21114 );
and ( n21868 , n21114 , n21222 );
and ( n21869 , n20907 , n21222 );
or ( n21870 , n21867 , n21868 , n21869 );
and ( n21871 , n20911 , n21034 );
and ( n21872 , n21034 , n21113 );
and ( n21873 , n20911 , n21113 );
or ( n21874 , n21871 , n21872 , n21873 );
and ( n21875 , n20915 , n20962 );
and ( n21876 , n20962 , n21033 );
and ( n21877 , n20915 , n21033 );
or ( n21878 , n21875 , n21876 , n21877 );
and ( n21879 , n20919 , n20923 );
and ( n21880 , n20923 , n20961 );
and ( n21881 , n20919 , n20961 );
or ( n21882 , n21879 , n21880 , n21881 );
and ( n21883 , n21048 , n21085 );
and ( n21884 , n21085 , n21111 );
and ( n21885 , n21048 , n21111 );
or ( n21886 , n21883 , n21884 , n21885 );
xor ( n21887 , n21882 , n21886 );
and ( n21888 , n21090 , n21094 );
and ( n21889 , n21094 , n21110 );
and ( n21890 , n21090 , n21110 );
or ( n21891 , n21888 , n21889 , n21890 );
and ( n21892 , n21072 , n21077 );
and ( n21893 , n21077 , n21083 );
and ( n21894 , n21072 , n21083 );
or ( n21895 , n21892 , n21893 , n21894 );
and ( n21896 , n21062 , n21063 );
and ( n21897 , n21063 , n21065 );
and ( n21898 , n21062 , n21065 );
or ( n21899 , n21896 , n21897 , n21898 );
and ( n21900 , n21073 , n21074 );
and ( n21901 , n21074 , n21076 );
and ( n21902 , n21073 , n21076 );
or ( n21903 , n21900 , n21901 , n21902 );
xor ( n21904 , n21899 , n21903 );
and ( n21905 , n7385 , n2739 );
and ( n21906 , n7808 , n2544 );
xor ( n21907 , n21905 , n21906 );
and ( n21908 , n8079 , n2298 );
xor ( n21909 , n21907 , n21908 );
xor ( n21910 , n21904 , n21909 );
xor ( n21911 , n21895 , n21910 );
and ( n21912 , n21079 , n21080 );
and ( n21913 , n21080 , n21082 );
and ( n21914 , n21079 , n21082 );
or ( n21915 , n21912 , n21913 , n21914 );
and ( n21916 , n6187 , n3495 );
and ( n21917 , n6569 , n3271 );
xor ( n21918 , n21916 , n21917 );
and ( n21919 , n6816 , n2981 );
xor ( n21920 , n21918 , n21919 );
xor ( n21921 , n21915 , n21920 );
and ( n21922 , n4959 , n4403 );
and ( n21923 , n5459 , n4102 );
xor ( n21924 , n21922 , n21923 );
and ( n21925 , n5819 , n3749 );
xor ( n21926 , n21924 , n21925 );
xor ( n21927 , n21921 , n21926 );
xor ( n21928 , n21911 , n21927 );
xor ( n21929 , n21891 , n21928 );
and ( n21930 , n21099 , n21103 );
and ( n21931 , n21103 , n21109 );
and ( n21932 , n21099 , n21109 );
or ( n21933 , n21930 , n21931 , n21932 );
and ( n21934 , n20932 , n20937 );
and ( n21935 , n20937 , n20943 );
and ( n21936 , n20932 , n20943 );
or ( n21937 , n21934 , n21935 , n21936 );
xor ( n21938 , n21933 , n21937 );
and ( n21939 , n20933 , n20934 );
and ( n21940 , n20934 , n20936 );
and ( n21941 , n20933 , n20936 );
or ( n21942 , n21939 , n21940 , n21941 );
and ( n21943 , n21105 , n21106 );
and ( n21944 , n21106 , n21108 );
and ( n21945 , n21105 , n21108 );
or ( n21946 , n21943 , n21944 , n21945 );
xor ( n21947 , n21942 , n21946 );
and ( n21948 , n4132 , n5408 );
and ( n21949 , n4438 , n5103 );
xor ( n21950 , n21948 , n21949 );
buf ( n21951 , n4766 );
xor ( n21952 , n21950 , n21951 );
xor ( n21953 , n21947 , n21952 );
xor ( n21954 , n21938 , n21953 );
xor ( n21955 , n21929 , n21954 );
xor ( n21956 , n21887 , n21955 );
xor ( n21957 , n21878 , n21956 );
and ( n21958 , n20967 , n21005 );
and ( n21959 , n21005 , n21032 );
and ( n21960 , n20967 , n21032 );
or ( n21961 , n21958 , n21959 , n21960 );
and ( n21962 , n21010 , n21014 );
and ( n21963 , n21014 , n21031 );
and ( n21964 , n21010 , n21031 );
or ( n21965 , n21962 , n21963 , n21964 );
and ( n21966 , n20928 , n20944 );
and ( n21967 , n20944 , n20960 );
and ( n21968 , n20928 , n20960 );
or ( n21969 , n21966 , n21967 , n21968 );
xor ( n21970 , n21965 , n21969 );
and ( n21971 , n20949 , n20953 );
and ( n21972 , n20953 , n20959 );
and ( n21973 , n20949 , n20959 );
or ( n21974 , n21971 , n21972 , n21973 );
and ( n21975 , n20939 , n20940 );
and ( n21976 , n20940 , n20942 );
and ( n21977 , n20939 , n20942 );
or ( n21978 , n21975 , n21976 , n21977 );
and ( n21979 , n2462 , n7662 );
and ( n21980 , n2779 , n7310 );
xor ( n21981 , n21979 , n21980 );
and ( n21982 , n3024 , n6971 );
xor ( n21983 , n21981 , n21982 );
xor ( n21984 , n21978 , n21983 );
and ( n21985 , n3182 , n6504 );
and ( n21986 , n3545 , n6132 );
xor ( n21987 , n21985 , n21986 );
and ( n21988 , n3801 , n5765 );
xor ( n21989 , n21987 , n21988 );
xor ( n21990 , n21984 , n21989 );
xor ( n21991 , n21974 , n21990 );
and ( n21992 , n20955 , n20956 );
and ( n21993 , n20956 , n20958 );
and ( n21994 , n20955 , n20958 );
or ( n21995 , n21992 , n21993 , n21994 );
and ( n21996 , n21026 , n21027 );
and ( n21997 , n21027 , n21029 );
and ( n21998 , n21026 , n21029 );
or ( n21999 , n21996 , n21997 , n21998 );
xor ( n22000 , n21995 , n21999 );
and ( n22001 , n1933 , n9348 );
and ( n22002 , n2120 , n8669 );
xor ( n22003 , n22001 , n22002 );
and ( n22004 , n2324 , n8243 );
xor ( n22005 , n22003 , n22004 );
xor ( n22006 , n22000 , n22005 );
xor ( n22007 , n21991 , n22006 );
xor ( n22008 , n21970 , n22007 );
xor ( n22009 , n21961 , n22008 );
and ( n22010 , n20971 , n20988 );
and ( n22011 , n20988 , n21004 );
and ( n22012 , n20971 , n21004 );
or ( n22013 , n22010 , n22011 , n22012 );
and ( n22014 , n20993 , n20997 );
and ( n22015 , n20997 , n21003 );
and ( n22016 , n20993 , n21003 );
or ( n22017 , n22014 , n22015 , n22016 );
and ( n22018 , n21019 , n21024 );
and ( n22019 , n21024 , n21030 );
and ( n22020 , n21019 , n21030 );
or ( n22021 , n22018 , n22019 , n22020 );
xor ( n22022 , n22017 , n22021 );
and ( n22023 , n21020 , n21021 );
and ( n22024 , n21021 , n21023 );
and ( n22025 , n21020 , n21023 );
or ( n22026 , n22023 , n22024 , n22025 );
and ( n22027 , n1047 , n14044 );
and ( n22028 , n1164 , n13256 );
xor ( n22029 , n22027 , n22028 );
and ( n22030 , n1287 , n12531 );
xor ( n22031 , n22029 , n22030 );
xor ( n22032 , n22026 , n22031 );
and ( n22033 , n1383 , n11718 );
and ( n22034 , n1580 , n10977 );
xor ( n22035 , n22033 , n22034 );
and ( n22036 , n1694 , n10239 );
xor ( n22037 , n22035 , n22036 );
xor ( n22038 , n22032 , n22037 );
xor ( n22039 , n22022 , n22038 );
xor ( n22040 , n22013 , n22039 );
and ( n22041 , n20975 , n20981 );
and ( n22042 , n20981 , n20987 );
and ( n22043 , n20975 , n20987 );
or ( n22044 , n22041 , n22042 , n22043 );
and ( n22045 , n20983 , n20984 );
and ( n22046 , n20984 , n20986 );
and ( n22047 , n20983 , n20986 );
or ( n22048 , n22045 , n22046 , n22047 );
and ( n22049 , n20999 , n21000 );
and ( n22050 , n21000 , n21002 );
and ( n22051 , n20999 , n21002 );
or ( n22052 , n22049 , n22050 , n22051 );
xor ( n22053 , n22048 , n22052 );
and ( n22054 , n783 , n16550 );
and ( n22055 , n856 , n15691 );
xor ( n22056 , n22054 , n22055 );
and ( n22057 , n925 , n14838 );
xor ( n22058 , n22056 , n22057 );
xor ( n22059 , n22053 , n22058 );
xor ( n22060 , n22044 , n22059 );
and ( n22061 , n20977 , n20978 );
and ( n22062 , n20978 , n20980 );
and ( n22063 , n20977 , n20980 );
or ( n22064 , n22061 , n22062 , n22063 );
buf ( n22065 , n418 );
and ( n22066 , n599 , n22065 );
and ( n22067 , n608 , n20976 );
xor ( n22068 , n22066 , n22067 );
and ( n22069 , n611 , n20156 );
xor ( n22070 , n22068 , n22069 );
xor ( n22071 , n22064 , n22070 );
and ( n22072 , n632 , n19222 );
and ( n22073 , n671 , n18407 );
xor ( n22074 , n22072 , n22073 );
and ( n22075 , n715 , n17422 );
xor ( n22076 , n22074 , n22075 );
xor ( n22077 , n22071 , n22076 );
xor ( n22078 , n22060 , n22077 );
xor ( n22079 , n22040 , n22078 );
xor ( n22080 , n22009 , n22079 );
xor ( n22081 , n21957 , n22080 );
xor ( n22082 , n21874 , n22081 );
and ( n22083 , n21039 , n21043 );
and ( n22084 , n21043 , n21112 );
and ( n22085 , n21039 , n21112 );
or ( n22086 , n22083 , n22084 , n22085 );
and ( n22087 , n21128 , n21164 );
and ( n22088 , n21164 , n21220 );
and ( n22089 , n21128 , n21220 );
or ( n22090 , n22087 , n22088 , n22089 );
xor ( n22091 , n22086 , n22090 );
and ( n22092 , n21132 , n21136 );
and ( n22093 , n21136 , n21163 );
and ( n22094 , n21132 , n21163 );
or ( n22095 , n22092 , n22093 , n22094 );
and ( n22096 , n21052 , n21067 );
and ( n22097 , n21067 , n21084 );
and ( n22098 , n21052 , n21084 );
or ( n22099 , n22096 , n22097 , n22098 );
and ( n22100 , n21141 , n21145 );
and ( n22101 , n21145 , n21162 );
and ( n22102 , n21141 , n21162 );
or ( n22103 , n22100 , n22101 , n22102 );
xor ( n22104 , n22099 , n22103 );
and ( n22105 , n21150 , n21155 );
and ( n22106 , n21155 , n21161 );
and ( n22107 , n21150 , n21161 );
or ( n22108 , n22105 , n22106 , n22107 );
and ( n22109 , n21056 , n21060 );
and ( n22110 , n21060 , n21066 );
and ( n22111 , n21056 , n21066 );
or ( n22112 , n22109 , n22110 , n22111 );
xor ( n22113 , n22108 , n22112 );
and ( n22114 , n21157 , n21158 );
and ( n22115 , n21158 , n21160 );
and ( n22116 , n21157 , n21160 );
or ( n22117 , n22114 , n22115 , n22116 );
and ( n22118 , n11015 , n1551 );
and ( n22119 , n11769 , n1424 );
xor ( n22120 , n22118 , n22119 );
and ( n22121 , n12320 , n1254 );
xor ( n22122 , n22120 , n22121 );
xor ( n22123 , n22117 , n22122 );
and ( n22124 , n8718 , n2100 );
and ( n22125 , n9400 , n1882 );
xor ( n22126 , n22124 , n22125 );
and ( n22127 , n10291 , n1738 );
xor ( n22128 , n22126 , n22127 );
xor ( n22129 , n22123 , n22128 );
xor ( n22130 , n22113 , n22129 );
xor ( n22131 , n22104 , n22130 );
xor ( n22132 , n22095 , n22131 );
and ( n22133 , n21173 , n21189 );
and ( n22134 , n21189 , n21205 );
and ( n22135 , n21173 , n21205 );
or ( n22136 , n22133 , n22134 , n22135 );
and ( n22137 , n21194 , n21198 );
and ( n22138 , n21198 , n21204 );
and ( n22139 , n21194 , n21204 );
or ( n22140 , n22137 , n22138 , n22139 );
and ( n22141 , n21184 , n21185 );
and ( n22142 , n21185 , n21187 );
and ( n22143 , n21184 , n21187 );
or ( n22144 , n22141 , n22142 , n22143 );
and ( n22145 , n18144 , n663 );
and ( n22146 , n19324 , n635 );
xor ( n22147 , n22145 , n22146 );
and ( n22148 , n20233 , n606 );
xor ( n22149 , n22147 , n22148 );
xor ( n22150 , n22144 , n22149 );
and ( n22151 , n15758 , n840 );
and ( n22152 , n16637 , n771 );
xor ( n22153 , n22151 , n22152 );
and ( n22154 , n17512 , n719 );
xor ( n22155 , n22153 , n22154 );
xor ( n22156 , n22150 , n22155 );
xor ( n22157 , n22140 , n22156 );
and ( n22158 , n21200 , n21201 );
and ( n22159 , n21201 , n21203 );
and ( n22160 , n21200 , n21203 );
or ( n22161 , n22158 , n22159 , n22160 );
and ( n22162 , n21151 , n21152 );
and ( n22163 , n21152 , n21154 );
and ( n22164 , n21151 , n21154 );
or ( n22165 , n22162 , n22163 , n22164 );
xor ( n22166 , n22161 , n22165 );
and ( n22167 , n13322 , n1134 );
and ( n22168 , n14118 , n1034 );
xor ( n22169 , n22167 , n22168 );
and ( n22170 , n14938 , n940 );
xor ( n22171 , n22169 , n22170 );
xor ( n22172 , n22166 , n22171 );
xor ( n22173 , n22157 , n22172 );
xor ( n22174 , n22136 , n22173 );
and ( n22175 , n21177 , n21182 );
and ( n22176 , n21182 , n21188 );
and ( n22177 , n21177 , n21188 );
or ( n22178 , n22175 , n22176 , n22177 );
and ( n22179 , n21215 , n21217 );
xor ( n22180 , n22178 , n22179 );
and ( n22181 , n21178 , n21179 );
and ( n22182 , n21179 , n21181 );
and ( n22183 , n21178 , n21181 );
or ( n22184 , n22181 , n22182 , n22183 );
and ( n22185 , n21216 , n615 );
buf ( n22186 , n418 );
and ( n22187 , n22186 , n612 );
xor ( n22188 , n22185 , n22187 );
xor ( n22189 , n22184 , n22188 );
xor ( n22190 , n22180 , n22189 );
xor ( n22191 , n22174 , n22190 );
xor ( n22192 , n22132 , n22191 );
xor ( n22193 , n22091 , n22192 );
xor ( n22194 , n22082 , n22193 );
xor ( n22195 , n21870 , n22194 );
and ( n22196 , n21119 , n21123 );
and ( n22197 , n21123 , n21221 );
and ( n22198 , n21119 , n21221 );
or ( n22199 , n22196 , n22197 , n22198 );
and ( n22200 , n21229 , n21233 );
and ( n22201 , n21211 , n21218 );
and ( n22202 , n21169 , n21206 );
and ( n22203 , n21206 , n21219 );
and ( n22204 , n21169 , n21219 );
or ( n22205 , n22202 , n22203 , n22204 );
xor ( n22206 , n22201 , n22205 );
xor ( n22207 , n22200 , n22206 );
xor ( n22208 , n22199 , n22207 );
xor ( n22209 , n22195 , n22208 );
xor ( n22210 , n21866 , n22209 );
and ( n22211 , n20894 , n20898 );
and ( n22212 , n20898 , n21236 );
and ( n22213 , n20894 , n21236 );
or ( n22214 , n22211 , n22212 , n22213 );
xor ( n22215 , n22210 , n22214 );
and ( n22216 , n21237 , n21241 );
and ( n22217 , n21242 , n21245 );
or ( n22218 , n22216 , n22217 );
xor ( n22219 , n22215 , n22218 );
buf ( n22220 , n22219 );
buf ( n22221 , n22220 );
not ( n22222 , n22221 );
nor ( n22223 , n22222 , n8739 );
xor ( n22224 , n21860 , n22223 );
and ( n22225 , n20893 , n21250 );
and ( n22226 , n21251 , n21254 );
or ( n22227 , n22225 , n22226 );
xor ( n22228 , n22224 , n22227 );
buf ( n22229 , n22228 );
buf ( n22230 , n22229 );
not ( n22231 , n22230 );
buf ( n22232 , n551 );
not ( n22233 , n22232 );
nor ( n22234 , n22231 , n22233 );
xor ( n22235 , n21560 , n22234 );
xor ( n22236 , n21266 , n21557 );
nor ( n22237 , n21258 , n22233 );
and ( n22238 , n22236 , n22237 );
xor ( n22239 , n22236 , n22237 );
xor ( n22240 , n21270 , n21555 );
nor ( n22241 , n20303 , n22233 );
and ( n22242 , n22240 , n22241 );
xor ( n22243 , n22240 , n22241 );
xor ( n22244 , n21274 , n21553 );
nor ( n22245 , n19365 , n22233 );
and ( n22246 , n22244 , n22245 );
xor ( n22247 , n22244 , n22245 );
xor ( n22248 , n21278 , n21551 );
nor ( n22249 , n18448 , n22233 );
and ( n22250 , n22248 , n22249 );
xor ( n22251 , n22248 , n22249 );
xor ( n22252 , n21282 , n21549 );
nor ( n22253 , n17548 , n22233 );
and ( n22254 , n22252 , n22253 );
xor ( n22255 , n22252 , n22253 );
xor ( n22256 , n21286 , n21547 );
nor ( n22257 , n16669 , n22233 );
and ( n22258 , n22256 , n22257 );
xor ( n22259 , n22256 , n22257 );
xor ( n22260 , n21290 , n21545 );
nor ( n22261 , n15809 , n22233 );
and ( n22262 , n22260 , n22261 );
xor ( n22263 , n22260 , n22261 );
xor ( n22264 , n21294 , n21543 );
nor ( n22265 , n14968 , n22233 );
and ( n22266 , n22264 , n22265 );
xor ( n22267 , n22264 , n22265 );
xor ( n22268 , n21298 , n21541 );
nor ( n22269 , n14147 , n22233 );
and ( n22270 , n22268 , n22269 );
xor ( n22271 , n22268 , n22269 );
xor ( n22272 , n21302 , n21539 );
nor ( n22273 , n13349 , n22233 );
and ( n22274 , n22272 , n22273 );
xor ( n22275 , n22272 , n22273 );
xor ( n22276 , n21306 , n21537 );
nor ( n22277 , n12564 , n22233 );
and ( n22278 , n22276 , n22277 );
xor ( n22279 , n22276 , n22277 );
xor ( n22280 , n21310 , n21535 );
nor ( n22281 , n11799 , n22233 );
and ( n22282 , n22280 , n22281 );
xor ( n22283 , n22280 , n22281 );
xor ( n22284 , n21314 , n21533 );
nor ( n22285 , n11050 , n22233 );
and ( n22286 , n22284 , n22285 );
xor ( n22287 , n22284 , n22285 );
xor ( n22288 , n21318 , n21531 );
nor ( n22289 , n10321 , n22233 );
and ( n22290 , n22288 , n22289 );
xor ( n22291 , n22288 , n22289 );
xor ( n22292 , n21322 , n21529 );
nor ( n22293 , n9429 , n22233 );
and ( n22294 , n22292 , n22293 );
xor ( n22295 , n22292 , n22293 );
xor ( n22296 , n21326 , n21527 );
nor ( n22297 , n8949 , n22233 );
and ( n22298 , n22296 , n22297 );
xor ( n22299 , n22296 , n22297 );
xor ( n22300 , n21330 , n21525 );
nor ( n22301 , n9437 , n22233 );
and ( n22302 , n22300 , n22301 );
xor ( n22303 , n22300 , n22301 );
xor ( n22304 , n21334 , n21523 );
nor ( n22305 , n9446 , n22233 );
and ( n22306 , n22304 , n22305 );
xor ( n22307 , n22304 , n22305 );
xor ( n22308 , n21338 , n21521 );
nor ( n22309 , n9455 , n22233 );
and ( n22310 , n22308 , n22309 );
xor ( n22311 , n22308 , n22309 );
xor ( n22312 , n21342 , n21519 );
nor ( n22313 , n9464 , n22233 );
and ( n22314 , n22312 , n22313 );
xor ( n22315 , n22312 , n22313 );
xor ( n22316 , n21346 , n21517 );
nor ( n22317 , n9473 , n22233 );
and ( n22318 , n22316 , n22317 );
xor ( n22319 , n22316 , n22317 );
xor ( n22320 , n21350 , n21515 );
nor ( n22321 , n9482 , n22233 );
and ( n22322 , n22320 , n22321 );
xor ( n22323 , n22320 , n22321 );
xor ( n22324 , n21354 , n21513 );
nor ( n22325 , n9491 , n22233 );
and ( n22326 , n22324 , n22325 );
xor ( n22327 , n22324 , n22325 );
xor ( n22328 , n21358 , n21511 );
nor ( n22329 , n9500 , n22233 );
and ( n22330 , n22328 , n22329 );
xor ( n22331 , n22328 , n22329 );
xor ( n22332 , n21362 , n21509 );
nor ( n22333 , n9509 , n22233 );
and ( n22334 , n22332 , n22333 );
xor ( n22335 , n22332 , n22333 );
xor ( n22336 , n21366 , n21507 );
nor ( n22337 , n9518 , n22233 );
and ( n22338 , n22336 , n22337 );
xor ( n22339 , n22336 , n22337 );
xor ( n22340 , n21370 , n21505 );
nor ( n22341 , n9527 , n22233 );
and ( n22342 , n22340 , n22341 );
xor ( n22343 , n22340 , n22341 );
xor ( n22344 , n21374 , n21503 );
nor ( n22345 , n9536 , n22233 );
and ( n22346 , n22344 , n22345 );
xor ( n22347 , n22344 , n22345 );
xor ( n22348 , n21378 , n21501 );
nor ( n22349 , n9545 , n22233 );
and ( n22350 , n22348 , n22349 );
xor ( n22351 , n22348 , n22349 );
xor ( n22352 , n21382 , n21499 );
nor ( n22353 , n9554 , n22233 );
and ( n22354 , n22352 , n22353 );
xor ( n22355 , n22352 , n22353 );
xor ( n22356 , n21386 , n21497 );
nor ( n22357 , n9563 , n22233 );
and ( n22358 , n22356 , n22357 );
xor ( n22359 , n22356 , n22357 );
xor ( n22360 , n21390 , n21495 );
nor ( n22361 , n9572 , n22233 );
and ( n22362 , n22360 , n22361 );
xor ( n22363 , n22360 , n22361 );
xor ( n22364 , n21394 , n21493 );
nor ( n22365 , n9581 , n22233 );
and ( n22366 , n22364 , n22365 );
xor ( n22367 , n22364 , n22365 );
xor ( n22368 , n21398 , n21491 );
nor ( n22369 , n9590 , n22233 );
and ( n22370 , n22368 , n22369 );
xor ( n22371 , n22368 , n22369 );
xor ( n22372 , n21402 , n21489 );
nor ( n22373 , n9599 , n22233 );
and ( n22374 , n22372 , n22373 );
xor ( n22375 , n22372 , n22373 );
xor ( n22376 , n21406 , n21487 );
nor ( n22377 , n9608 , n22233 );
and ( n22378 , n22376 , n22377 );
xor ( n22379 , n22376 , n22377 );
xor ( n22380 , n21410 , n21485 );
nor ( n22381 , n9617 , n22233 );
and ( n22382 , n22380 , n22381 );
xor ( n22383 , n22380 , n22381 );
xor ( n22384 , n21414 , n21483 );
nor ( n22385 , n9626 , n22233 );
and ( n22386 , n22384 , n22385 );
xor ( n22387 , n22384 , n22385 );
xor ( n22388 , n21418 , n21481 );
nor ( n22389 , n9635 , n22233 );
and ( n22390 , n22388 , n22389 );
xor ( n22391 , n22388 , n22389 );
xor ( n22392 , n21422 , n21479 );
nor ( n22393 , n9644 , n22233 );
and ( n22394 , n22392 , n22393 );
xor ( n22395 , n22392 , n22393 );
xor ( n22396 , n21426 , n21477 );
nor ( n22397 , n9653 , n22233 );
and ( n22398 , n22396 , n22397 );
xor ( n22399 , n22396 , n22397 );
xor ( n22400 , n21430 , n21475 );
nor ( n22401 , n9662 , n22233 );
and ( n22402 , n22400 , n22401 );
xor ( n22403 , n22400 , n22401 );
xor ( n22404 , n21434 , n21473 );
nor ( n22405 , n9671 , n22233 );
and ( n22406 , n22404 , n22405 );
xor ( n22407 , n22404 , n22405 );
xor ( n22408 , n21438 , n21471 );
nor ( n22409 , n9680 , n22233 );
and ( n22410 , n22408 , n22409 );
xor ( n22411 , n22408 , n22409 );
xor ( n22412 , n21442 , n21469 );
nor ( n22413 , n9689 , n22233 );
and ( n22414 , n22412 , n22413 );
xor ( n22415 , n22412 , n22413 );
xor ( n22416 , n21446 , n21467 );
nor ( n22417 , n9698 , n22233 );
and ( n22418 , n22416 , n22417 );
xor ( n22419 , n22416 , n22417 );
xor ( n22420 , n21450 , n21465 );
nor ( n22421 , n9707 , n22233 );
and ( n22422 , n22420 , n22421 );
xor ( n22423 , n22420 , n22421 );
xor ( n22424 , n21454 , n21463 );
nor ( n22425 , n9716 , n22233 );
and ( n22426 , n22424 , n22425 );
xor ( n22427 , n22424 , n22425 );
xor ( n22428 , n21458 , n21461 );
nor ( n22429 , n9725 , n22233 );
and ( n22430 , n22428 , n22429 );
xor ( n22431 , n22428 , n22429 );
xor ( n22432 , n21459 , n21460 );
nor ( n22433 , n9734 , n22233 );
and ( n22434 , n22432 , n22433 );
xor ( n22435 , n22432 , n22433 );
nor ( n22436 , n9752 , n21260 );
nor ( n22437 , n9743 , n22233 );
and ( n22438 , n22436 , n22437 );
and ( n22439 , n22435 , n22438 );
or ( n22440 , n22434 , n22439 );
and ( n22441 , n22431 , n22440 );
or ( n22442 , n22430 , n22441 );
and ( n22443 , n22427 , n22442 );
or ( n22444 , n22426 , n22443 );
and ( n22445 , n22423 , n22444 );
or ( n22446 , n22422 , n22445 );
and ( n22447 , n22419 , n22446 );
or ( n22448 , n22418 , n22447 );
and ( n22449 , n22415 , n22448 );
or ( n22450 , n22414 , n22449 );
and ( n22451 , n22411 , n22450 );
or ( n22452 , n22410 , n22451 );
and ( n22453 , n22407 , n22452 );
or ( n22454 , n22406 , n22453 );
and ( n22455 , n22403 , n22454 );
or ( n22456 , n22402 , n22455 );
and ( n22457 , n22399 , n22456 );
or ( n22458 , n22398 , n22457 );
and ( n22459 , n22395 , n22458 );
or ( n22460 , n22394 , n22459 );
and ( n22461 , n22391 , n22460 );
or ( n22462 , n22390 , n22461 );
and ( n22463 , n22387 , n22462 );
or ( n22464 , n22386 , n22463 );
and ( n22465 , n22383 , n22464 );
or ( n22466 , n22382 , n22465 );
and ( n22467 , n22379 , n22466 );
or ( n22468 , n22378 , n22467 );
and ( n22469 , n22375 , n22468 );
or ( n22470 , n22374 , n22469 );
and ( n22471 , n22371 , n22470 );
or ( n22472 , n22370 , n22471 );
and ( n22473 , n22367 , n22472 );
or ( n22474 , n22366 , n22473 );
and ( n22475 , n22363 , n22474 );
or ( n22476 , n22362 , n22475 );
and ( n22477 , n22359 , n22476 );
or ( n22478 , n22358 , n22477 );
and ( n22479 , n22355 , n22478 );
or ( n22480 , n22354 , n22479 );
and ( n22481 , n22351 , n22480 );
or ( n22482 , n22350 , n22481 );
and ( n22483 , n22347 , n22482 );
or ( n22484 , n22346 , n22483 );
and ( n22485 , n22343 , n22484 );
or ( n22486 , n22342 , n22485 );
and ( n22487 , n22339 , n22486 );
or ( n22488 , n22338 , n22487 );
and ( n22489 , n22335 , n22488 );
or ( n22490 , n22334 , n22489 );
and ( n22491 , n22331 , n22490 );
or ( n22492 , n22330 , n22491 );
and ( n22493 , n22327 , n22492 );
or ( n22494 , n22326 , n22493 );
and ( n22495 , n22323 , n22494 );
or ( n22496 , n22322 , n22495 );
and ( n22497 , n22319 , n22496 );
or ( n22498 , n22318 , n22497 );
and ( n22499 , n22315 , n22498 );
or ( n22500 , n22314 , n22499 );
and ( n22501 , n22311 , n22500 );
or ( n22502 , n22310 , n22501 );
and ( n22503 , n22307 , n22502 );
or ( n22504 , n22306 , n22503 );
and ( n22505 , n22303 , n22504 );
or ( n22506 , n22302 , n22505 );
and ( n22507 , n22299 , n22506 );
or ( n22508 , n22298 , n22507 );
and ( n22509 , n22295 , n22508 );
or ( n22510 , n22294 , n22509 );
and ( n22511 , n22291 , n22510 );
or ( n22512 , n22290 , n22511 );
and ( n22513 , n22287 , n22512 );
or ( n22514 , n22286 , n22513 );
and ( n22515 , n22283 , n22514 );
or ( n22516 , n22282 , n22515 );
and ( n22517 , n22279 , n22516 );
or ( n22518 , n22278 , n22517 );
and ( n22519 , n22275 , n22518 );
or ( n22520 , n22274 , n22519 );
and ( n22521 , n22271 , n22520 );
or ( n22522 , n22270 , n22521 );
and ( n22523 , n22267 , n22522 );
or ( n22524 , n22266 , n22523 );
and ( n22525 , n22263 , n22524 );
or ( n22526 , n22262 , n22525 );
and ( n22527 , n22259 , n22526 );
or ( n22528 , n22258 , n22527 );
and ( n22529 , n22255 , n22528 );
or ( n22530 , n22254 , n22529 );
and ( n22531 , n22251 , n22530 );
or ( n22532 , n22250 , n22531 );
and ( n22533 , n22247 , n22532 );
or ( n22534 , n22246 , n22533 );
and ( n22535 , n22243 , n22534 );
or ( n22536 , n22242 , n22535 );
and ( n22537 , n22239 , n22536 );
or ( n22538 , n22238 , n22537 );
xor ( n22539 , n22235 , n22538 );
buf ( n22540 , n481 );
not ( n22541 , n22540 );
nor ( n22542 , n601 , n22541 );
buf ( n22543 , n22542 );
nor ( n22544 , n622 , n20601 );
xor ( n22545 , n22543 , n22544 );
buf ( n22546 , n22545 );
nor ( n22547 , n646 , n19657 );
xor ( n22548 , n22546 , n22547 );
and ( n22549 , n21564 , n21565 );
buf ( n22550 , n22549 );
xor ( n22551 , n22548 , n22550 );
nor ( n22552 , n684 , n18734 );
xor ( n22553 , n22551 , n22552 );
and ( n22554 , n21567 , n21568 );
and ( n22555 , n21569 , n21571 );
or ( n22556 , n22554 , n22555 );
xor ( n22557 , n22553 , n22556 );
nor ( n22558 , n733 , n17828 );
xor ( n22559 , n22557 , n22558 );
and ( n22560 , n21572 , n21573 );
and ( n22561 , n21574 , n21577 );
or ( n22562 , n22560 , n22561 );
xor ( n22563 , n22559 , n22562 );
nor ( n22564 , n796 , n16943 );
xor ( n22565 , n22563 , n22564 );
and ( n22566 , n21578 , n21579 );
and ( n22567 , n21580 , n21583 );
or ( n22568 , n22566 , n22567 );
xor ( n22569 , n22565 , n22568 );
nor ( n22570 , n868 , n16077 );
xor ( n22571 , n22569 , n22570 );
and ( n22572 , n21584 , n21585 );
and ( n22573 , n21586 , n21589 );
or ( n22574 , n22572 , n22573 );
xor ( n22575 , n22571 , n22574 );
nor ( n22576 , n958 , n15230 );
xor ( n22577 , n22575 , n22576 );
and ( n22578 , n21590 , n21591 );
and ( n22579 , n21592 , n21595 );
or ( n22580 , n22578 , n22579 );
xor ( n22581 , n22577 , n22580 );
nor ( n22582 , n1062 , n14403 );
xor ( n22583 , n22581 , n22582 );
and ( n22584 , n21596 , n21597 );
and ( n22585 , n21598 , n21601 );
or ( n22586 , n22584 , n22585 );
xor ( n22587 , n22583 , n22586 );
nor ( n22588 , n1176 , n13599 );
xor ( n22589 , n22587 , n22588 );
and ( n22590 , n21602 , n21603 );
and ( n22591 , n21604 , n21607 );
or ( n22592 , n22590 , n22591 );
xor ( n22593 , n22589 , n22592 );
nor ( n22594 , n1303 , n12808 );
xor ( n22595 , n22593 , n22594 );
and ( n22596 , n21608 , n21609 );
and ( n22597 , n21610 , n21613 );
or ( n22598 , n22596 , n22597 );
xor ( n22599 , n22595 , n22598 );
nor ( n22600 , n1445 , n12037 );
xor ( n22601 , n22599 , n22600 );
and ( n22602 , n21614 , n21615 );
and ( n22603 , n21616 , n21619 );
or ( n22604 , n22602 , n22603 );
xor ( n22605 , n22601 , n22604 );
nor ( n22606 , n1598 , n11282 );
xor ( n22607 , n22605 , n22606 );
and ( n22608 , n21620 , n21621 );
and ( n22609 , n21622 , n21625 );
or ( n22610 , n22608 , n22609 );
xor ( n22611 , n22607 , n22610 );
nor ( n22612 , n1766 , n10547 );
xor ( n22613 , n22611 , n22612 );
and ( n22614 , n21626 , n21627 );
and ( n22615 , n21628 , n21631 );
or ( n22616 , n22614 , n22615 );
xor ( n22617 , n22613 , n22616 );
nor ( n22618 , n1945 , n9829 );
xor ( n22619 , n22617 , n22618 );
and ( n22620 , n21632 , n21633 );
and ( n22621 , n21634 , n21637 );
or ( n22622 , n22620 , n22621 );
xor ( n22623 , n22619 , n22622 );
nor ( n22624 , n2137 , n8955 );
xor ( n22625 , n22623 , n22624 );
and ( n22626 , n21638 , n21639 );
and ( n22627 , n21640 , n21643 );
or ( n22628 , n22626 , n22627 );
xor ( n22629 , n22625 , n22628 );
nor ( n22630 , n2343 , n603 );
xor ( n22631 , n22629 , n22630 );
and ( n22632 , n21644 , n21645 );
and ( n22633 , n21646 , n21649 );
or ( n22634 , n22632 , n22633 );
xor ( n22635 , n22631 , n22634 );
nor ( n22636 , n2566 , n652 );
xor ( n22637 , n22635 , n22636 );
and ( n22638 , n21650 , n21651 );
and ( n22639 , n21652 , n21655 );
or ( n22640 , n22638 , n22639 );
xor ( n22641 , n22637 , n22640 );
nor ( n22642 , n2797 , n624 );
xor ( n22643 , n22641 , n22642 );
and ( n22644 , n21656 , n21657 );
and ( n22645 , n21658 , n21661 );
or ( n22646 , n22644 , n22645 );
xor ( n22647 , n22643 , n22646 );
nor ( n22648 , n3043 , n648 );
xor ( n22649 , n22647 , n22648 );
and ( n22650 , n21662 , n21663 );
and ( n22651 , n21664 , n21667 );
or ( n22652 , n22650 , n22651 );
xor ( n22653 , n22649 , n22652 );
nor ( n22654 , n3300 , n686 );
xor ( n22655 , n22653 , n22654 );
and ( n22656 , n21668 , n21669 );
and ( n22657 , n21670 , n21673 );
or ( n22658 , n22656 , n22657 );
xor ( n22659 , n22655 , n22658 );
nor ( n22660 , n3570 , n735 );
xor ( n22661 , n22659 , n22660 );
and ( n22662 , n21674 , n21675 );
and ( n22663 , n21676 , n21679 );
or ( n22664 , n22662 , n22663 );
xor ( n22665 , n22661 , n22664 );
nor ( n22666 , n3853 , n798 );
xor ( n22667 , n22665 , n22666 );
and ( n22668 , n21680 , n21681 );
and ( n22669 , n21682 , n21685 );
or ( n22670 , n22668 , n22669 );
xor ( n22671 , n22667 , n22670 );
nor ( n22672 , n4151 , n870 );
xor ( n22673 , n22671 , n22672 );
and ( n22674 , n21686 , n21687 );
and ( n22675 , n21688 , n21691 );
or ( n22676 , n22674 , n22675 );
xor ( n22677 , n22673 , n22676 );
nor ( n22678 , n4458 , n960 );
xor ( n22679 , n22677 , n22678 );
and ( n22680 , n21692 , n21693 );
and ( n22681 , n21694 , n21697 );
or ( n22682 , n22680 , n22681 );
xor ( n22683 , n22679 , n22682 );
nor ( n22684 , n4786 , n1064 );
xor ( n22685 , n22683 , n22684 );
and ( n22686 , n21698 , n21699 );
and ( n22687 , n21700 , n21703 );
or ( n22688 , n22686 , n22687 );
xor ( n22689 , n22685 , n22688 );
nor ( n22690 , n5126 , n1178 );
xor ( n22691 , n22689 , n22690 );
and ( n22692 , n21704 , n21705 );
and ( n22693 , n21706 , n21709 );
or ( n22694 , n22692 , n22693 );
xor ( n22695 , n22691 , n22694 );
nor ( n22696 , n5477 , n1305 );
xor ( n22697 , n22695 , n22696 );
and ( n22698 , n21710 , n21711 );
and ( n22699 , n21712 , n21715 );
or ( n22700 , n22698 , n22699 );
xor ( n22701 , n22697 , n22700 );
nor ( n22702 , n5838 , n1447 );
xor ( n22703 , n22701 , n22702 );
and ( n22704 , n21716 , n21717 );
and ( n22705 , n21718 , n21721 );
or ( n22706 , n22704 , n22705 );
xor ( n22707 , n22703 , n22706 );
nor ( n22708 , n6212 , n1600 );
xor ( n22709 , n22707 , n22708 );
and ( n22710 , n21722 , n21723 );
and ( n22711 , n21724 , n21727 );
or ( n22712 , n22710 , n22711 );
xor ( n22713 , n22709 , n22712 );
nor ( n22714 , n6596 , n1768 );
xor ( n22715 , n22713 , n22714 );
and ( n22716 , n21728 , n21729 );
and ( n22717 , n21730 , n21733 );
or ( n22718 , n22716 , n22717 );
xor ( n22719 , n22715 , n22718 );
nor ( n22720 , n6997 , n1947 );
xor ( n22721 , n22719 , n22720 );
and ( n22722 , n21734 , n21735 );
and ( n22723 , n21736 , n21739 );
or ( n22724 , n22722 , n22723 );
xor ( n22725 , n22721 , n22724 );
nor ( n22726 , n7413 , n2139 );
xor ( n22727 , n22725 , n22726 );
and ( n22728 , n21740 , n21741 );
and ( n22729 , n21742 , n21745 );
or ( n22730 , n22728 , n22729 );
xor ( n22731 , n22727 , n22730 );
nor ( n22732 , n7841 , n2345 );
xor ( n22733 , n22731 , n22732 );
and ( n22734 , n21746 , n21747 );
and ( n22735 , n21748 , n21751 );
or ( n22736 , n22734 , n22735 );
xor ( n22737 , n22733 , n22736 );
nor ( n22738 , n8281 , n2568 );
xor ( n22739 , n22737 , n22738 );
and ( n22740 , n21752 , n21753 );
and ( n22741 , n21754 , n21757 );
or ( n22742 , n22740 , n22741 );
xor ( n22743 , n22739 , n22742 );
nor ( n22744 , n8737 , n2799 );
xor ( n22745 , n22743 , n22744 );
and ( n22746 , n21758 , n21759 );
and ( n22747 , n21760 , n21763 );
or ( n22748 , n22746 , n22747 );
xor ( n22749 , n22745 , n22748 );
nor ( n22750 , n9420 , n3045 );
xor ( n22751 , n22749 , n22750 );
and ( n22752 , n21764 , n21765 );
and ( n22753 , n21766 , n21769 );
or ( n22754 , n22752 , n22753 );
xor ( n22755 , n22751 , n22754 );
nor ( n22756 , n10312 , n3302 );
xor ( n22757 , n22755 , n22756 );
and ( n22758 , n21770 , n21771 );
and ( n22759 , n21772 , n21775 );
or ( n22760 , n22758 , n22759 );
xor ( n22761 , n22757 , n22760 );
nor ( n22762 , n11041 , n3572 );
xor ( n22763 , n22761 , n22762 );
and ( n22764 , n21776 , n21777 );
and ( n22765 , n21778 , n21781 );
or ( n22766 , n22764 , n22765 );
xor ( n22767 , n22763 , n22766 );
nor ( n22768 , n11790 , n3855 );
xor ( n22769 , n22767 , n22768 );
and ( n22770 , n21782 , n21783 );
and ( n22771 , n21784 , n21787 );
or ( n22772 , n22770 , n22771 );
xor ( n22773 , n22769 , n22772 );
nor ( n22774 , n12555 , n4153 );
xor ( n22775 , n22773 , n22774 );
and ( n22776 , n21788 , n21789 );
and ( n22777 , n21790 , n21793 );
or ( n22778 , n22776 , n22777 );
xor ( n22779 , n22775 , n22778 );
nor ( n22780 , n13340 , n4460 );
xor ( n22781 , n22779 , n22780 );
and ( n22782 , n21794 , n21795 );
and ( n22783 , n21796 , n21799 );
or ( n22784 , n22782 , n22783 );
xor ( n22785 , n22781 , n22784 );
nor ( n22786 , n14138 , n4788 );
xor ( n22787 , n22785 , n22786 );
and ( n22788 , n21800 , n21801 );
and ( n22789 , n21802 , n21805 );
or ( n22790 , n22788 , n22789 );
xor ( n22791 , n22787 , n22790 );
nor ( n22792 , n14959 , n5128 );
xor ( n22793 , n22791 , n22792 );
and ( n22794 , n21806 , n21807 );
and ( n22795 , n21808 , n21811 );
or ( n22796 , n22794 , n22795 );
xor ( n22797 , n22793 , n22796 );
nor ( n22798 , n15800 , n5479 );
xor ( n22799 , n22797 , n22798 );
and ( n22800 , n21812 , n21813 );
and ( n22801 , n21814 , n21817 );
or ( n22802 , n22800 , n22801 );
xor ( n22803 , n22799 , n22802 );
nor ( n22804 , n16660 , n5840 );
xor ( n22805 , n22803 , n22804 );
and ( n22806 , n21818 , n21819 );
and ( n22807 , n21820 , n21823 );
or ( n22808 , n22806 , n22807 );
xor ( n22809 , n22805 , n22808 );
nor ( n22810 , n17539 , n6214 );
xor ( n22811 , n22809 , n22810 );
and ( n22812 , n21824 , n21825 );
and ( n22813 , n21826 , n21829 );
or ( n22814 , n22812 , n22813 );
xor ( n22815 , n22811 , n22814 );
nor ( n22816 , n18439 , n6598 );
xor ( n22817 , n22815 , n22816 );
and ( n22818 , n21830 , n21831 );
and ( n22819 , n21832 , n21835 );
or ( n22820 , n22818 , n22819 );
xor ( n22821 , n22817 , n22820 );
nor ( n22822 , n19356 , n6999 );
xor ( n22823 , n22821 , n22822 );
and ( n22824 , n21836 , n21837 );
and ( n22825 , n21838 , n21841 );
or ( n22826 , n22824 , n22825 );
xor ( n22827 , n22823 , n22826 );
nor ( n22828 , n20294 , n7415 );
xor ( n22829 , n22827 , n22828 );
and ( n22830 , n21842 , n21843 );
and ( n22831 , n21844 , n21847 );
or ( n22832 , n22830 , n22831 );
xor ( n22833 , n22829 , n22832 );
nor ( n22834 , n21249 , n7843 );
xor ( n22835 , n22833 , n22834 );
and ( n22836 , n21848 , n21849 );
and ( n22837 , n21850 , n21853 );
or ( n22838 , n22836 , n22837 );
xor ( n22839 , n22835 , n22838 );
nor ( n22840 , n22222 , n8283 );
xor ( n22841 , n22839 , n22840 );
and ( n22842 , n21854 , n21855 );
and ( n22843 , n21856 , n21859 );
or ( n22844 , n22842 , n22843 );
xor ( n22845 , n22841 , n22844 );
and ( n22846 , n22199 , n22207 );
and ( n22847 , n21870 , n22194 );
and ( n22848 , n22194 , n22208 );
and ( n22849 , n21870 , n22208 );
or ( n22850 , n22847 , n22848 , n22849 );
xor ( n22851 , n22846 , n22850 );
and ( n22852 , n21874 , n22081 );
and ( n22853 , n22081 , n22193 );
and ( n22854 , n21874 , n22193 );
or ( n22855 , n22852 , n22853 , n22854 );
and ( n22856 , n21878 , n21956 );
and ( n22857 , n21956 , n22080 );
and ( n22858 , n21878 , n22080 );
or ( n22859 , n22856 , n22857 , n22858 );
and ( n22860 , n21882 , n21886 );
and ( n22861 , n21886 , n21955 );
and ( n22862 , n21882 , n21955 );
or ( n22863 , n22860 , n22861 , n22862 );
and ( n22864 , n22095 , n22131 );
and ( n22865 , n22131 , n22191 );
and ( n22866 , n22095 , n22191 );
or ( n22867 , n22864 , n22865 , n22866 );
xor ( n22868 , n22863 , n22867 );
and ( n22869 , n22099 , n22103 );
and ( n22870 , n22103 , n22130 );
and ( n22871 , n22099 , n22130 );
or ( n22872 , n22869 , n22870 , n22871 );
and ( n22873 , n22140 , n22156 );
and ( n22874 , n22156 , n22172 );
and ( n22875 , n22140 , n22172 );
or ( n22876 , n22873 , n22874 , n22875 );
and ( n22877 , n22144 , n22149 );
and ( n22878 , n22149 , n22155 );
and ( n22879 , n22144 , n22155 );
or ( n22880 , n22877 , n22878 , n22879 );
and ( n22881 , n22184 , n22188 );
xor ( n22882 , n22880 , n22881 );
and ( n22883 , n22145 , n22146 );
and ( n22884 , n22146 , n22148 );
and ( n22885 , n22145 , n22148 );
or ( n22886 , n22883 , n22884 , n22885 );
and ( n22887 , n22185 , n22187 );
xor ( n22888 , n22886 , n22887 );
and ( n22889 , n21216 , n606 );
and ( n22890 , n22186 , n615 );
xor ( n22891 , n22889 , n22890 );
buf ( n22892 , n417 );
and ( n22893 , n22892 , n612 );
xor ( n22894 , n22891 , n22893 );
xor ( n22895 , n22888 , n22894 );
xor ( n22896 , n22882 , n22895 );
xor ( n22897 , n22876 , n22896 );
and ( n22898 , n22161 , n22165 );
and ( n22899 , n22165 , n22171 );
and ( n22900 , n22161 , n22171 );
or ( n22901 , n22898 , n22899 , n22900 );
and ( n22902 , n22151 , n22152 );
and ( n22903 , n22152 , n22154 );
and ( n22904 , n22151 , n22154 );
or ( n22905 , n22902 , n22903 , n22904 );
and ( n22906 , n18144 , n719 );
and ( n22907 , n19324 , n663 );
xor ( n22908 , n22906 , n22907 );
and ( n22909 , n20233 , n635 );
xor ( n22910 , n22908 , n22909 );
xor ( n22911 , n22905 , n22910 );
and ( n22912 , n15758 , n940 );
and ( n22913 , n16637 , n840 );
xor ( n22914 , n22912 , n22913 );
and ( n22915 , n17512 , n771 );
xor ( n22916 , n22914 , n22915 );
xor ( n22917 , n22911 , n22916 );
xor ( n22918 , n22901 , n22917 );
and ( n22919 , n22167 , n22168 );
and ( n22920 , n22168 , n22170 );
and ( n22921 , n22167 , n22170 );
or ( n22922 , n22919 , n22920 , n22921 );
and ( n22923 , n22118 , n22119 );
and ( n22924 , n22119 , n22121 );
and ( n22925 , n22118 , n22121 );
or ( n22926 , n22923 , n22924 , n22925 );
xor ( n22927 , n22922 , n22926 );
and ( n22928 , n13322 , n1254 );
and ( n22929 , n14118 , n1134 );
xor ( n22930 , n22928 , n22929 );
and ( n22931 , n14938 , n1034 );
xor ( n22932 , n22930 , n22931 );
xor ( n22933 , n22927 , n22932 );
xor ( n22934 , n22918 , n22933 );
xor ( n22935 , n22897 , n22934 );
xor ( n22936 , n22872 , n22935 );
and ( n22937 , n22108 , n22112 );
and ( n22938 , n22112 , n22129 );
and ( n22939 , n22108 , n22129 );
or ( n22940 , n22937 , n22938 , n22939 );
and ( n22941 , n21895 , n21910 );
and ( n22942 , n21910 , n21927 );
and ( n22943 , n21895 , n21927 );
or ( n22944 , n22941 , n22942 , n22943 );
xor ( n22945 , n22940 , n22944 );
and ( n22946 , n22117 , n22122 );
and ( n22947 , n22122 , n22128 );
and ( n22948 , n22117 , n22128 );
or ( n22949 , n22946 , n22947 , n22948 );
and ( n22950 , n21899 , n21903 );
and ( n22951 , n21903 , n21909 );
and ( n22952 , n21899 , n21909 );
or ( n22953 , n22950 , n22951 , n22952 );
xor ( n22954 , n22949 , n22953 );
and ( n22955 , n22124 , n22125 );
and ( n22956 , n22125 , n22127 );
and ( n22957 , n22124 , n22127 );
or ( n22958 , n22955 , n22956 , n22957 );
and ( n22959 , n11015 , n1738 );
and ( n22960 , n11769 , n1551 );
xor ( n22961 , n22959 , n22960 );
and ( n22962 , n12320 , n1424 );
xor ( n22963 , n22961 , n22962 );
xor ( n22964 , n22958 , n22963 );
and ( n22965 , n8718 , n2298 );
and ( n22966 , n9400 , n2100 );
xor ( n22967 , n22965 , n22966 );
and ( n22968 , n10291 , n1882 );
xor ( n22969 , n22967 , n22968 );
xor ( n22970 , n22964 , n22969 );
xor ( n22971 , n22954 , n22970 );
xor ( n22972 , n22945 , n22971 );
xor ( n22973 , n22936 , n22972 );
xor ( n22974 , n22868 , n22973 );
xor ( n22975 , n22859 , n22974 );
and ( n22976 , n21961 , n22008 );
and ( n22977 , n22008 , n22079 );
and ( n22978 , n21961 , n22079 );
or ( n22979 , n22976 , n22977 , n22978 );
and ( n22980 , n21891 , n21928 );
and ( n22981 , n21928 , n21954 );
and ( n22982 , n21891 , n21954 );
or ( n22983 , n22980 , n22981 , n22982 );
and ( n22984 , n21965 , n21969 );
and ( n22985 , n21969 , n22007 );
and ( n22986 , n21965 , n22007 );
or ( n22987 , n22984 , n22985 , n22986 );
xor ( n22988 , n22983 , n22987 );
and ( n22989 , n21933 , n21937 );
and ( n22990 , n21937 , n21953 );
and ( n22991 , n21933 , n21953 );
or ( n22992 , n22989 , n22990 , n22991 );
and ( n22993 , n21942 , n21946 );
and ( n22994 , n21946 , n21952 );
and ( n22995 , n21942 , n21952 );
or ( n22996 , n22993 , n22994 , n22995 );
and ( n22997 , n21978 , n21983 );
and ( n22998 , n21983 , n21989 );
and ( n22999 , n21978 , n21989 );
or ( n23000 , n22997 , n22998 , n22999 );
xor ( n23001 , n22996 , n23000 );
and ( n23002 , n21948 , n21949 );
and ( n23003 , n21949 , n21951 );
and ( n23004 , n21948 , n21951 );
or ( n23005 , n23002 , n23003 , n23004 );
and ( n23006 , n21985 , n21986 );
and ( n23007 , n21986 , n21988 );
and ( n23008 , n21985 , n21988 );
or ( n23009 , n23006 , n23007 , n23008 );
xor ( n23010 , n23005 , n23009 );
and ( n23011 , n4132 , n5765 );
and ( n23012 , n4438 , n5408 );
xor ( n23013 , n23011 , n23012 );
and ( n23014 , n4766 , n5103 );
xor ( n23015 , n23013 , n23014 );
xor ( n23016 , n23010 , n23015 );
xor ( n23017 , n23001 , n23016 );
xor ( n23018 , n22992 , n23017 );
and ( n23019 , n21915 , n21920 );
and ( n23020 , n21920 , n21926 );
and ( n23021 , n21915 , n21926 );
or ( n23022 , n23019 , n23020 , n23021 );
and ( n23023 , n21905 , n21906 );
and ( n23024 , n21906 , n21908 );
and ( n23025 , n21905 , n21908 );
or ( n23026 , n23023 , n23024 , n23025 );
and ( n23027 , n21916 , n21917 );
and ( n23028 , n21917 , n21919 );
and ( n23029 , n21916 , n21919 );
or ( n23030 , n23027 , n23028 , n23029 );
xor ( n23031 , n23026 , n23030 );
and ( n23032 , n7385 , n2981 );
and ( n23033 , n7808 , n2739 );
xor ( n23034 , n23032 , n23033 );
and ( n23035 , n8079 , n2544 );
xor ( n23036 , n23034 , n23035 );
xor ( n23037 , n23031 , n23036 );
xor ( n23038 , n23022 , n23037 );
and ( n23039 , n21922 , n21923 );
and ( n23040 , n21923 , n21925 );
and ( n23041 , n21922 , n21925 );
or ( n23042 , n23039 , n23040 , n23041 );
and ( n23043 , n6187 , n3749 );
and ( n23044 , n6569 , n3495 );
xor ( n23045 , n23043 , n23044 );
and ( n23046 , n6816 , n3271 );
xor ( n23047 , n23045 , n23046 );
xor ( n23048 , n23042 , n23047 );
and ( n23049 , n4959 , n4730 );
and ( n23050 , n5459 , n4403 );
xor ( n23051 , n23049 , n23050 );
and ( n23052 , n5819 , n4102 );
xor ( n23053 , n23051 , n23052 );
xor ( n23054 , n23048 , n23053 );
xor ( n23055 , n23038 , n23054 );
xor ( n23056 , n23018 , n23055 );
xor ( n23057 , n22988 , n23056 );
xor ( n23058 , n22979 , n23057 );
and ( n23059 , n22013 , n22039 );
and ( n23060 , n22039 , n22078 );
and ( n23061 , n22013 , n22078 );
or ( n23062 , n23059 , n23060 , n23061 );
and ( n23063 , n22044 , n22059 );
and ( n23064 , n22059 , n22077 );
and ( n23065 , n22044 , n22077 );
or ( n23066 , n23063 , n23064 , n23065 );
and ( n23067 , n22064 , n22070 );
and ( n23068 , n22070 , n22076 );
and ( n23069 , n22064 , n22076 );
or ( n23070 , n23067 , n23068 , n23069 );
and ( n23071 , n22066 , n22067 );
and ( n23072 , n22067 , n22069 );
and ( n23073 , n22066 , n22069 );
or ( n23074 , n23071 , n23072 , n23073 );
buf ( n23075 , n417 );
and ( n23076 , n599 , n23075 );
and ( n23077 , n608 , n22065 );
xor ( n23078 , n23076 , n23077 );
and ( n23079 , n611 , n20976 );
xor ( n23080 , n23078 , n23079 );
xor ( n23081 , n23074 , n23080 );
and ( n23082 , n632 , n20156 );
and ( n23083 , n671 , n19222 );
xor ( n23084 , n23082 , n23083 );
and ( n23085 , n715 , n18407 );
xor ( n23086 , n23084 , n23085 );
xor ( n23087 , n23081 , n23086 );
xor ( n23088 , n23070 , n23087 );
and ( n23089 , n22072 , n22073 );
and ( n23090 , n22073 , n22075 );
and ( n23091 , n22072 , n22075 );
or ( n23092 , n23089 , n23090 , n23091 );
and ( n23093 , n22054 , n22055 );
and ( n23094 , n22055 , n22057 );
and ( n23095 , n22054 , n22057 );
or ( n23096 , n23093 , n23094 , n23095 );
xor ( n23097 , n23092 , n23096 );
and ( n23098 , n783 , n17422 );
and ( n23099 , n856 , n16550 );
xor ( n23100 , n23098 , n23099 );
and ( n23101 , n925 , n15691 );
xor ( n23102 , n23100 , n23101 );
xor ( n23103 , n23097 , n23102 );
xor ( n23104 , n23088 , n23103 );
xor ( n23105 , n23066 , n23104 );
and ( n23106 , n22026 , n22031 );
and ( n23107 , n22031 , n22037 );
and ( n23108 , n22026 , n22037 );
or ( n23109 , n23106 , n23107 , n23108 );
and ( n23110 , n22048 , n22052 );
and ( n23111 , n22052 , n22058 );
and ( n23112 , n22048 , n22058 );
or ( n23113 , n23110 , n23111 , n23112 );
xor ( n23114 , n23109 , n23113 );
and ( n23115 , n22027 , n22028 );
and ( n23116 , n22028 , n22030 );
and ( n23117 , n22027 , n22030 );
or ( n23118 , n23115 , n23116 , n23117 );
and ( n23119 , n1383 , n12531 );
and ( n23120 , n1580 , n11718 );
xor ( n23121 , n23119 , n23120 );
and ( n23122 , n1694 , n10977 );
xor ( n23123 , n23121 , n23122 );
xor ( n23124 , n23118 , n23123 );
and ( n23125 , n1047 , n14838 );
and ( n23126 , n1164 , n14044 );
xor ( n23127 , n23125 , n23126 );
and ( n23128 , n1287 , n13256 );
xor ( n23129 , n23127 , n23128 );
xor ( n23130 , n23124 , n23129 );
xor ( n23131 , n23114 , n23130 );
xor ( n23132 , n23105 , n23131 );
xor ( n23133 , n23062 , n23132 );
and ( n23134 , n21974 , n21990 );
and ( n23135 , n21990 , n22006 );
and ( n23136 , n21974 , n22006 );
or ( n23137 , n23134 , n23135 , n23136 );
and ( n23138 , n22017 , n22021 );
and ( n23139 , n22021 , n22038 );
and ( n23140 , n22017 , n22038 );
or ( n23141 , n23138 , n23139 , n23140 );
xor ( n23142 , n23137 , n23141 );
and ( n23143 , n21995 , n21999 );
and ( n23144 , n21999 , n22005 );
and ( n23145 , n21995 , n22005 );
or ( n23146 , n23143 , n23144 , n23145 );
and ( n23147 , n22001 , n22002 );
and ( n23148 , n22002 , n22004 );
and ( n23149 , n22001 , n22004 );
or ( n23150 , n23147 , n23148 , n23149 );
and ( n23151 , n22033 , n22034 );
and ( n23152 , n22034 , n22036 );
and ( n23153 , n22033 , n22036 );
or ( n23154 , n23151 , n23152 , n23153 );
xor ( n23155 , n23150 , n23154 );
and ( n23156 , n1933 , n10239 );
and ( n23157 , n2120 , n9348 );
xor ( n23158 , n23156 , n23157 );
and ( n23159 , n2324 , n8669 );
xor ( n23160 , n23158 , n23159 );
xor ( n23161 , n23155 , n23160 );
xor ( n23162 , n23146 , n23161 );
and ( n23163 , n21979 , n21980 );
and ( n23164 , n21980 , n21982 );
and ( n23165 , n21979 , n21982 );
or ( n23166 , n23163 , n23164 , n23165 );
and ( n23167 , n2462 , n8243 );
and ( n23168 , n2779 , n7662 );
xor ( n23169 , n23167 , n23168 );
and ( n23170 , n3024 , n7310 );
xor ( n23171 , n23169 , n23170 );
xor ( n23172 , n23166 , n23171 );
and ( n23173 , n3182 , n6971 );
and ( n23174 , n3545 , n6504 );
xor ( n23175 , n23173 , n23174 );
and ( n23176 , n3801 , n6132 );
xor ( n23177 , n23175 , n23176 );
xor ( n23178 , n23172 , n23177 );
xor ( n23179 , n23162 , n23178 );
xor ( n23180 , n23142 , n23179 );
xor ( n23181 , n23133 , n23180 );
xor ( n23182 , n23058 , n23181 );
xor ( n23183 , n22975 , n23182 );
xor ( n23184 , n22855 , n23183 );
and ( n23185 , n22086 , n22090 );
and ( n23186 , n22090 , n22192 );
and ( n23187 , n22086 , n22192 );
or ( n23188 , n23185 , n23186 , n23187 );
and ( n23189 , n22200 , n22206 );
xor ( n23190 , n23188 , n23189 );
and ( n23191 , n22201 , n22205 );
and ( n23192 , n22178 , n22179 );
and ( n23193 , n22179 , n22189 );
and ( n23194 , n22178 , n22189 );
or ( n23195 , n23192 , n23193 , n23194 );
and ( n23196 , n22136 , n22173 );
and ( n23197 , n22173 , n22190 );
and ( n23198 , n22136 , n22190 );
or ( n23199 , n23196 , n23197 , n23198 );
xor ( n23200 , n23195 , n23199 );
xor ( n23201 , n23191 , n23200 );
xor ( n23202 , n23190 , n23201 );
xor ( n23203 , n23184 , n23202 );
xor ( n23204 , n22851 , n23203 );
and ( n23205 , n21861 , n21865 );
and ( n23206 , n21865 , n22209 );
and ( n23207 , n21861 , n22209 );
or ( n23208 , n23205 , n23206 , n23207 );
xor ( n23209 , n23204 , n23208 );
and ( n23210 , n22210 , n22214 );
and ( n23211 , n22215 , n22218 );
or ( n23212 , n23210 , n23211 );
xor ( n23213 , n23209 , n23212 );
buf ( n23214 , n23213 );
buf ( n23215 , n23214 );
not ( n23216 , n23215 );
nor ( n23217 , n23216 , n8739 );
xor ( n23218 , n22845 , n23217 );
and ( n23219 , n21860 , n22223 );
and ( n23220 , n22224 , n22227 );
or ( n23221 , n23219 , n23220 );
xor ( n23222 , n23218 , n23221 );
buf ( n23223 , n23222 );
buf ( n23224 , n23223 );
not ( n23225 , n23224 );
buf ( n23226 , n552 );
not ( n23227 , n23226 );
nor ( n23228 , n23225 , n23227 );
xor ( n23229 , n22539 , n23228 );
xor ( n23230 , n22239 , n22536 );
nor ( n23231 , n22231 , n23227 );
and ( n23232 , n23230 , n23231 );
xor ( n23233 , n23230 , n23231 );
xor ( n23234 , n22243 , n22534 );
nor ( n23235 , n21258 , n23227 );
and ( n23236 , n23234 , n23235 );
xor ( n23237 , n23234 , n23235 );
xor ( n23238 , n22247 , n22532 );
nor ( n23239 , n20303 , n23227 );
and ( n23240 , n23238 , n23239 );
xor ( n23241 , n23238 , n23239 );
xor ( n23242 , n22251 , n22530 );
nor ( n23243 , n19365 , n23227 );
and ( n23244 , n23242 , n23243 );
xor ( n23245 , n23242 , n23243 );
xor ( n23246 , n22255 , n22528 );
nor ( n23247 , n18448 , n23227 );
and ( n23248 , n23246 , n23247 );
xor ( n23249 , n23246 , n23247 );
xor ( n23250 , n22259 , n22526 );
nor ( n23251 , n17548 , n23227 );
and ( n23252 , n23250 , n23251 );
xor ( n23253 , n23250 , n23251 );
xor ( n23254 , n22263 , n22524 );
nor ( n23255 , n16669 , n23227 );
and ( n23256 , n23254 , n23255 );
xor ( n23257 , n23254 , n23255 );
xor ( n23258 , n22267 , n22522 );
nor ( n23259 , n15809 , n23227 );
and ( n23260 , n23258 , n23259 );
xor ( n23261 , n23258 , n23259 );
xor ( n23262 , n22271 , n22520 );
nor ( n23263 , n14968 , n23227 );
and ( n23264 , n23262 , n23263 );
xor ( n23265 , n23262 , n23263 );
xor ( n23266 , n22275 , n22518 );
nor ( n23267 , n14147 , n23227 );
and ( n23268 , n23266 , n23267 );
xor ( n23269 , n23266 , n23267 );
xor ( n23270 , n22279 , n22516 );
nor ( n23271 , n13349 , n23227 );
and ( n23272 , n23270 , n23271 );
xor ( n23273 , n23270 , n23271 );
xor ( n23274 , n22283 , n22514 );
nor ( n23275 , n12564 , n23227 );
and ( n23276 , n23274 , n23275 );
xor ( n23277 , n23274 , n23275 );
xor ( n23278 , n22287 , n22512 );
nor ( n23279 , n11799 , n23227 );
and ( n23280 , n23278 , n23279 );
xor ( n23281 , n23278 , n23279 );
xor ( n23282 , n22291 , n22510 );
nor ( n23283 , n11050 , n23227 );
and ( n23284 , n23282 , n23283 );
xor ( n23285 , n23282 , n23283 );
xor ( n23286 , n22295 , n22508 );
nor ( n23287 , n10321 , n23227 );
and ( n23288 , n23286 , n23287 );
xor ( n23289 , n23286 , n23287 );
xor ( n23290 , n22299 , n22506 );
nor ( n23291 , n9429 , n23227 );
and ( n23292 , n23290 , n23291 );
xor ( n23293 , n23290 , n23291 );
xor ( n23294 , n22303 , n22504 );
nor ( n23295 , n8949 , n23227 );
and ( n23296 , n23294 , n23295 );
xor ( n23297 , n23294 , n23295 );
xor ( n23298 , n22307 , n22502 );
nor ( n23299 , n9437 , n23227 );
and ( n23300 , n23298 , n23299 );
xor ( n23301 , n23298 , n23299 );
xor ( n23302 , n22311 , n22500 );
nor ( n23303 , n9446 , n23227 );
and ( n23304 , n23302 , n23303 );
xor ( n23305 , n23302 , n23303 );
xor ( n23306 , n22315 , n22498 );
nor ( n23307 , n9455 , n23227 );
and ( n23308 , n23306 , n23307 );
xor ( n23309 , n23306 , n23307 );
xor ( n23310 , n22319 , n22496 );
nor ( n23311 , n9464 , n23227 );
and ( n23312 , n23310 , n23311 );
xor ( n23313 , n23310 , n23311 );
xor ( n23314 , n22323 , n22494 );
nor ( n23315 , n9473 , n23227 );
and ( n23316 , n23314 , n23315 );
xor ( n23317 , n23314 , n23315 );
xor ( n23318 , n22327 , n22492 );
nor ( n23319 , n9482 , n23227 );
and ( n23320 , n23318 , n23319 );
xor ( n23321 , n23318 , n23319 );
xor ( n23322 , n22331 , n22490 );
nor ( n23323 , n9491 , n23227 );
and ( n23324 , n23322 , n23323 );
xor ( n23325 , n23322 , n23323 );
xor ( n23326 , n22335 , n22488 );
nor ( n23327 , n9500 , n23227 );
and ( n23328 , n23326 , n23327 );
xor ( n23329 , n23326 , n23327 );
xor ( n23330 , n22339 , n22486 );
nor ( n23331 , n9509 , n23227 );
and ( n23332 , n23330 , n23331 );
xor ( n23333 , n23330 , n23331 );
xor ( n23334 , n22343 , n22484 );
nor ( n23335 , n9518 , n23227 );
and ( n23336 , n23334 , n23335 );
xor ( n23337 , n23334 , n23335 );
xor ( n23338 , n22347 , n22482 );
nor ( n23339 , n9527 , n23227 );
and ( n23340 , n23338 , n23339 );
xor ( n23341 , n23338 , n23339 );
xor ( n23342 , n22351 , n22480 );
nor ( n23343 , n9536 , n23227 );
and ( n23344 , n23342 , n23343 );
xor ( n23345 , n23342 , n23343 );
xor ( n23346 , n22355 , n22478 );
nor ( n23347 , n9545 , n23227 );
and ( n23348 , n23346 , n23347 );
xor ( n23349 , n23346 , n23347 );
xor ( n23350 , n22359 , n22476 );
nor ( n23351 , n9554 , n23227 );
and ( n23352 , n23350 , n23351 );
xor ( n23353 , n23350 , n23351 );
xor ( n23354 , n22363 , n22474 );
nor ( n23355 , n9563 , n23227 );
and ( n23356 , n23354 , n23355 );
xor ( n23357 , n23354 , n23355 );
xor ( n23358 , n22367 , n22472 );
nor ( n23359 , n9572 , n23227 );
and ( n23360 , n23358 , n23359 );
xor ( n23361 , n23358 , n23359 );
xor ( n23362 , n22371 , n22470 );
nor ( n23363 , n9581 , n23227 );
and ( n23364 , n23362 , n23363 );
xor ( n23365 , n23362 , n23363 );
xor ( n23366 , n22375 , n22468 );
nor ( n23367 , n9590 , n23227 );
and ( n23368 , n23366 , n23367 );
xor ( n23369 , n23366 , n23367 );
xor ( n23370 , n22379 , n22466 );
nor ( n23371 , n9599 , n23227 );
and ( n23372 , n23370 , n23371 );
xor ( n23373 , n23370 , n23371 );
xor ( n23374 , n22383 , n22464 );
nor ( n23375 , n9608 , n23227 );
and ( n23376 , n23374 , n23375 );
xor ( n23377 , n23374 , n23375 );
xor ( n23378 , n22387 , n22462 );
nor ( n23379 , n9617 , n23227 );
and ( n23380 , n23378 , n23379 );
xor ( n23381 , n23378 , n23379 );
xor ( n23382 , n22391 , n22460 );
nor ( n23383 , n9626 , n23227 );
and ( n23384 , n23382 , n23383 );
xor ( n23385 , n23382 , n23383 );
xor ( n23386 , n22395 , n22458 );
nor ( n23387 , n9635 , n23227 );
and ( n23388 , n23386 , n23387 );
xor ( n23389 , n23386 , n23387 );
xor ( n23390 , n22399 , n22456 );
nor ( n23391 , n9644 , n23227 );
and ( n23392 , n23390 , n23391 );
xor ( n23393 , n23390 , n23391 );
xor ( n23394 , n22403 , n22454 );
nor ( n23395 , n9653 , n23227 );
and ( n23396 , n23394 , n23395 );
xor ( n23397 , n23394 , n23395 );
xor ( n23398 , n22407 , n22452 );
nor ( n23399 , n9662 , n23227 );
and ( n23400 , n23398 , n23399 );
xor ( n23401 , n23398 , n23399 );
xor ( n23402 , n22411 , n22450 );
nor ( n23403 , n9671 , n23227 );
and ( n23404 , n23402 , n23403 );
xor ( n23405 , n23402 , n23403 );
xor ( n23406 , n22415 , n22448 );
nor ( n23407 , n9680 , n23227 );
and ( n23408 , n23406 , n23407 );
xor ( n23409 , n23406 , n23407 );
xor ( n23410 , n22419 , n22446 );
nor ( n23411 , n9689 , n23227 );
and ( n23412 , n23410 , n23411 );
xor ( n23413 , n23410 , n23411 );
xor ( n23414 , n22423 , n22444 );
nor ( n23415 , n9698 , n23227 );
and ( n23416 , n23414 , n23415 );
xor ( n23417 , n23414 , n23415 );
xor ( n23418 , n22427 , n22442 );
nor ( n23419 , n9707 , n23227 );
and ( n23420 , n23418 , n23419 );
xor ( n23421 , n23418 , n23419 );
xor ( n23422 , n22431 , n22440 );
nor ( n23423 , n9716 , n23227 );
and ( n23424 , n23422 , n23423 );
xor ( n23425 , n23422 , n23423 );
xor ( n23426 , n22435 , n22438 );
nor ( n23427 , n9725 , n23227 );
and ( n23428 , n23426 , n23427 );
xor ( n23429 , n23426 , n23427 );
xor ( n23430 , n22436 , n22437 );
nor ( n23431 , n9734 , n23227 );
and ( n23432 , n23430 , n23431 );
xor ( n23433 , n23430 , n23431 );
nor ( n23434 , n9752 , n22233 );
nor ( n23435 , n9743 , n23227 );
and ( n23436 , n23434 , n23435 );
and ( n23437 , n23433 , n23436 );
or ( n23438 , n23432 , n23437 );
and ( n23439 , n23429 , n23438 );
or ( n23440 , n23428 , n23439 );
and ( n23441 , n23425 , n23440 );
or ( n23442 , n23424 , n23441 );
and ( n23443 , n23421 , n23442 );
or ( n23444 , n23420 , n23443 );
and ( n23445 , n23417 , n23444 );
or ( n23446 , n23416 , n23445 );
and ( n23447 , n23413 , n23446 );
or ( n23448 , n23412 , n23447 );
and ( n23449 , n23409 , n23448 );
or ( n23450 , n23408 , n23449 );
and ( n23451 , n23405 , n23450 );
or ( n23452 , n23404 , n23451 );
and ( n23453 , n23401 , n23452 );
or ( n23454 , n23400 , n23453 );
and ( n23455 , n23397 , n23454 );
or ( n23456 , n23396 , n23455 );
and ( n23457 , n23393 , n23456 );
or ( n23458 , n23392 , n23457 );
and ( n23459 , n23389 , n23458 );
or ( n23460 , n23388 , n23459 );
and ( n23461 , n23385 , n23460 );
or ( n23462 , n23384 , n23461 );
and ( n23463 , n23381 , n23462 );
or ( n23464 , n23380 , n23463 );
and ( n23465 , n23377 , n23464 );
or ( n23466 , n23376 , n23465 );
and ( n23467 , n23373 , n23466 );
or ( n23468 , n23372 , n23467 );
and ( n23469 , n23369 , n23468 );
or ( n23470 , n23368 , n23469 );
and ( n23471 , n23365 , n23470 );
or ( n23472 , n23364 , n23471 );
and ( n23473 , n23361 , n23472 );
or ( n23474 , n23360 , n23473 );
and ( n23475 , n23357 , n23474 );
or ( n23476 , n23356 , n23475 );
and ( n23477 , n23353 , n23476 );
or ( n23478 , n23352 , n23477 );
and ( n23479 , n23349 , n23478 );
or ( n23480 , n23348 , n23479 );
and ( n23481 , n23345 , n23480 );
or ( n23482 , n23344 , n23481 );
and ( n23483 , n23341 , n23482 );
or ( n23484 , n23340 , n23483 );
and ( n23485 , n23337 , n23484 );
or ( n23486 , n23336 , n23485 );
and ( n23487 , n23333 , n23486 );
or ( n23488 , n23332 , n23487 );
and ( n23489 , n23329 , n23488 );
or ( n23490 , n23328 , n23489 );
and ( n23491 , n23325 , n23490 );
or ( n23492 , n23324 , n23491 );
and ( n23493 , n23321 , n23492 );
or ( n23494 , n23320 , n23493 );
and ( n23495 , n23317 , n23494 );
or ( n23496 , n23316 , n23495 );
and ( n23497 , n23313 , n23496 );
or ( n23498 , n23312 , n23497 );
and ( n23499 , n23309 , n23498 );
or ( n23500 , n23308 , n23499 );
and ( n23501 , n23305 , n23500 );
or ( n23502 , n23304 , n23501 );
and ( n23503 , n23301 , n23502 );
or ( n23504 , n23300 , n23503 );
and ( n23505 , n23297 , n23504 );
or ( n23506 , n23296 , n23505 );
and ( n23507 , n23293 , n23506 );
or ( n23508 , n23292 , n23507 );
and ( n23509 , n23289 , n23508 );
or ( n23510 , n23288 , n23509 );
and ( n23511 , n23285 , n23510 );
or ( n23512 , n23284 , n23511 );
and ( n23513 , n23281 , n23512 );
or ( n23514 , n23280 , n23513 );
and ( n23515 , n23277 , n23514 );
or ( n23516 , n23276 , n23515 );
and ( n23517 , n23273 , n23516 );
or ( n23518 , n23272 , n23517 );
and ( n23519 , n23269 , n23518 );
or ( n23520 , n23268 , n23519 );
and ( n23521 , n23265 , n23520 );
or ( n23522 , n23264 , n23521 );
and ( n23523 , n23261 , n23522 );
or ( n23524 , n23260 , n23523 );
and ( n23525 , n23257 , n23524 );
or ( n23526 , n23256 , n23525 );
and ( n23527 , n23253 , n23526 );
or ( n23528 , n23252 , n23527 );
and ( n23529 , n23249 , n23528 );
or ( n23530 , n23248 , n23529 );
and ( n23531 , n23245 , n23530 );
or ( n23532 , n23244 , n23531 );
and ( n23533 , n23241 , n23532 );
or ( n23534 , n23240 , n23533 );
and ( n23535 , n23237 , n23534 );
or ( n23536 , n23236 , n23535 );
and ( n23537 , n23233 , n23536 );
or ( n23538 , n23232 , n23537 );
xor ( n23539 , n23229 , n23538 );
buf ( n23540 , n480 );
not ( n23541 , n23540 );
nor ( n23542 , n601 , n23541 );
buf ( n23543 , n23542 );
nor ( n23544 , n622 , n21562 );
xor ( n23545 , n23543 , n23544 );
buf ( n23546 , n23545 );
nor ( n23547 , n646 , n20601 );
xor ( n23548 , n23546 , n23547 );
and ( n23549 , n22543 , n22544 );
buf ( n23550 , n23549 );
xor ( n23551 , n23548 , n23550 );
nor ( n23552 , n684 , n19657 );
xor ( n23553 , n23551 , n23552 );
and ( n23554 , n22546 , n22547 );
and ( n23555 , n22548 , n22550 );
or ( n23556 , n23554 , n23555 );
xor ( n23557 , n23553 , n23556 );
nor ( n23558 , n733 , n18734 );
xor ( n23559 , n23557 , n23558 );
and ( n23560 , n22551 , n22552 );
and ( n23561 , n22553 , n22556 );
or ( n23562 , n23560 , n23561 );
xor ( n23563 , n23559 , n23562 );
nor ( n23564 , n796 , n17828 );
xor ( n23565 , n23563 , n23564 );
and ( n23566 , n22557 , n22558 );
and ( n23567 , n22559 , n22562 );
or ( n23568 , n23566 , n23567 );
xor ( n23569 , n23565 , n23568 );
nor ( n23570 , n868 , n16943 );
xor ( n23571 , n23569 , n23570 );
and ( n23572 , n22563 , n22564 );
and ( n23573 , n22565 , n22568 );
or ( n23574 , n23572 , n23573 );
xor ( n23575 , n23571 , n23574 );
nor ( n23576 , n958 , n16077 );
xor ( n23577 , n23575 , n23576 );
and ( n23578 , n22569 , n22570 );
and ( n23579 , n22571 , n22574 );
or ( n23580 , n23578 , n23579 );
xor ( n23581 , n23577 , n23580 );
nor ( n23582 , n1062 , n15230 );
xor ( n23583 , n23581 , n23582 );
and ( n23584 , n22575 , n22576 );
and ( n23585 , n22577 , n22580 );
or ( n23586 , n23584 , n23585 );
xor ( n23587 , n23583 , n23586 );
nor ( n23588 , n1176 , n14403 );
xor ( n23589 , n23587 , n23588 );
and ( n23590 , n22581 , n22582 );
and ( n23591 , n22583 , n22586 );
or ( n23592 , n23590 , n23591 );
xor ( n23593 , n23589 , n23592 );
nor ( n23594 , n1303 , n13599 );
xor ( n23595 , n23593 , n23594 );
and ( n23596 , n22587 , n22588 );
and ( n23597 , n22589 , n22592 );
or ( n23598 , n23596 , n23597 );
xor ( n23599 , n23595 , n23598 );
nor ( n23600 , n1445 , n12808 );
xor ( n23601 , n23599 , n23600 );
and ( n23602 , n22593 , n22594 );
and ( n23603 , n22595 , n22598 );
or ( n23604 , n23602 , n23603 );
xor ( n23605 , n23601 , n23604 );
nor ( n23606 , n1598 , n12037 );
xor ( n23607 , n23605 , n23606 );
and ( n23608 , n22599 , n22600 );
and ( n23609 , n22601 , n22604 );
or ( n23610 , n23608 , n23609 );
xor ( n23611 , n23607 , n23610 );
nor ( n23612 , n1766 , n11282 );
xor ( n23613 , n23611 , n23612 );
and ( n23614 , n22605 , n22606 );
and ( n23615 , n22607 , n22610 );
or ( n23616 , n23614 , n23615 );
xor ( n23617 , n23613 , n23616 );
nor ( n23618 , n1945 , n10547 );
xor ( n23619 , n23617 , n23618 );
and ( n23620 , n22611 , n22612 );
and ( n23621 , n22613 , n22616 );
or ( n23622 , n23620 , n23621 );
xor ( n23623 , n23619 , n23622 );
nor ( n23624 , n2137 , n9829 );
xor ( n23625 , n23623 , n23624 );
and ( n23626 , n22617 , n22618 );
and ( n23627 , n22619 , n22622 );
or ( n23628 , n23626 , n23627 );
xor ( n23629 , n23625 , n23628 );
nor ( n23630 , n2343 , n8955 );
xor ( n23631 , n23629 , n23630 );
and ( n23632 , n22623 , n22624 );
and ( n23633 , n22625 , n22628 );
or ( n23634 , n23632 , n23633 );
xor ( n23635 , n23631 , n23634 );
nor ( n23636 , n2566 , n603 );
xor ( n23637 , n23635 , n23636 );
and ( n23638 , n22629 , n22630 );
and ( n23639 , n22631 , n22634 );
or ( n23640 , n23638 , n23639 );
xor ( n23641 , n23637 , n23640 );
nor ( n23642 , n2797 , n652 );
xor ( n23643 , n23641 , n23642 );
and ( n23644 , n22635 , n22636 );
and ( n23645 , n22637 , n22640 );
or ( n23646 , n23644 , n23645 );
xor ( n23647 , n23643 , n23646 );
nor ( n23648 , n3043 , n624 );
xor ( n23649 , n23647 , n23648 );
and ( n23650 , n22641 , n22642 );
and ( n23651 , n22643 , n22646 );
or ( n23652 , n23650 , n23651 );
xor ( n23653 , n23649 , n23652 );
nor ( n23654 , n3300 , n648 );
xor ( n23655 , n23653 , n23654 );
and ( n23656 , n22647 , n22648 );
and ( n23657 , n22649 , n22652 );
or ( n23658 , n23656 , n23657 );
xor ( n23659 , n23655 , n23658 );
nor ( n23660 , n3570 , n686 );
xor ( n23661 , n23659 , n23660 );
and ( n23662 , n22653 , n22654 );
and ( n23663 , n22655 , n22658 );
or ( n23664 , n23662 , n23663 );
xor ( n23665 , n23661 , n23664 );
nor ( n23666 , n3853 , n735 );
xor ( n23667 , n23665 , n23666 );
and ( n23668 , n22659 , n22660 );
and ( n23669 , n22661 , n22664 );
or ( n23670 , n23668 , n23669 );
xor ( n23671 , n23667 , n23670 );
nor ( n23672 , n4151 , n798 );
xor ( n23673 , n23671 , n23672 );
and ( n23674 , n22665 , n22666 );
and ( n23675 , n22667 , n22670 );
or ( n23676 , n23674 , n23675 );
xor ( n23677 , n23673 , n23676 );
nor ( n23678 , n4458 , n870 );
xor ( n23679 , n23677 , n23678 );
and ( n23680 , n22671 , n22672 );
and ( n23681 , n22673 , n22676 );
or ( n23682 , n23680 , n23681 );
xor ( n23683 , n23679 , n23682 );
nor ( n23684 , n4786 , n960 );
xor ( n23685 , n23683 , n23684 );
and ( n23686 , n22677 , n22678 );
and ( n23687 , n22679 , n22682 );
or ( n23688 , n23686 , n23687 );
xor ( n23689 , n23685 , n23688 );
nor ( n23690 , n5126 , n1064 );
xor ( n23691 , n23689 , n23690 );
and ( n23692 , n22683 , n22684 );
and ( n23693 , n22685 , n22688 );
or ( n23694 , n23692 , n23693 );
xor ( n23695 , n23691 , n23694 );
nor ( n23696 , n5477 , n1178 );
xor ( n23697 , n23695 , n23696 );
and ( n23698 , n22689 , n22690 );
and ( n23699 , n22691 , n22694 );
or ( n23700 , n23698 , n23699 );
xor ( n23701 , n23697 , n23700 );
nor ( n23702 , n5838 , n1305 );
xor ( n23703 , n23701 , n23702 );
and ( n23704 , n22695 , n22696 );
and ( n23705 , n22697 , n22700 );
or ( n23706 , n23704 , n23705 );
xor ( n23707 , n23703 , n23706 );
nor ( n23708 , n6212 , n1447 );
xor ( n23709 , n23707 , n23708 );
and ( n23710 , n22701 , n22702 );
and ( n23711 , n22703 , n22706 );
or ( n23712 , n23710 , n23711 );
xor ( n23713 , n23709 , n23712 );
nor ( n23714 , n6596 , n1600 );
xor ( n23715 , n23713 , n23714 );
and ( n23716 , n22707 , n22708 );
and ( n23717 , n22709 , n22712 );
or ( n23718 , n23716 , n23717 );
xor ( n23719 , n23715 , n23718 );
nor ( n23720 , n6997 , n1768 );
xor ( n23721 , n23719 , n23720 );
and ( n23722 , n22713 , n22714 );
and ( n23723 , n22715 , n22718 );
or ( n23724 , n23722 , n23723 );
xor ( n23725 , n23721 , n23724 );
nor ( n23726 , n7413 , n1947 );
xor ( n23727 , n23725 , n23726 );
and ( n23728 , n22719 , n22720 );
and ( n23729 , n22721 , n22724 );
or ( n23730 , n23728 , n23729 );
xor ( n23731 , n23727 , n23730 );
nor ( n23732 , n7841 , n2139 );
xor ( n23733 , n23731 , n23732 );
and ( n23734 , n22725 , n22726 );
and ( n23735 , n22727 , n22730 );
or ( n23736 , n23734 , n23735 );
xor ( n23737 , n23733 , n23736 );
nor ( n23738 , n8281 , n2345 );
xor ( n23739 , n23737 , n23738 );
and ( n23740 , n22731 , n22732 );
and ( n23741 , n22733 , n22736 );
or ( n23742 , n23740 , n23741 );
xor ( n23743 , n23739 , n23742 );
nor ( n23744 , n8737 , n2568 );
xor ( n23745 , n23743 , n23744 );
and ( n23746 , n22737 , n22738 );
and ( n23747 , n22739 , n22742 );
or ( n23748 , n23746 , n23747 );
xor ( n23749 , n23745 , n23748 );
nor ( n23750 , n9420 , n2799 );
xor ( n23751 , n23749 , n23750 );
and ( n23752 , n22743 , n22744 );
and ( n23753 , n22745 , n22748 );
or ( n23754 , n23752 , n23753 );
xor ( n23755 , n23751 , n23754 );
nor ( n23756 , n10312 , n3045 );
xor ( n23757 , n23755 , n23756 );
and ( n23758 , n22749 , n22750 );
and ( n23759 , n22751 , n22754 );
or ( n23760 , n23758 , n23759 );
xor ( n23761 , n23757 , n23760 );
nor ( n23762 , n11041 , n3302 );
xor ( n23763 , n23761 , n23762 );
and ( n23764 , n22755 , n22756 );
and ( n23765 , n22757 , n22760 );
or ( n23766 , n23764 , n23765 );
xor ( n23767 , n23763 , n23766 );
nor ( n23768 , n11790 , n3572 );
xor ( n23769 , n23767 , n23768 );
and ( n23770 , n22761 , n22762 );
and ( n23771 , n22763 , n22766 );
or ( n23772 , n23770 , n23771 );
xor ( n23773 , n23769 , n23772 );
nor ( n23774 , n12555 , n3855 );
xor ( n23775 , n23773 , n23774 );
and ( n23776 , n22767 , n22768 );
and ( n23777 , n22769 , n22772 );
or ( n23778 , n23776 , n23777 );
xor ( n23779 , n23775 , n23778 );
nor ( n23780 , n13340 , n4153 );
xor ( n23781 , n23779 , n23780 );
and ( n23782 , n22773 , n22774 );
and ( n23783 , n22775 , n22778 );
or ( n23784 , n23782 , n23783 );
xor ( n23785 , n23781 , n23784 );
nor ( n23786 , n14138 , n4460 );
xor ( n23787 , n23785 , n23786 );
and ( n23788 , n22779 , n22780 );
and ( n23789 , n22781 , n22784 );
or ( n23790 , n23788 , n23789 );
xor ( n23791 , n23787 , n23790 );
nor ( n23792 , n14959 , n4788 );
xor ( n23793 , n23791 , n23792 );
and ( n23794 , n22785 , n22786 );
and ( n23795 , n22787 , n22790 );
or ( n23796 , n23794 , n23795 );
xor ( n23797 , n23793 , n23796 );
nor ( n23798 , n15800 , n5128 );
xor ( n23799 , n23797 , n23798 );
and ( n23800 , n22791 , n22792 );
and ( n23801 , n22793 , n22796 );
or ( n23802 , n23800 , n23801 );
xor ( n23803 , n23799 , n23802 );
nor ( n23804 , n16660 , n5479 );
xor ( n23805 , n23803 , n23804 );
and ( n23806 , n22797 , n22798 );
and ( n23807 , n22799 , n22802 );
or ( n23808 , n23806 , n23807 );
xor ( n23809 , n23805 , n23808 );
nor ( n23810 , n17539 , n5840 );
xor ( n23811 , n23809 , n23810 );
and ( n23812 , n22803 , n22804 );
and ( n23813 , n22805 , n22808 );
or ( n23814 , n23812 , n23813 );
xor ( n23815 , n23811 , n23814 );
nor ( n23816 , n18439 , n6214 );
xor ( n23817 , n23815 , n23816 );
and ( n23818 , n22809 , n22810 );
and ( n23819 , n22811 , n22814 );
or ( n23820 , n23818 , n23819 );
xor ( n23821 , n23817 , n23820 );
nor ( n23822 , n19356 , n6598 );
xor ( n23823 , n23821 , n23822 );
and ( n23824 , n22815 , n22816 );
and ( n23825 , n22817 , n22820 );
or ( n23826 , n23824 , n23825 );
xor ( n23827 , n23823 , n23826 );
nor ( n23828 , n20294 , n6999 );
xor ( n23829 , n23827 , n23828 );
and ( n23830 , n22821 , n22822 );
and ( n23831 , n22823 , n22826 );
or ( n23832 , n23830 , n23831 );
xor ( n23833 , n23829 , n23832 );
nor ( n23834 , n21249 , n7415 );
xor ( n23835 , n23833 , n23834 );
and ( n23836 , n22827 , n22828 );
and ( n23837 , n22829 , n22832 );
or ( n23838 , n23836 , n23837 );
xor ( n23839 , n23835 , n23838 );
nor ( n23840 , n22222 , n7843 );
xor ( n23841 , n23839 , n23840 );
and ( n23842 , n22833 , n22834 );
and ( n23843 , n22835 , n22838 );
or ( n23844 , n23842 , n23843 );
xor ( n23845 , n23841 , n23844 );
nor ( n23846 , n23216 , n8283 );
xor ( n23847 , n23845 , n23846 );
and ( n23848 , n22839 , n22840 );
and ( n23849 , n22841 , n22844 );
or ( n23850 , n23848 , n23849 );
xor ( n23851 , n23847 , n23850 );
and ( n23852 , n23188 , n23189 );
and ( n23853 , n23189 , n23201 );
and ( n23854 , n23188 , n23201 );
or ( n23855 , n23852 , n23853 , n23854 );
and ( n23856 , n22855 , n23183 );
and ( n23857 , n23183 , n23202 );
and ( n23858 , n22855 , n23202 );
or ( n23859 , n23856 , n23857 , n23858 );
xor ( n23860 , n23855 , n23859 );
and ( n23861 , n22859 , n22974 );
and ( n23862 , n22974 , n23182 );
and ( n23863 , n22859 , n23182 );
or ( n23864 , n23861 , n23862 , n23863 );
and ( n23865 , n22979 , n23057 );
and ( n23866 , n23057 , n23181 );
and ( n23867 , n22979 , n23181 );
or ( n23868 , n23865 , n23866 , n23867 );
and ( n23869 , n22983 , n22987 );
and ( n23870 , n22987 , n23056 );
and ( n23871 , n22983 , n23056 );
or ( n23872 , n23869 , n23870 , n23871 );
and ( n23873 , n22872 , n22935 );
and ( n23874 , n22935 , n22972 );
and ( n23875 , n22872 , n22972 );
or ( n23876 , n23873 , n23874 , n23875 );
xor ( n23877 , n23872 , n23876 );
and ( n23878 , n22940 , n22944 );
and ( n23879 , n22944 , n22971 );
and ( n23880 , n22940 , n22971 );
or ( n23881 , n23878 , n23879 , n23880 );
and ( n23882 , n22901 , n22917 );
and ( n23883 , n22917 , n22933 );
and ( n23884 , n22901 , n22933 );
or ( n23885 , n23882 , n23883 , n23884 );
and ( n23886 , n22886 , n22887 );
and ( n23887 , n22887 , n22894 );
and ( n23888 , n22886 , n22894 );
or ( n23889 , n23886 , n23887 , n23888 );
and ( n23890 , n22905 , n22910 );
and ( n23891 , n22910 , n22916 );
and ( n23892 , n22905 , n22916 );
or ( n23893 , n23890 , n23891 , n23892 );
xor ( n23894 , n23889 , n23893 );
and ( n23895 , n22889 , n22890 );
and ( n23896 , n22890 , n22893 );
and ( n23897 , n22889 , n22893 );
or ( n23898 , n23895 , n23896 , n23897 );
and ( n23899 , n22906 , n22907 );
and ( n23900 , n22907 , n22909 );
and ( n23901 , n22906 , n22909 );
or ( n23902 , n23899 , n23900 , n23901 );
xor ( n23903 , n23898 , n23902 );
and ( n23904 , n21216 , n635 );
and ( n23905 , n22186 , n606 );
xor ( n23906 , n23904 , n23905 );
and ( n23907 , n22892 , n615 );
xor ( n23908 , n23906 , n23907 );
xor ( n23909 , n23903 , n23908 );
xor ( n23910 , n23894 , n23909 );
xor ( n23911 , n23885 , n23910 );
and ( n23912 , n22922 , n22926 );
and ( n23913 , n22926 , n22932 );
and ( n23914 , n22922 , n22932 );
or ( n23915 , n23912 , n23913 , n23914 );
and ( n23916 , n22912 , n22913 );
and ( n23917 , n22913 , n22915 );
and ( n23918 , n22912 , n22915 );
or ( n23919 , n23916 , n23917 , n23918 );
and ( n23920 , n18144 , n771 );
and ( n23921 , n19324 , n719 );
xor ( n23922 , n23920 , n23921 );
and ( n23923 , n20233 , n663 );
xor ( n23924 , n23922 , n23923 );
xor ( n23925 , n23919 , n23924 );
and ( n23926 , n15758 , n1034 );
and ( n23927 , n16637 , n940 );
xor ( n23928 , n23926 , n23927 );
and ( n23929 , n17512 , n840 );
xor ( n23930 , n23928 , n23929 );
xor ( n23931 , n23925 , n23930 );
xor ( n23932 , n23915 , n23931 );
and ( n23933 , n22928 , n22929 );
and ( n23934 , n22929 , n22931 );
and ( n23935 , n22928 , n22931 );
or ( n23936 , n23933 , n23934 , n23935 );
and ( n23937 , n22959 , n22960 );
and ( n23938 , n22960 , n22962 );
and ( n23939 , n22959 , n22962 );
or ( n23940 , n23937 , n23938 , n23939 );
xor ( n23941 , n23936 , n23940 );
and ( n23942 , n13322 , n1424 );
and ( n23943 , n14118 , n1254 );
xor ( n23944 , n23942 , n23943 );
and ( n23945 , n14938 , n1134 );
xor ( n23946 , n23944 , n23945 );
xor ( n23947 , n23941 , n23946 );
xor ( n23948 , n23932 , n23947 );
xor ( n23949 , n23911 , n23948 );
xor ( n23950 , n23881 , n23949 );
and ( n23951 , n22949 , n22953 );
and ( n23952 , n22953 , n22970 );
and ( n23953 , n22949 , n22970 );
or ( n23954 , n23951 , n23952 , n23953 );
and ( n23955 , n23022 , n23037 );
and ( n23956 , n23037 , n23054 );
and ( n23957 , n23022 , n23054 );
or ( n23958 , n23955 , n23956 , n23957 );
xor ( n23959 , n23954 , n23958 );
and ( n23960 , n22958 , n22963 );
and ( n23961 , n22963 , n22969 );
and ( n23962 , n22958 , n22969 );
or ( n23963 , n23960 , n23961 , n23962 );
and ( n23964 , n23026 , n23030 );
and ( n23965 , n23030 , n23036 );
and ( n23966 , n23026 , n23036 );
or ( n23967 , n23964 , n23965 , n23966 );
xor ( n23968 , n23963 , n23967 );
and ( n23969 , n22965 , n22966 );
and ( n23970 , n22966 , n22968 );
and ( n23971 , n22965 , n22968 );
or ( n23972 , n23969 , n23970 , n23971 );
and ( n23973 , n11015 , n1882 );
and ( n23974 , n11769 , n1738 );
xor ( n23975 , n23973 , n23974 );
and ( n23976 , n12320 , n1551 );
xor ( n23977 , n23975 , n23976 );
xor ( n23978 , n23972 , n23977 );
and ( n23979 , n8718 , n2544 );
and ( n23980 , n9400 , n2298 );
xor ( n23981 , n23979 , n23980 );
and ( n23982 , n10291 , n2100 );
xor ( n23983 , n23981 , n23982 );
xor ( n23984 , n23978 , n23983 );
xor ( n23985 , n23968 , n23984 );
xor ( n23986 , n23959 , n23985 );
xor ( n23987 , n23950 , n23986 );
xor ( n23988 , n23877 , n23987 );
xor ( n23989 , n23868 , n23988 );
and ( n23990 , n23062 , n23132 );
and ( n23991 , n23132 , n23180 );
and ( n23992 , n23062 , n23180 );
or ( n23993 , n23990 , n23991 , n23992 );
and ( n23994 , n22992 , n23017 );
and ( n23995 , n23017 , n23055 );
and ( n23996 , n22992 , n23055 );
or ( n23997 , n23994 , n23995 , n23996 );
and ( n23998 , n23137 , n23141 );
and ( n23999 , n23141 , n23179 );
and ( n24000 , n23137 , n23179 );
or ( n24001 , n23998 , n23999 , n24000 );
xor ( n24002 , n23997 , n24001 );
and ( n24003 , n22996 , n23000 );
and ( n24004 , n23000 , n23016 );
and ( n24005 , n22996 , n23016 );
or ( n24006 , n24003 , n24004 , n24005 );
and ( n24007 , n23005 , n23009 );
and ( n24008 , n23009 , n23015 );
and ( n24009 , n23005 , n23015 );
or ( n24010 , n24007 , n24008 , n24009 );
and ( n24011 , n23166 , n23171 );
and ( n24012 , n23171 , n23177 );
and ( n24013 , n23166 , n23177 );
or ( n24014 , n24011 , n24012 , n24013 );
xor ( n24015 , n24010 , n24014 );
and ( n24016 , n23011 , n23012 );
and ( n24017 , n23012 , n23014 );
and ( n24018 , n23011 , n23014 );
or ( n24019 , n24016 , n24017 , n24018 );
and ( n24020 , n23173 , n23174 );
and ( n24021 , n23174 , n23176 );
and ( n24022 , n23173 , n23176 );
or ( n24023 , n24020 , n24021 , n24022 );
xor ( n24024 , n24019 , n24023 );
and ( n24025 , n4132 , n6132 );
and ( n24026 , n4438 , n5765 );
xor ( n24027 , n24025 , n24026 );
and ( n24028 , n4766 , n5408 );
xor ( n24029 , n24027 , n24028 );
xor ( n24030 , n24024 , n24029 );
xor ( n24031 , n24015 , n24030 );
xor ( n24032 , n24006 , n24031 );
and ( n24033 , n23042 , n23047 );
and ( n24034 , n23047 , n23053 );
and ( n24035 , n23042 , n23053 );
or ( n24036 , n24033 , n24034 , n24035 );
and ( n24037 , n23032 , n23033 );
and ( n24038 , n23033 , n23035 );
and ( n24039 , n23032 , n23035 );
or ( n24040 , n24037 , n24038 , n24039 );
and ( n24041 , n23043 , n23044 );
and ( n24042 , n23044 , n23046 );
and ( n24043 , n23043 , n23046 );
or ( n24044 , n24041 , n24042 , n24043 );
xor ( n24045 , n24040 , n24044 );
and ( n24046 , n7385 , n3271 );
and ( n24047 , n7808 , n2981 );
xor ( n24048 , n24046 , n24047 );
and ( n24049 , n8079 , n2739 );
xor ( n24050 , n24048 , n24049 );
xor ( n24051 , n24045 , n24050 );
xor ( n24052 , n24036 , n24051 );
and ( n24053 , n23049 , n23050 );
and ( n24054 , n23050 , n23052 );
and ( n24055 , n23049 , n23052 );
or ( n24056 , n24053 , n24054 , n24055 );
and ( n24057 , n6187 , n4102 );
and ( n24058 , n6569 , n3749 );
xor ( n24059 , n24057 , n24058 );
and ( n24060 , n6816 , n3495 );
xor ( n24061 , n24059 , n24060 );
xor ( n24062 , n24056 , n24061 );
buf ( n24063 , n4959 );
and ( n24064 , n5459 , n4730 );
xor ( n24065 , n24063 , n24064 );
and ( n24066 , n5819 , n4403 );
xor ( n24067 , n24065 , n24066 );
xor ( n24068 , n24062 , n24067 );
xor ( n24069 , n24052 , n24068 );
xor ( n24070 , n24032 , n24069 );
xor ( n24071 , n24002 , n24070 );
xor ( n24072 , n23993 , n24071 );
and ( n24073 , n23066 , n23104 );
and ( n24074 , n23104 , n23131 );
and ( n24075 , n23066 , n23131 );
or ( n24076 , n24073 , n24074 , n24075 );
and ( n24077 , n23109 , n23113 );
and ( n24078 , n23113 , n23130 );
and ( n24079 , n23109 , n23130 );
or ( n24080 , n24077 , n24078 , n24079 );
and ( n24081 , n23146 , n23161 );
and ( n24082 , n23161 , n23178 );
and ( n24083 , n23146 , n23178 );
or ( n24084 , n24081 , n24082 , n24083 );
xor ( n24085 , n24080 , n24084 );
and ( n24086 , n23150 , n23154 );
and ( n24087 , n23154 , n23160 );
and ( n24088 , n23150 , n23160 );
or ( n24089 , n24086 , n24087 , n24088 );
and ( n24090 , n23156 , n23157 );
and ( n24091 , n23157 , n23159 );
and ( n24092 , n23156 , n23159 );
or ( n24093 , n24090 , n24091 , n24092 );
and ( n24094 , n23119 , n23120 );
and ( n24095 , n23120 , n23122 );
and ( n24096 , n23119 , n23122 );
or ( n24097 , n24094 , n24095 , n24096 );
xor ( n24098 , n24093 , n24097 );
and ( n24099 , n1933 , n10977 );
and ( n24100 , n2120 , n10239 );
xor ( n24101 , n24099 , n24100 );
and ( n24102 , n2324 , n9348 );
xor ( n24103 , n24101 , n24102 );
xor ( n24104 , n24098 , n24103 );
xor ( n24105 , n24089 , n24104 );
and ( n24106 , n23167 , n23168 );
and ( n24107 , n23168 , n23170 );
and ( n24108 , n23167 , n23170 );
or ( n24109 , n24106 , n24107 , n24108 );
and ( n24110 , n2462 , n8669 );
and ( n24111 , n2779 , n8243 );
xor ( n24112 , n24110 , n24111 );
and ( n24113 , n3024 , n7662 );
xor ( n24114 , n24112 , n24113 );
xor ( n24115 , n24109 , n24114 );
and ( n24116 , n3182 , n7310 );
and ( n24117 , n3545 , n6971 );
xor ( n24118 , n24116 , n24117 );
and ( n24119 , n3801 , n6504 );
xor ( n24120 , n24118 , n24119 );
xor ( n24121 , n24115 , n24120 );
xor ( n24122 , n24105 , n24121 );
xor ( n24123 , n24085 , n24122 );
xor ( n24124 , n24076 , n24123 );
and ( n24125 , n23070 , n23087 );
and ( n24126 , n23087 , n23103 );
and ( n24127 , n23070 , n23103 );
or ( n24128 , n24125 , n24126 , n24127 );
and ( n24129 , n23074 , n23080 );
and ( n24130 , n23080 , n23086 );
and ( n24131 , n23074 , n23086 );
or ( n24132 , n24129 , n24130 , n24131 );
and ( n24133 , n23076 , n23077 );
and ( n24134 , n23077 , n23079 );
and ( n24135 , n23076 , n23079 );
or ( n24136 , n24133 , n24134 , n24135 );
buf ( n24137 , n416 );
and ( n24138 , n599 , n24137 );
and ( n24139 , n608 , n23075 );
xor ( n24140 , n24138 , n24139 );
and ( n24141 , n611 , n22065 );
xor ( n24142 , n24140 , n24141 );
xor ( n24143 , n24136 , n24142 );
and ( n24144 , n632 , n20976 );
and ( n24145 , n671 , n20156 );
xor ( n24146 , n24144 , n24145 );
and ( n24147 , n715 , n19222 );
xor ( n24148 , n24146 , n24147 );
xor ( n24149 , n24143 , n24148 );
xor ( n24150 , n24132 , n24149 );
and ( n24151 , n23082 , n23083 );
and ( n24152 , n23083 , n23085 );
and ( n24153 , n23082 , n23085 );
or ( n24154 , n24151 , n24152 , n24153 );
and ( n24155 , n23098 , n23099 );
and ( n24156 , n23099 , n23101 );
and ( n24157 , n23098 , n23101 );
or ( n24158 , n24155 , n24156 , n24157 );
xor ( n24159 , n24154 , n24158 );
and ( n24160 , n783 , n18407 );
and ( n24161 , n856 , n17422 );
xor ( n24162 , n24160 , n24161 );
and ( n24163 , n925 , n16550 );
xor ( n24164 , n24162 , n24163 );
xor ( n24165 , n24159 , n24164 );
xor ( n24166 , n24150 , n24165 );
xor ( n24167 , n24128 , n24166 );
and ( n24168 , n23092 , n23096 );
and ( n24169 , n23096 , n23102 );
and ( n24170 , n23092 , n23102 );
or ( n24171 , n24168 , n24169 , n24170 );
and ( n24172 , n23118 , n23123 );
and ( n24173 , n23123 , n23129 );
and ( n24174 , n23118 , n23129 );
or ( n24175 , n24172 , n24173 , n24174 );
xor ( n24176 , n24171 , n24175 );
and ( n24177 , n23125 , n23126 );
and ( n24178 , n23126 , n23128 );
and ( n24179 , n23125 , n23128 );
or ( n24180 , n24177 , n24178 , n24179 );
and ( n24181 , n1383 , n13256 );
and ( n24182 , n1580 , n12531 );
xor ( n24183 , n24181 , n24182 );
and ( n24184 , n1694 , n11718 );
xor ( n24185 , n24183 , n24184 );
xor ( n24186 , n24180 , n24185 );
and ( n24187 , n1047 , n15691 );
and ( n24188 , n1164 , n14838 );
xor ( n24189 , n24187 , n24188 );
and ( n24190 , n1287 , n14044 );
xor ( n24191 , n24189 , n24190 );
xor ( n24192 , n24186 , n24191 );
xor ( n24193 , n24176 , n24192 );
xor ( n24194 , n24167 , n24193 );
xor ( n24195 , n24124 , n24194 );
xor ( n24196 , n24072 , n24195 );
xor ( n24197 , n23989 , n24196 );
xor ( n24198 , n23864 , n24197 );
and ( n24199 , n22863 , n22867 );
and ( n24200 , n22867 , n22973 );
and ( n24201 , n22863 , n22973 );
or ( n24202 , n24199 , n24200 , n24201 );
and ( n24203 , n23191 , n23200 );
xor ( n24204 , n24202 , n24203 );
and ( n24205 , n23195 , n23199 );
and ( n24206 , n22876 , n22896 );
and ( n24207 , n22896 , n22934 );
and ( n24208 , n22876 , n22934 );
or ( n24209 , n24206 , n24207 , n24208 );
and ( n24210 , n22880 , n22881 );
and ( n24211 , n22881 , n22895 );
and ( n24212 , n22880 , n22895 );
or ( n24213 , n24210 , n24211 , n24212 );
buf ( n24214 , n416 );
and ( n24215 , n24214 , n612 );
xor ( n24216 , n24213 , n24215 );
xor ( n24217 , n24209 , n24216 );
xor ( n24218 , n24205 , n24217 );
xor ( n24219 , n24204 , n24218 );
xor ( n24220 , n24198 , n24219 );
xor ( n24221 , n23860 , n24220 );
and ( n24222 , n22846 , n22850 );
and ( n24223 , n22850 , n23203 );
and ( n24224 , n22846 , n23203 );
or ( n24225 , n24222 , n24223 , n24224 );
xor ( n24226 , n24221 , n24225 );
and ( n24227 , n23204 , n23208 );
and ( n24228 , n23209 , n23212 );
or ( n24229 , n24227 , n24228 );
xor ( n24230 , n24226 , n24229 );
buf ( n24231 , n24230 );
buf ( n24232 , n24231 );
not ( n24233 , n24232 );
nor ( n24234 , n24233 , n8739 );
xor ( n24235 , n23851 , n24234 );
and ( n24236 , n22845 , n23217 );
and ( n24237 , n23218 , n23221 );
or ( n24238 , n24236 , n24237 );
xor ( n24239 , n24235 , n24238 );
buf ( n24240 , n24239 );
buf ( n24241 , n24240 );
not ( n24242 , n24241 );
buf ( n24243 , n553 );
not ( n24244 , n24243 );
nor ( n24245 , n24242 , n24244 );
xor ( n24246 , n23539 , n24245 );
xor ( n24247 , n23233 , n23536 );
nor ( n24248 , n23225 , n24244 );
and ( n24249 , n24247 , n24248 );
xor ( n24250 , n24247 , n24248 );
xor ( n24251 , n23237 , n23534 );
nor ( n24252 , n22231 , n24244 );
and ( n24253 , n24251 , n24252 );
xor ( n24254 , n24251 , n24252 );
xor ( n24255 , n23241 , n23532 );
nor ( n24256 , n21258 , n24244 );
and ( n24257 , n24255 , n24256 );
xor ( n24258 , n24255 , n24256 );
xor ( n24259 , n23245 , n23530 );
nor ( n24260 , n20303 , n24244 );
and ( n24261 , n24259 , n24260 );
xor ( n24262 , n24259 , n24260 );
xor ( n24263 , n23249 , n23528 );
nor ( n24264 , n19365 , n24244 );
and ( n24265 , n24263 , n24264 );
xor ( n24266 , n24263 , n24264 );
xor ( n24267 , n23253 , n23526 );
nor ( n24268 , n18448 , n24244 );
and ( n24269 , n24267 , n24268 );
xor ( n24270 , n24267 , n24268 );
xor ( n24271 , n23257 , n23524 );
nor ( n24272 , n17548 , n24244 );
and ( n24273 , n24271 , n24272 );
xor ( n24274 , n24271 , n24272 );
xor ( n24275 , n23261 , n23522 );
nor ( n24276 , n16669 , n24244 );
and ( n24277 , n24275 , n24276 );
xor ( n24278 , n24275 , n24276 );
xor ( n24279 , n23265 , n23520 );
nor ( n24280 , n15809 , n24244 );
and ( n24281 , n24279 , n24280 );
xor ( n24282 , n24279 , n24280 );
xor ( n24283 , n23269 , n23518 );
nor ( n24284 , n14968 , n24244 );
and ( n24285 , n24283 , n24284 );
xor ( n24286 , n24283 , n24284 );
xor ( n24287 , n23273 , n23516 );
nor ( n24288 , n14147 , n24244 );
and ( n24289 , n24287 , n24288 );
xor ( n24290 , n24287 , n24288 );
xor ( n24291 , n23277 , n23514 );
nor ( n24292 , n13349 , n24244 );
and ( n24293 , n24291 , n24292 );
xor ( n24294 , n24291 , n24292 );
xor ( n24295 , n23281 , n23512 );
nor ( n24296 , n12564 , n24244 );
and ( n24297 , n24295 , n24296 );
xor ( n24298 , n24295 , n24296 );
xor ( n24299 , n23285 , n23510 );
nor ( n24300 , n11799 , n24244 );
and ( n24301 , n24299 , n24300 );
xor ( n24302 , n24299 , n24300 );
xor ( n24303 , n23289 , n23508 );
nor ( n24304 , n11050 , n24244 );
and ( n24305 , n24303 , n24304 );
xor ( n24306 , n24303 , n24304 );
xor ( n24307 , n23293 , n23506 );
nor ( n24308 , n10321 , n24244 );
and ( n24309 , n24307 , n24308 );
xor ( n24310 , n24307 , n24308 );
xor ( n24311 , n23297 , n23504 );
nor ( n24312 , n9429 , n24244 );
and ( n24313 , n24311 , n24312 );
xor ( n24314 , n24311 , n24312 );
xor ( n24315 , n23301 , n23502 );
nor ( n24316 , n8949 , n24244 );
and ( n24317 , n24315 , n24316 );
xor ( n24318 , n24315 , n24316 );
xor ( n24319 , n23305 , n23500 );
nor ( n24320 , n9437 , n24244 );
and ( n24321 , n24319 , n24320 );
xor ( n24322 , n24319 , n24320 );
xor ( n24323 , n23309 , n23498 );
nor ( n24324 , n9446 , n24244 );
and ( n24325 , n24323 , n24324 );
xor ( n24326 , n24323 , n24324 );
xor ( n24327 , n23313 , n23496 );
nor ( n24328 , n9455 , n24244 );
and ( n24329 , n24327 , n24328 );
xor ( n24330 , n24327 , n24328 );
xor ( n24331 , n23317 , n23494 );
nor ( n24332 , n9464 , n24244 );
and ( n24333 , n24331 , n24332 );
xor ( n24334 , n24331 , n24332 );
xor ( n24335 , n23321 , n23492 );
nor ( n24336 , n9473 , n24244 );
and ( n24337 , n24335 , n24336 );
xor ( n24338 , n24335 , n24336 );
xor ( n24339 , n23325 , n23490 );
nor ( n24340 , n9482 , n24244 );
and ( n24341 , n24339 , n24340 );
xor ( n24342 , n24339 , n24340 );
xor ( n24343 , n23329 , n23488 );
nor ( n24344 , n9491 , n24244 );
and ( n24345 , n24343 , n24344 );
xor ( n24346 , n24343 , n24344 );
xor ( n24347 , n23333 , n23486 );
nor ( n24348 , n9500 , n24244 );
and ( n24349 , n24347 , n24348 );
xor ( n24350 , n24347 , n24348 );
xor ( n24351 , n23337 , n23484 );
nor ( n24352 , n9509 , n24244 );
and ( n24353 , n24351 , n24352 );
xor ( n24354 , n24351 , n24352 );
xor ( n24355 , n23341 , n23482 );
nor ( n24356 , n9518 , n24244 );
and ( n24357 , n24355 , n24356 );
xor ( n24358 , n24355 , n24356 );
xor ( n24359 , n23345 , n23480 );
nor ( n24360 , n9527 , n24244 );
and ( n24361 , n24359 , n24360 );
xor ( n24362 , n24359 , n24360 );
xor ( n24363 , n23349 , n23478 );
nor ( n24364 , n9536 , n24244 );
and ( n24365 , n24363 , n24364 );
xor ( n24366 , n24363 , n24364 );
xor ( n24367 , n23353 , n23476 );
nor ( n24368 , n9545 , n24244 );
and ( n24369 , n24367 , n24368 );
xor ( n24370 , n24367 , n24368 );
xor ( n24371 , n23357 , n23474 );
nor ( n24372 , n9554 , n24244 );
and ( n24373 , n24371 , n24372 );
xor ( n24374 , n24371 , n24372 );
xor ( n24375 , n23361 , n23472 );
nor ( n24376 , n9563 , n24244 );
and ( n24377 , n24375 , n24376 );
xor ( n24378 , n24375 , n24376 );
xor ( n24379 , n23365 , n23470 );
nor ( n24380 , n9572 , n24244 );
and ( n24381 , n24379 , n24380 );
xor ( n24382 , n24379 , n24380 );
xor ( n24383 , n23369 , n23468 );
nor ( n24384 , n9581 , n24244 );
and ( n24385 , n24383 , n24384 );
xor ( n24386 , n24383 , n24384 );
xor ( n24387 , n23373 , n23466 );
nor ( n24388 , n9590 , n24244 );
and ( n24389 , n24387 , n24388 );
xor ( n24390 , n24387 , n24388 );
xor ( n24391 , n23377 , n23464 );
nor ( n24392 , n9599 , n24244 );
and ( n24393 , n24391 , n24392 );
xor ( n24394 , n24391 , n24392 );
xor ( n24395 , n23381 , n23462 );
nor ( n24396 , n9608 , n24244 );
and ( n24397 , n24395 , n24396 );
xor ( n24398 , n24395 , n24396 );
xor ( n24399 , n23385 , n23460 );
nor ( n24400 , n9617 , n24244 );
and ( n24401 , n24399 , n24400 );
xor ( n24402 , n24399 , n24400 );
xor ( n24403 , n23389 , n23458 );
nor ( n24404 , n9626 , n24244 );
and ( n24405 , n24403 , n24404 );
xor ( n24406 , n24403 , n24404 );
xor ( n24407 , n23393 , n23456 );
nor ( n24408 , n9635 , n24244 );
and ( n24409 , n24407 , n24408 );
xor ( n24410 , n24407 , n24408 );
xor ( n24411 , n23397 , n23454 );
nor ( n24412 , n9644 , n24244 );
and ( n24413 , n24411 , n24412 );
xor ( n24414 , n24411 , n24412 );
xor ( n24415 , n23401 , n23452 );
nor ( n24416 , n9653 , n24244 );
and ( n24417 , n24415 , n24416 );
xor ( n24418 , n24415 , n24416 );
xor ( n24419 , n23405 , n23450 );
nor ( n24420 , n9662 , n24244 );
and ( n24421 , n24419 , n24420 );
xor ( n24422 , n24419 , n24420 );
xor ( n24423 , n23409 , n23448 );
nor ( n24424 , n9671 , n24244 );
and ( n24425 , n24423 , n24424 );
xor ( n24426 , n24423 , n24424 );
xor ( n24427 , n23413 , n23446 );
nor ( n24428 , n9680 , n24244 );
and ( n24429 , n24427 , n24428 );
xor ( n24430 , n24427 , n24428 );
xor ( n24431 , n23417 , n23444 );
nor ( n24432 , n9689 , n24244 );
and ( n24433 , n24431 , n24432 );
xor ( n24434 , n24431 , n24432 );
xor ( n24435 , n23421 , n23442 );
nor ( n24436 , n9698 , n24244 );
and ( n24437 , n24435 , n24436 );
xor ( n24438 , n24435 , n24436 );
xor ( n24439 , n23425 , n23440 );
nor ( n24440 , n9707 , n24244 );
and ( n24441 , n24439 , n24440 );
xor ( n24442 , n24439 , n24440 );
xor ( n24443 , n23429 , n23438 );
nor ( n24444 , n9716 , n24244 );
and ( n24445 , n24443 , n24444 );
xor ( n24446 , n24443 , n24444 );
xor ( n24447 , n23433 , n23436 );
nor ( n24448 , n9725 , n24244 );
and ( n24449 , n24447 , n24448 );
xor ( n24450 , n24447 , n24448 );
xor ( n24451 , n23434 , n23435 );
nor ( n24452 , n9734 , n24244 );
and ( n24453 , n24451 , n24452 );
xor ( n24454 , n24451 , n24452 );
nor ( n24455 , n9752 , n23227 );
nor ( n24456 , n9743 , n24244 );
and ( n24457 , n24455 , n24456 );
and ( n24458 , n24454 , n24457 );
or ( n24459 , n24453 , n24458 );
and ( n24460 , n24450 , n24459 );
or ( n24461 , n24449 , n24460 );
and ( n24462 , n24446 , n24461 );
or ( n24463 , n24445 , n24462 );
and ( n24464 , n24442 , n24463 );
or ( n24465 , n24441 , n24464 );
and ( n24466 , n24438 , n24465 );
or ( n24467 , n24437 , n24466 );
and ( n24468 , n24434 , n24467 );
or ( n24469 , n24433 , n24468 );
and ( n24470 , n24430 , n24469 );
or ( n24471 , n24429 , n24470 );
and ( n24472 , n24426 , n24471 );
or ( n24473 , n24425 , n24472 );
and ( n24474 , n24422 , n24473 );
or ( n24475 , n24421 , n24474 );
and ( n24476 , n24418 , n24475 );
or ( n24477 , n24417 , n24476 );
and ( n24478 , n24414 , n24477 );
or ( n24479 , n24413 , n24478 );
and ( n24480 , n24410 , n24479 );
or ( n24481 , n24409 , n24480 );
and ( n24482 , n24406 , n24481 );
or ( n24483 , n24405 , n24482 );
and ( n24484 , n24402 , n24483 );
or ( n24485 , n24401 , n24484 );
and ( n24486 , n24398 , n24485 );
or ( n24487 , n24397 , n24486 );
and ( n24488 , n24394 , n24487 );
or ( n24489 , n24393 , n24488 );
and ( n24490 , n24390 , n24489 );
or ( n24491 , n24389 , n24490 );
and ( n24492 , n24386 , n24491 );
or ( n24493 , n24385 , n24492 );
and ( n24494 , n24382 , n24493 );
or ( n24495 , n24381 , n24494 );
and ( n24496 , n24378 , n24495 );
or ( n24497 , n24377 , n24496 );
and ( n24498 , n24374 , n24497 );
or ( n24499 , n24373 , n24498 );
and ( n24500 , n24370 , n24499 );
or ( n24501 , n24369 , n24500 );
and ( n24502 , n24366 , n24501 );
or ( n24503 , n24365 , n24502 );
and ( n24504 , n24362 , n24503 );
or ( n24505 , n24361 , n24504 );
and ( n24506 , n24358 , n24505 );
or ( n24507 , n24357 , n24506 );
and ( n24508 , n24354 , n24507 );
or ( n24509 , n24353 , n24508 );
and ( n24510 , n24350 , n24509 );
or ( n24511 , n24349 , n24510 );
and ( n24512 , n24346 , n24511 );
or ( n24513 , n24345 , n24512 );
and ( n24514 , n24342 , n24513 );
or ( n24515 , n24341 , n24514 );
and ( n24516 , n24338 , n24515 );
or ( n24517 , n24337 , n24516 );
and ( n24518 , n24334 , n24517 );
or ( n24519 , n24333 , n24518 );
and ( n24520 , n24330 , n24519 );
or ( n24521 , n24329 , n24520 );
and ( n24522 , n24326 , n24521 );
or ( n24523 , n24325 , n24522 );
and ( n24524 , n24322 , n24523 );
or ( n24525 , n24321 , n24524 );
and ( n24526 , n24318 , n24525 );
or ( n24527 , n24317 , n24526 );
and ( n24528 , n24314 , n24527 );
or ( n24529 , n24313 , n24528 );
and ( n24530 , n24310 , n24529 );
or ( n24531 , n24309 , n24530 );
and ( n24532 , n24306 , n24531 );
or ( n24533 , n24305 , n24532 );
and ( n24534 , n24302 , n24533 );
or ( n24535 , n24301 , n24534 );
and ( n24536 , n24298 , n24535 );
or ( n24537 , n24297 , n24536 );
and ( n24538 , n24294 , n24537 );
or ( n24539 , n24293 , n24538 );
and ( n24540 , n24290 , n24539 );
or ( n24541 , n24289 , n24540 );
and ( n24542 , n24286 , n24541 );
or ( n24543 , n24285 , n24542 );
and ( n24544 , n24282 , n24543 );
or ( n24545 , n24281 , n24544 );
and ( n24546 , n24278 , n24545 );
or ( n24547 , n24277 , n24546 );
and ( n24548 , n24274 , n24547 );
or ( n24549 , n24273 , n24548 );
and ( n24550 , n24270 , n24549 );
or ( n24551 , n24269 , n24550 );
and ( n24552 , n24266 , n24551 );
or ( n24553 , n24265 , n24552 );
and ( n24554 , n24262 , n24553 );
or ( n24555 , n24261 , n24554 );
and ( n24556 , n24258 , n24555 );
or ( n24557 , n24257 , n24556 );
and ( n24558 , n24254 , n24557 );
or ( n24559 , n24253 , n24558 );
and ( n24560 , n24250 , n24559 );
or ( n24561 , n24249 , n24560 );
xor ( n24562 , n24246 , n24561 );
buf ( n24563 , n479 );
not ( n24564 , n24563 );
nor ( n24565 , n601 , n24564 );
buf ( n24566 , n24565 );
nor ( n24567 , n622 , n22541 );
xor ( n24568 , n24566 , n24567 );
buf ( n24569 , n24568 );
nor ( n24570 , n646 , n21562 );
xor ( n24571 , n24569 , n24570 );
and ( n24572 , n23543 , n23544 );
buf ( n24573 , n24572 );
xor ( n24574 , n24571 , n24573 );
nor ( n24575 , n684 , n20601 );
xor ( n24576 , n24574 , n24575 );
and ( n24577 , n23546 , n23547 );
and ( n24578 , n23548 , n23550 );
or ( n24579 , n24577 , n24578 );
xor ( n24580 , n24576 , n24579 );
nor ( n24581 , n733 , n19657 );
xor ( n24582 , n24580 , n24581 );
and ( n24583 , n23551 , n23552 );
and ( n24584 , n23553 , n23556 );
or ( n24585 , n24583 , n24584 );
xor ( n24586 , n24582 , n24585 );
nor ( n24587 , n796 , n18734 );
xor ( n24588 , n24586 , n24587 );
and ( n24589 , n23557 , n23558 );
and ( n24590 , n23559 , n23562 );
or ( n24591 , n24589 , n24590 );
xor ( n24592 , n24588 , n24591 );
nor ( n24593 , n868 , n17828 );
xor ( n24594 , n24592 , n24593 );
and ( n24595 , n23563 , n23564 );
and ( n24596 , n23565 , n23568 );
or ( n24597 , n24595 , n24596 );
xor ( n24598 , n24594 , n24597 );
nor ( n24599 , n958 , n16943 );
xor ( n24600 , n24598 , n24599 );
and ( n24601 , n23569 , n23570 );
and ( n24602 , n23571 , n23574 );
or ( n24603 , n24601 , n24602 );
xor ( n24604 , n24600 , n24603 );
nor ( n24605 , n1062 , n16077 );
xor ( n24606 , n24604 , n24605 );
and ( n24607 , n23575 , n23576 );
and ( n24608 , n23577 , n23580 );
or ( n24609 , n24607 , n24608 );
xor ( n24610 , n24606 , n24609 );
nor ( n24611 , n1176 , n15230 );
xor ( n24612 , n24610 , n24611 );
and ( n24613 , n23581 , n23582 );
and ( n24614 , n23583 , n23586 );
or ( n24615 , n24613 , n24614 );
xor ( n24616 , n24612 , n24615 );
nor ( n24617 , n1303 , n14403 );
xor ( n24618 , n24616 , n24617 );
and ( n24619 , n23587 , n23588 );
and ( n24620 , n23589 , n23592 );
or ( n24621 , n24619 , n24620 );
xor ( n24622 , n24618 , n24621 );
nor ( n24623 , n1445 , n13599 );
xor ( n24624 , n24622 , n24623 );
and ( n24625 , n23593 , n23594 );
and ( n24626 , n23595 , n23598 );
or ( n24627 , n24625 , n24626 );
xor ( n24628 , n24624 , n24627 );
nor ( n24629 , n1598 , n12808 );
xor ( n24630 , n24628 , n24629 );
and ( n24631 , n23599 , n23600 );
and ( n24632 , n23601 , n23604 );
or ( n24633 , n24631 , n24632 );
xor ( n24634 , n24630 , n24633 );
nor ( n24635 , n1766 , n12037 );
xor ( n24636 , n24634 , n24635 );
and ( n24637 , n23605 , n23606 );
and ( n24638 , n23607 , n23610 );
or ( n24639 , n24637 , n24638 );
xor ( n24640 , n24636 , n24639 );
nor ( n24641 , n1945 , n11282 );
xor ( n24642 , n24640 , n24641 );
and ( n24643 , n23611 , n23612 );
and ( n24644 , n23613 , n23616 );
or ( n24645 , n24643 , n24644 );
xor ( n24646 , n24642 , n24645 );
nor ( n24647 , n2137 , n10547 );
xor ( n24648 , n24646 , n24647 );
and ( n24649 , n23617 , n23618 );
and ( n24650 , n23619 , n23622 );
or ( n24651 , n24649 , n24650 );
xor ( n24652 , n24648 , n24651 );
nor ( n24653 , n2343 , n9829 );
xor ( n24654 , n24652 , n24653 );
and ( n24655 , n23623 , n23624 );
and ( n24656 , n23625 , n23628 );
or ( n24657 , n24655 , n24656 );
xor ( n24658 , n24654 , n24657 );
nor ( n24659 , n2566 , n8955 );
xor ( n24660 , n24658 , n24659 );
and ( n24661 , n23629 , n23630 );
and ( n24662 , n23631 , n23634 );
or ( n24663 , n24661 , n24662 );
xor ( n24664 , n24660 , n24663 );
nor ( n24665 , n2797 , n603 );
xor ( n24666 , n24664 , n24665 );
and ( n24667 , n23635 , n23636 );
and ( n24668 , n23637 , n23640 );
or ( n24669 , n24667 , n24668 );
xor ( n24670 , n24666 , n24669 );
nor ( n24671 , n3043 , n652 );
xor ( n24672 , n24670 , n24671 );
and ( n24673 , n23641 , n23642 );
and ( n24674 , n23643 , n23646 );
or ( n24675 , n24673 , n24674 );
xor ( n24676 , n24672 , n24675 );
nor ( n24677 , n3300 , n624 );
xor ( n24678 , n24676 , n24677 );
and ( n24679 , n23647 , n23648 );
and ( n24680 , n23649 , n23652 );
or ( n24681 , n24679 , n24680 );
xor ( n24682 , n24678 , n24681 );
nor ( n24683 , n3570 , n648 );
xor ( n24684 , n24682 , n24683 );
and ( n24685 , n23653 , n23654 );
and ( n24686 , n23655 , n23658 );
or ( n24687 , n24685 , n24686 );
xor ( n24688 , n24684 , n24687 );
nor ( n24689 , n3853 , n686 );
xor ( n24690 , n24688 , n24689 );
and ( n24691 , n23659 , n23660 );
and ( n24692 , n23661 , n23664 );
or ( n24693 , n24691 , n24692 );
xor ( n24694 , n24690 , n24693 );
nor ( n24695 , n4151 , n735 );
xor ( n24696 , n24694 , n24695 );
and ( n24697 , n23665 , n23666 );
and ( n24698 , n23667 , n23670 );
or ( n24699 , n24697 , n24698 );
xor ( n24700 , n24696 , n24699 );
nor ( n24701 , n4458 , n798 );
xor ( n24702 , n24700 , n24701 );
and ( n24703 , n23671 , n23672 );
and ( n24704 , n23673 , n23676 );
or ( n24705 , n24703 , n24704 );
xor ( n24706 , n24702 , n24705 );
nor ( n24707 , n4786 , n870 );
xor ( n24708 , n24706 , n24707 );
and ( n24709 , n23677 , n23678 );
and ( n24710 , n23679 , n23682 );
or ( n24711 , n24709 , n24710 );
xor ( n24712 , n24708 , n24711 );
nor ( n24713 , n5126 , n960 );
xor ( n24714 , n24712 , n24713 );
and ( n24715 , n23683 , n23684 );
and ( n24716 , n23685 , n23688 );
or ( n24717 , n24715 , n24716 );
xor ( n24718 , n24714 , n24717 );
nor ( n24719 , n5477 , n1064 );
xor ( n24720 , n24718 , n24719 );
and ( n24721 , n23689 , n23690 );
and ( n24722 , n23691 , n23694 );
or ( n24723 , n24721 , n24722 );
xor ( n24724 , n24720 , n24723 );
nor ( n24725 , n5838 , n1178 );
xor ( n24726 , n24724 , n24725 );
and ( n24727 , n23695 , n23696 );
and ( n24728 , n23697 , n23700 );
or ( n24729 , n24727 , n24728 );
xor ( n24730 , n24726 , n24729 );
nor ( n24731 , n6212 , n1305 );
xor ( n24732 , n24730 , n24731 );
and ( n24733 , n23701 , n23702 );
and ( n24734 , n23703 , n23706 );
or ( n24735 , n24733 , n24734 );
xor ( n24736 , n24732 , n24735 );
nor ( n24737 , n6596 , n1447 );
xor ( n24738 , n24736 , n24737 );
and ( n24739 , n23707 , n23708 );
and ( n24740 , n23709 , n23712 );
or ( n24741 , n24739 , n24740 );
xor ( n24742 , n24738 , n24741 );
nor ( n24743 , n6997 , n1600 );
xor ( n24744 , n24742 , n24743 );
and ( n24745 , n23713 , n23714 );
and ( n24746 , n23715 , n23718 );
or ( n24747 , n24745 , n24746 );
xor ( n24748 , n24744 , n24747 );
nor ( n24749 , n7413 , n1768 );
xor ( n24750 , n24748 , n24749 );
and ( n24751 , n23719 , n23720 );
and ( n24752 , n23721 , n23724 );
or ( n24753 , n24751 , n24752 );
xor ( n24754 , n24750 , n24753 );
nor ( n24755 , n7841 , n1947 );
xor ( n24756 , n24754 , n24755 );
and ( n24757 , n23725 , n23726 );
and ( n24758 , n23727 , n23730 );
or ( n24759 , n24757 , n24758 );
xor ( n24760 , n24756 , n24759 );
nor ( n24761 , n8281 , n2139 );
xor ( n24762 , n24760 , n24761 );
and ( n24763 , n23731 , n23732 );
and ( n24764 , n23733 , n23736 );
or ( n24765 , n24763 , n24764 );
xor ( n24766 , n24762 , n24765 );
nor ( n24767 , n8737 , n2345 );
xor ( n24768 , n24766 , n24767 );
and ( n24769 , n23737 , n23738 );
and ( n24770 , n23739 , n23742 );
or ( n24771 , n24769 , n24770 );
xor ( n24772 , n24768 , n24771 );
nor ( n24773 , n9420 , n2568 );
xor ( n24774 , n24772 , n24773 );
and ( n24775 , n23743 , n23744 );
and ( n24776 , n23745 , n23748 );
or ( n24777 , n24775 , n24776 );
xor ( n24778 , n24774 , n24777 );
nor ( n24779 , n10312 , n2799 );
xor ( n24780 , n24778 , n24779 );
and ( n24781 , n23749 , n23750 );
and ( n24782 , n23751 , n23754 );
or ( n24783 , n24781 , n24782 );
xor ( n24784 , n24780 , n24783 );
nor ( n24785 , n11041 , n3045 );
xor ( n24786 , n24784 , n24785 );
and ( n24787 , n23755 , n23756 );
and ( n24788 , n23757 , n23760 );
or ( n24789 , n24787 , n24788 );
xor ( n24790 , n24786 , n24789 );
nor ( n24791 , n11790 , n3302 );
xor ( n24792 , n24790 , n24791 );
and ( n24793 , n23761 , n23762 );
and ( n24794 , n23763 , n23766 );
or ( n24795 , n24793 , n24794 );
xor ( n24796 , n24792 , n24795 );
nor ( n24797 , n12555 , n3572 );
xor ( n24798 , n24796 , n24797 );
and ( n24799 , n23767 , n23768 );
and ( n24800 , n23769 , n23772 );
or ( n24801 , n24799 , n24800 );
xor ( n24802 , n24798 , n24801 );
nor ( n24803 , n13340 , n3855 );
xor ( n24804 , n24802 , n24803 );
and ( n24805 , n23773 , n23774 );
and ( n24806 , n23775 , n23778 );
or ( n24807 , n24805 , n24806 );
xor ( n24808 , n24804 , n24807 );
nor ( n24809 , n14138 , n4153 );
xor ( n24810 , n24808 , n24809 );
and ( n24811 , n23779 , n23780 );
and ( n24812 , n23781 , n23784 );
or ( n24813 , n24811 , n24812 );
xor ( n24814 , n24810 , n24813 );
nor ( n24815 , n14959 , n4460 );
xor ( n24816 , n24814 , n24815 );
and ( n24817 , n23785 , n23786 );
and ( n24818 , n23787 , n23790 );
or ( n24819 , n24817 , n24818 );
xor ( n24820 , n24816 , n24819 );
nor ( n24821 , n15800 , n4788 );
xor ( n24822 , n24820 , n24821 );
and ( n24823 , n23791 , n23792 );
and ( n24824 , n23793 , n23796 );
or ( n24825 , n24823 , n24824 );
xor ( n24826 , n24822 , n24825 );
nor ( n24827 , n16660 , n5128 );
xor ( n24828 , n24826 , n24827 );
and ( n24829 , n23797 , n23798 );
and ( n24830 , n23799 , n23802 );
or ( n24831 , n24829 , n24830 );
xor ( n24832 , n24828 , n24831 );
nor ( n24833 , n17539 , n5479 );
xor ( n24834 , n24832 , n24833 );
and ( n24835 , n23803 , n23804 );
and ( n24836 , n23805 , n23808 );
or ( n24837 , n24835 , n24836 );
xor ( n24838 , n24834 , n24837 );
nor ( n24839 , n18439 , n5840 );
xor ( n24840 , n24838 , n24839 );
and ( n24841 , n23809 , n23810 );
and ( n24842 , n23811 , n23814 );
or ( n24843 , n24841 , n24842 );
xor ( n24844 , n24840 , n24843 );
nor ( n24845 , n19356 , n6214 );
xor ( n24846 , n24844 , n24845 );
and ( n24847 , n23815 , n23816 );
and ( n24848 , n23817 , n23820 );
or ( n24849 , n24847 , n24848 );
xor ( n24850 , n24846 , n24849 );
nor ( n24851 , n20294 , n6598 );
xor ( n24852 , n24850 , n24851 );
and ( n24853 , n23821 , n23822 );
and ( n24854 , n23823 , n23826 );
or ( n24855 , n24853 , n24854 );
xor ( n24856 , n24852 , n24855 );
nor ( n24857 , n21249 , n6999 );
xor ( n24858 , n24856 , n24857 );
and ( n24859 , n23827 , n23828 );
and ( n24860 , n23829 , n23832 );
or ( n24861 , n24859 , n24860 );
xor ( n24862 , n24858 , n24861 );
nor ( n24863 , n22222 , n7415 );
xor ( n24864 , n24862 , n24863 );
and ( n24865 , n23833 , n23834 );
and ( n24866 , n23835 , n23838 );
or ( n24867 , n24865 , n24866 );
xor ( n24868 , n24864 , n24867 );
nor ( n24869 , n23216 , n7843 );
xor ( n24870 , n24868 , n24869 );
and ( n24871 , n23839 , n23840 );
and ( n24872 , n23841 , n23844 );
or ( n24873 , n24871 , n24872 );
xor ( n24874 , n24870 , n24873 );
nor ( n24875 , n24233 , n8283 );
xor ( n24876 , n24874 , n24875 );
and ( n24877 , n23845 , n23846 );
and ( n24878 , n23847 , n23850 );
or ( n24879 , n24877 , n24878 );
xor ( n24880 , n24876 , n24879 );
and ( n24881 , n24202 , n24203 );
and ( n24882 , n24203 , n24218 );
and ( n24883 , n24202 , n24218 );
or ( n24884 , n24881 , n24882 , n24883 );
and ( n24885 , n23864 , n24197 );
and ( n24886 , n24197 , n24219 );
and ( n24887 , n23864 , n24219 );
or ( n24888 , n24885 , n24886 , n24887 );
xor ( n24889 , n24884 , n24888 );
and ( n24890 , n23868 , n23988 );
and ( n24891 , n23988 , n24196 );
and ( n24892 , n23868 , n24196 );
or ( n24893 , n24890 , n24891 , n24892 );
and ( n24894 , n23993 , n24071 );
and ( n24895 , n24071 , n24195 );
and ( n24896 , n23993 , n24195 );
or ( n24897 , n24894 , n24895 , n24896 );
and ( n24898 , n23881 , n23949 );
and ( n24899 , n23949 , n23986 );
and ( n24900 , n23881 , n23986 );
or ( n24901 , n24898 , n24899 , n24900 );
and ( n24902 , n23997 , n24001 );
and ( n24903 , n24001 , n24070 );
and ( n24904 , n23997 , n24070 );
or ( n24905 , n24902 , n24903 , n24904 );
xor ( n24906 , n24901 , n24905 );
and ( n24907 , n23954 , n23958 );
and ( n24908 , n23958 , n23985 );
and ( n24909 , n23954 , n23985 );
or ( n24910 , n24907 , n24908 , n24909 );
and ( n24911 , n23915 , n23931 );
and ( n24912 , n23931 , n23947 );
and ( n24913 , n23915 , n23947 );
or ( n24914 , n24911 , n24912 , n24913 );
and ( n24915 , n23898 , n23902 );
and ( n24916 , n23902 , n23908 );
and ( n24917 , n23898 , n23908 );
or ( n24918 , n24915 , n24916 , n24917 );
and ( n24919 , n23919 , n23924 );
and ( n24920 , n23924 , n23930 );
and ( n24921 , n23919 , n23930 );
or ( n24922 , n24919 , n24920 , n24921 );
xor ( n24923 , n24918 , n24922 );
and ( n24924 , n23904 , n23905 );
and ( n24925 , n23905 , n23907 );
and ( n24926 , n23904 , n23907 );
or ( n24927 , n24924 , n24925 , n24926 );
and ( n24928 , n23920 , n23921 );
and ( n24929 , n23921 , n23923 );
and ( n24930 , n23920 , n23923 );
or ( n24931 , n24928 , n24929 , n24930 );
xor ( n24932 , n24927 , n24931 );
and ( n24933 , n21216 , n663 );
and ( n24934 , n22186 , n635 );
xor ( n24935 , n24933 , n24934 );
and ( n24936 , n22892 , n606 );
xor ( n24937 , n24935 , n24936 );
xor ( n24938 , n24932 , n24937 );
xor ( n24939 , n24923 , n24938 );
xor ( n24940 , n24914 , n24939 );
and ( n24941 , n23936 , n23940 );
and ( n24942 , n23940 , n23946 );
and ( n24943 , n23936 , n23946 );
or ( n24944 , n24941 , n24942 , n24943 );
and ( n24945 , n23926 , n23927 );
and ( n24946 , n23927 , n23929 );
and ( n24947 , n23926 , n23929 );
or ( n24948 , n24945 , n24946 , n24947 );
and ( n24949 , n18144 , n840 );
and ( n24950 , n19324 , n771 );
xor ( n24951 , n24949 , n24950 );
and ( n24952 , n20233 , n719 );
xor ( n24953 , n24951 , n24952 );
xor ( n24954 , n24948 , n24953 );
and ( n24955 , n15758 , n1134 );
and ( n24956 , n16637 , n1034 );
xor ( n24957 , n24955 , n24956 );
and ( n24958 , n17512 , n940 );
xor ( n24959 , n24957 , n24958 );
xor ( n24960 , n24954 , n24959 );
xor ( n24961 , n24944 , n24960 );
and ( n24962 , n23942 , n23943 );
and ( n24963 , n23943 , n23945 );
and ( n24964 , n23942 , n23945 );
or ( n24965 , n24962 , n24963 , n24964 );
and ( n24966 , n23973 , n23974 );
and ( n24967 , n23974 , n23976 );
and ( n24968 , n23973 , n23976 );
or ( n24969 , n24966 , n24967 , n24968 );
xor ( n24970 , n24965 , n24969 );
and ( n24971 , n13322 , n1551 );
and ( n24972 , n14118 , n1424 );
xor ( n24973 , n24971 , n24972 );
and ( n24974 , n14938 , n1254 );
xor ( n24975 , n24973 , n24974 );
xor ( n24976 , n24970 , n24975 );
xor ( n24977 , n24961 , n24976 );
xor ( n24978 , n24940 , n24977 );
xor ( n24979 , n24910 , n24978 );
and ( n24980 , n23963 , n23967 );
and ( n24981 , n23967 , n23984 );
and ( n24982 , n23963 , n23984 );
or ( n24983 , n24980 , n24981 , n24982 );
and ( n24984 , n24036 , n24051 );
and ( n24985 , n24051 , n24068 );
and ( n24986 , n24036 , n24068 );
or ( n24987 , n24984 , n24985 , n24986 );
xor ( n24988 , n24983 , n24987 );
and ( n24989 , n23972 , n23977 );
and ( n24990 , n23977 , n23983 );
and ( n24991 , n23972 , n23983 );
or ( n24992 , n24989 , n24990 , n24991 );
and ( n24993 , n24040 , n24044 );
and ( n24994 , n24044 , n24050 );
and ( n24995 , n24040 , n24050 );
or ( n24996 , n24993 , n24994 , n24995 );
xor ( n24997 , n24992 , n24996 );
and ( n24998 , n23979 , n23980 );
and ( n24999 , n23980 , n23982 );
and ( n25000 , n23979 , n23982 );
or ( n25001 , n24998 , n24999 , n25000 );
and ( n25002 , n11015 , n2100 );
and ( n25003 , n11769 , n1882 );
xor ( n25004 , n25002 , n25003 );
and ( n25005 , n12320 , n1738 );
xor ( n25006 , n25004 , n25005 );
xor ( n25007 , n25001 , n25006 );
and ( n25008 , n8718 , n2739 );
and ( n25009 , n9400 , n2544 );
xor ( n25010 , n25008 , n25009 );
and ( n25011 , n10291 , n2298 );
xor ( n25012 , n25010 , n25011 );
xor ( n25013 , n25007 , n25012 );
xor ( n25014 , n24997 , n25013 );
xor ( n25015 , n24988 , n25014 );
xor ( n25016 , n24979 , n25015 );
xor ( n25017 , n24906 , n25016 );
xor ( n25018 , n24897 , n25017 );
and ( n25019 , n24076 , n24123 );
and ( n25020 , n24123 , n24194 );
and ( n25021 , n24076 , n24194 );
or ( n25022 , n25019 , n25020 , n25021 );
and ( n25023 , n24006 , n24031 );
and ( n25024 , n24031 , n24069 );
and ( n25025 , n24006 , n24069 );
or ( n25026 , n25023 , n25024 , n25025 );
and ( n25027 , n24080 , n24084 );
and ( n25028 , n24084 , n24122 );
and ( n25029 , n24080 , n24122 );
or ( n25030 , n25027 , n25028 , n25029 );
xor ( n25031 , n25026 , n25030 );
and ( n25032 , n24010 , n24014 );
and ( n25033 , n24014 , n24030 );
and ( n25034 , n24010 , n24030 );
or ( n25035 , n25032 , n25033 , n25034 );
and ( n25036 , n24109 , n24114 );
and ( n25037 , n24114 , n24120 );
and ( n25038 , n24109 , n24120 );
or ( n25039 , n25036 , n25037 , n25038 );
and ( n25040 , n24019 , n24023 );
and ( n25041 , n24023 , n24029 );
and ( n25042 , n24019 , n24029 );
or ( n25043 , n25040 , n25041 , n25042 );
xor ( n25044 , n25039 , n25043 );
and ( n25045 , n24025 , n24026 );
and ( n25046 , n24026 , n24028 );
and ( n25047 , n24025 , n24028 );
or ( n25048 , n25045 , n25046 , n25047 );
and ( n25049 , n24116 , n24117 );
and ( n25050 , n24117 , n24119 );
and ( n25051 , n24116 , n24119 );
or ( n25052 , n25049 , n25050 , n25051 );
xor ( n25053 , n25048 , n25052 );
and ( n25054 , n4132 , n6504 );
and ( n25055 , n4438 , n6132 );
xor ( n25056 , n25054 , n25055 );
and ( n25057 , n4766 , n5765 );
xor ( n25058 , n25056 , n25057 );
xor ( n25059 , n25053 , n25058 );
xor ( n25060 , n25044 , n25059 );
xor ( n25061 , n25035 , n25060 );
and ( n25062 , n24056 , n24061 );
and ( n25063 , n24061 , n24067 );
and ( n25064 , n24056 , n24067 );
or ( n25065 , n25062 , n25063 , n25064 );
and ( n25066 , n24046 , n24047 );
and ( n25067 , n24047 , n24049 );
and ( n25068 , n24046 , n24049 );
or ( n25069 , n25066 , n25067 , n25068 );
and ( n25070 , n24057 , n24058 );
and ( n25071 , n24058 , n24060 );
and ( n25072 , n24057 , n24060 );
or ( n25073 , n25070 , n25071 , n25072 );
xor ( n25074 , n25069 , n25073 );
and ( n25075 , n7385 , n3495 );
and ( n25076 , n7808 , n3271 );
xor ( n25077 , n25075 , n25076 );
and ( n25078 , n8079 , n2981 );
xor ( n25079 , n25077 , n25078 );
xor ( n25080 , n25074 , n25079 );
xor ( n25081 , n25065 , n25080 );
and ( n25082 , n24063 , n24064 );
and ( n25083 , n24064 , n24066 );
and ( n25084 , n24063 , n24066 );
or ( n25085 , n25082 , n25083 , n25084 );
and ( n25086 , n6187 , n4403 );
and ( n25087 , n6569 , n4102 );
xor ( n25088 , n25086 , n25087 );
and ( n25089 , n6816 , n3749 );
xor ( n25090 , n25088 , n25089 );
xor ( n25091 , n25085 , n25090 );
and ( n25092 , n5819 , n4730 );
buf ( n25093 , n25092 );
xor ( n25094 , n25091 , n25093 );
xor ( n25095 , n25081 , n25094 );
xor ( n25096 , n25061 , n25095 );
xor ( n25097 , n25031 , n25096 );
xor ( n25098 , n25022 , n25097 );
and ( n25099 , n24128 , n24166 );
and ( n25100 , n24166 , n24193 );
and ( n25101 , n24128 , n24193 );
or ( n25102 , n25099 , n25100 , n25101 );
and ( n25103 , n24089 , n24104 );
and ( n25104 , n24104 , n24121 );
and ( n25105 , n24089 , n24121 );
or ( n25106 , n25103 , n25104 , n25105 );
and ( n25107 , n24171 , n24175 );
and ( n25108 , n24175 , n24192 );
and ( n25109 , n24171 , n24192 );
or ( n25110 , n25107 , n25108 , n25109 );
xor ( n25111 , n25106 , n25110 );
and ( n25112 , n24093 , n24097 );
and ( n25113 , n24097 , n24103 );
and ( n25114 , n24093 , n24103 );
or ( n25115 , n25112 , n25113 , n25114 );
and ( n25116 , n24110 , n24111 );
and ( n25117 , n24111 , n24113 );
and ( n25118 , n24110 , n24113 );
or ( n25119 , n25116 , n25117 , n25118 );
and ( n25120 , n2462 , n9348 );
and ( n25121 , n2779 , n8669 );
xor ( n25122 , n25120 , n25121 );
and ( n25123 , n3024 , n8243 );
xor ( n25124 , n25122 , n25123 );
xor ( n25125 , n25119 , n25124 );
and ( n25126 , n3182 , n7662 );
and ( n25127 , n3545 , n7310 );
xor ( n25128 , n25126 , n25127 );
and ( n25129 , n3801 , n6971 );
xor ( n25130 , n25128 , n25129 );
xor ( n25131 , n25125 , n25130 );
xor ( n25132 , n25115 , n25131 );
and ( n25133 , n24099 , n24100 );
and ( n25134 , n24100 , n24102 );
and ( n25135 , n24099 , n24102 );
or ( n25136 , n25133 , n25134 , n25135 );
and ( n25137 , n24181 , n24182 );
and ( n25138 , n24182 , n24184 );
and ( n25139 , n24181 , n24184 );
or ( n25140 , n25137 , n25138 , n25139 );
xor ( n25141 , n25136 , n25140 );
and ( n25142 , n1933 , n11718 );
and ( n25143 , n2120 , n10977 );
xor ( n25144 , n25142 , n25143 );
and ( n25145 , n2324 , n10239 );
xor ( n25146 , n25144 , n25145 );
xor ( n25147 , n25141 , n25146 );
xor ( n25148 , n25132 , n25147 );
xor ( n25149 , n25111 , n25148 );
xor ( n25150 , n25102 , n25149 );
and ( n25151 , n24132 , n24149 );
and ( n25152 , n24149 , n24165 );
and ( n25153 , n24132 , n24165 );
or ( n25154 , n25151 , n25152 , n25153 );
and ( n25155 , n24136 , n24142 );
and ( n25156 , n24142 , n24148 );
and ( n25157 , n24136 , n24148 );
or ( n25158 , n25155 , n25156 , n25157 );
and ( n25159 , n24138 , n24139 );
and ( n25160 , n24139 , n24141 );
and ( n25161 , n24138 , n24141 );
or ( n25162 , n25159 , n25160 , n25161 );
buf ( n25163 , n415 );
and ( n25164 , n599 , n25163 );
and ( n25165 , n608 , n24137 );
xor ( n25166 , n25164 , n25165 );
and ( n25167 , n611 , n23075 );
xor ( n25168 , n25166 , n25167 );
xor ( n25169 , n25162 , n25168 );
and ( n25170 , n632 , n22065 );
and ( n25171 , n671 , n20976 );
xor ( n25172 , n25170 , n25171 );
and ( n25173 , n715 , n20156 );
xor ( n25174 , n25172 , n25173 );
xor ( n25175 , n25169 , n25174 );
xor ( n25176 , n25158 , n25175 );
and ( n25177 , n24160 , n24161 );
and ( n25178 , n24161 , n24163 );
and ( n25179 , n24160 , n24163 );
or ( n25180 , n25177 , n25178 , n25179 );
and ( n25181 , n24144 , n24145 );
and ( n25182 , n24145 , n24147 );
and ( n25183 , n24144 , n24147 );
or ( n25184 , n25181 , n25182 , n25183 );
xor ( n25185 , n25180 , n25184 );
and ( n25186 , n783 , n19222 );
and ( n25187 , n856 , n18407 );
xor ( n25188 , n25186 , n25187 );
and ( n25189 , n925 , n17422 );
xor ( n25190 , n25188 , n25189 );
xor ( n25191 , n25185 , n25190 );
xor ( n25192 , n25176 , n25191 );
xor ( n25193 , n25154 , n25192 );
and ( n25194 , n24154 , n24158 );
and ( n25195 , n24158 , n24164 );
and ( n25196 , n24154 , n24164 );
or ( n25197 , n25194 , n25195 , n25196 );
and ( n25198 , n24180 , n24185 );
and ( n25199 , n24185 , n24191 );
and ( n25200 , n24180 , n24191 );
or ( n25201 , n25198 , n25199 , n25200 );
xor ( n25202 , n25197 , n25201 );
and ( n25203 , n24187 , n24188 );
and ( n25204 , n24188 , n24190 );
and ( n25205 , n24187 , n24190 );
or ( n25206 , n25203 , n25204 , n25205 );
and ( n25207 , n1047 , n16550 );
and ( n25208 , n1164 , n15691 );
xor ( n25209 , n25207 , n25208 );
and ( n25210 , n1287 , n14838 );
xor ( n25211 , n25209 , n25210 );
xor ( n25212 , n25206 , n25211 );
and ( n25213 , n1383 , n14044 );
and ( n25214 , n1580 , n13256 );
xor ( n25215 , n25213 , n25214 );
and ( n25216 , n1694 , n12531 );
xor ( n25217 , n25215 , n25216 );
xor ( n25218 , n25212 , n25217 );
xor ( n25219 , n25202 , n25218 );
xor ( n25220 , n25193 , n25219 );
xor ( n25221 , n25150 , n25220 );
xor ( n25222 , n25098 , n25221 );
xor ( n25223 , n25018 , n25222 );
xor ( n25224 , n24893 , n25223 );
and ( n25225 , n23872 , n23876 );
and ( n25226 , n23876 , n23987 );
and ( n25227 , n23872 , n23987 );
or ( n25228 , n25225 , n25226 , n25227 );
and ( n25229 , n24205 , n24217 );
xor ( n25230 , n25228 , n25229 );
and ( n25231 , n24209 , n24216 );
and ( n25232 , n23885 , n23910 );
and ( n25233 , n23910 , n23948 );
and ( n25234 , n23885 , n23948 );
or ( n25235 , n25232 , n25233 , n25234 );
and ( n25236 , n24213 , n24215 );
xor ( n25237 , n25235 , n25236 );
and ( n25238 , n23889 , n23893 );
and ( n25239 , n23893 , n23909 );
and ( n25240 , n23889 , n23909 );
or ( n25241 , n25238 , n25239 , n25240 );
and ( n25242 , n24214 , n615 );
buf ( n25243 , n415 );
and ( n25244 , n25243 , n612 );
xor ( n25245 , n25242 , n25244 );
xor ( n25246 , n25241 , n25245 );
xor ( n25247 , n25237 , n25246 );
xor ( n25248 , n25231 , n25247 );
xor ( n25249 , n25230 , n25248 );
xor ( n25250 , n25224 , n25249 );
xor ( n25251 , n24889 , n25250 );
and ( n25252 , n23855 , n23859 );
and ( n25253 , n23859 , n24220 );
and ( n25254 , n23855 , n24220 );
or ( n25255 , n25252 , n25253 , n25254 );
xor ( n25256 , n25251 , n25255 );
and ( n25257 , n24221 , n24225 );
and ( n25258 , n24226 , n24229 );
or ( n25259 , n25257 , n25258 );
xor ( n25260 , n25256 , n25259 );
buf ( n25261 , n25260 );
buf ( n25262 , n25261 );
not ( n25263 , n25262 );
nor ( n25264 , n25263 , n8739 );
xor ( n25265 , n24880 , n25264 );
and ( n25266 , n23851 , n24234 );
and ( n25267 , n24235 , n24238 );
or ( n25268 , n25266 , n25267 );
xor ( n25269 , n25265 , n25268 );
buf ( n25270 , n25269 );
buf ( n25271 , n25270 );
not ( n25272 , n25271 );
buf ( n25273 , n554 );
not ( n25274 , n25273 );
nor ( n25275 , n25272 , n25274 );
xor ( n25276 , n24562 , n25275 );
xor ( n25277 , n24250 , n24559 );
nor ( n25278 , n24242 , n25274 );
and ( n25279 , n25277 , n25278 );
xor ( n25280 , n25277 , n25278 );
xor ( n25281 , n24254 , n24557 );
nor ( n25282 , n23225 , n25274 );
and ( n25283 , n25281 , n25282 );
xor ( n25284 , n25281 , n25282 );
xor ( n25285 , n24258 , n24555 );
nor ( n25286 , n22231 , n25274 );
and ( n25287 , n25285 , n25286 );
xor ( n25288 , n25285 , n25286 );
xor ( n25289 , n24262 , n24553 );
nor ( n25290 , n21258 , n25274 );
and ( n25291 , n25289 , n25290 );
xor ( n25292 , n25289 , n25290 );
xor ( n25293 , n24266 , n24551 );
nor ( n25294 , n20303 , n25274 );
and ( n25295 , n25293 , n25294 );
xor ( n25296 , n25293 , n25294 );
xor ( n25297 , n24270 , n24549 );
nor ( n25298 , n19365 , n25274 );
and ( n25299 , n25297 , n25298 );
xor ( n25300 , n25297 , n25298 );
xor ( n25301 , n24274 , n24547 );
nor ( n25302 , n18448 , n25274 );
and ( n25303 , n25301 , n25302 );
xor ( n25304 , n25301 , n25302 );
xor ( n25305 , n24278 , n24545 );
nor ( n25306 , n17548 , n25274 );
and ( n25307 , n25305 , n25306 );
xor ( n25308 , n25305 , n25306 );
xor ( n25309 , n24282 , n24543 );
nor ( n25310 , n16669 , n25274 );
and ( n25311 , n25309 , n25310 );
xor ( n25312 , n25309 , n25310 );
xor ( n25313 , n24286 , n24541 );
nor ( n25314 , n15809 , n25274 );
and ( n25315 , n25313 , n25314 );
xor ( n25316 , n25313 , n25314 );
xor ( n25317 , n24290 , n24539 );
nor ( n25318 , n14968 , n25274 );
and ( n25319 , n25317 , n25318 );
xor ( n25320 , n25317 , n25318 );
xor ( n25321 , n24294 , n24537 );
nor ( n25322 , n14147 , n25274 );
and ( n25323 , n25321 , n25322 );
xor ( n25324 , n25321 , n25322 );
xor ( n25325 , n24298 , n24535 );
nor ( n25326 , n13349 , n25274 );
and ( n25327 , n25325 , n25326 );
xor ( n25328 , n25325 , n25326 );
xor ( n25329 , n24302 , n24533 );
nor ( n25330 , n12564 , n25274 );
and ( n25331 , n25329 , n25330 );
xor ( n25332 , n25329 , n25330 );
xor ( n25333 , n24306 , n24531 );
nor ( n25334 , n11799 , n25274 );
and ( n25335 , n25333 , n25334 );
xor ( n25336 , n25333 , n25334 );
xor ( n25337 , n24310 , n24529 );
nor ( n25338 , n11050 , n25274 );
and ( n25339 , n25337 , n25338 );
xor ( n25340 , n25337 , n25338 );
xor ( n25341 , n24314 , n24527 );
nor ( n25342 , n10321 , n25274 );
and ( n25343 , n25341 , n25342 );
xor ( n25344 , n25341 , n25342 );
xor ( n25345 , n24318 , n24525 );
nor ( n25346 , n9429 , n25274 );
and ( n25347 , n25345 , n25346 );
xor ( n25348 , n25345 , n25346 );
xor ( n25349 , n24322 , n24523 );
nor ( n25350 , n8949 , n25274 );
and ( n25351 , n25349 , n25350 );
xor ( n25352 , n25349 , n25350 );
xor ( n25353 , n24326 , n24521 );
nor ( n25354 , n9437 , n25274 );
and ( n25355 , n25353 , n25354 );
xor ( n25356 , n25353 , n25354 );
xor ( n25357 , n24330 , n24519 );
nor ( n25358 , n9446 , n25274 );
and ( n25359 , n25357 , n25358 );
xor ( n25360 , n25357 , n25358 );
xor ( n25361 , n24334 , n24517 );
nor ( n25362 , n9455 , n25274 );
and ( n25363 , n25361 , n25362 );
xor ( n25364 , n25361 , n25362 );
xor ( n25365 , n24338 , n24515 );
nor ( n25366 , n9464 , n25274 );
and ( n25367 , n25365 , n25366 );
xor ( n25368 , n25365 , n25366 );
xor ( n25369 , n24342 , n24513 );
nor ( n25370 , n9473 , n25274 );
and ( n25371 , n25369 , n25370 );
xor ( n25372 , n25369 , n25370 );
xor ( n25373 , n24346 , n24511 );
nor ( n25374 , n9482 , n25274 );
and ( n25375 , n25373 , n25374 );
xor ( n25376 , n25373 , n25374 );
xor ( n25377 , n24350 , n24509 );
nor ( n25378 , n9491 , n25274 );
and ( n25379 , n25377 , n25378 );
xor ( n25380 , n25377 , n25378 );
xor ( n25381 , n24354 , n24507 );
nor ( n25382 , n9500 , n25274 );
and ( n25383 , n25381 , n25382 );
xor ( n25384 , n25381 , n25382 );
xor ( n25385 , n24358 , n24505 );
nor ( n25386 , n9509 , n25274 );
and ( n25387 , n25385 , n25386 );
xor ( n25388 , n25385 , n25386 );
xor ( n25389 , n24362 , n24503 );
nor ( n25390 , n9518 , n25274 );
and ( n25391 , n25389 , n25390 );
xor ( n25392 , n25389 , n25390 );
xor ( n25393 , n24366 , n24501 );
nor ( n25394 , n9527 , n25274 );
and ( n25395 , n25393 , n25394 );
xor ( n25396 , n25393 , n25394 );
xor ( n25397 , n24370 , n24499 );
nor ( n25398 , n9536 , n25274 );
and ( n25399 , n25397 , n25398 );
xor ( n25400 , n25397 , n25398 );
xor ( n25401 , n24374 , n24497 );
nor ( n25402 , n9545 , n25274 );
and ( n25403 , n25401 , n25402 );
xor ( n25404 , n25401 , n25402 );
xor ( n25405 , n24378 , n24495 );
nor ( n25406 , n9554 , n25274 );
and ( n25407 , n25405 , n25406 );
xor ( n25408 , n25405 , n25406 );
xor ( n25409 , n24382 , n24493 );
nor ( n25410 , n9563 , n25274 );
and ( n25411 , n25409 , n25410 );
xor ( n25412 , n25409 , n25410 );
xor ( n25413 , n24386 , n24491 );
nor ( n25414 , n9572 , n25274 );
and ( n25415 , n25413 , n25414 );
xor ( n25416 , n25413 , n25414 );
xor ( n25417 , n24390 , n24489 );
nor ( n25418 , n9581 , n25274 );
and ( n25419 , n25417 , n25418 );
xor ( n25420 , n25417 , n25418 );
xor ( n25421 , n24394 , n24487 );
nor ( n25422 , n9590 , n25274 );
and ( n25423 , n25421 , n25422 );
xor ( n25424 , n25421 , n25422 );
xor ( n25425 , n24398 , n24485 );
nor ( n25426 , n9599 , n25274 );
and ( n25427 , n25425 , n25426 );
xor ( n25428 , n25425 , n25426 );
xor ( n25429 , n24402 , n24483 );
nor ( n25430 , n9608 , n25274 );
and ( n25431 , n25429 , n25430 );
xor ( n25432 , n25429 , n25430 );
xor ( n25433 , n24406 , n24481 );
nor ( n25434 , n9617 , n25274 );
and ( n25435 , n25433 , n25434 );
xor ( n25436 , n25433 , n25434 );
xor ( n25437 , n24410 , n24479 );
nor ( n25438 , n9626 , n25274 );
and ( n25439 , n25437 , n25438 );
xor ( n25440 , n25437 , n25438 );
xor ( n25441 , n24414 , n24477 );
nor ( n25442 , n9635 , n25274 );
and ( n25443 , n25441 , n25442 );
xor ( n25444 , n25441 , n25442 );
xor ( n25445 , n24418 , n24475 );
nor ( n25446 , n9644 , n25274 );
and ( n25447 , n25445 , n25446 );
xor ( n25448 , n25445 , n25446 );
xor ( n25449 , n24422 , n24473 );
nor ( n25450 , n9653 , n25274 );
and ( n25451 , n25449 , n25450 );
xor ( n25452 , n25449 , n25450 );
xor ( n25453 , n24426 , n24471 );
nor ( n25454 , n9662 , n25274 );
and ( n25455 , n25453 , n25454 );
xor ( n25456 , n25453 , n25454 );
xor ( n25457 , n24430 , n24469 );
nor ( n25458 , n9671 , n25274 );
and ( n25459 , n25457 , n25458 );
xor ( n25460 , n25457 , n25458 );
xor ( n25461 , n24434 , n24467 );
nor ( n25462 , n9680 , n25274 );
and ( n25463 , n25461 , n25462 );
xor ( n25464 , n25461 , n25462 );
xor ( n25465 , n24438 , n24465 );
nor ( n25466 , n9689 , n25274 );
and ( n25467 , n25465 , n25466 );
xor ( n25468 , n25465 , n25466 );
xor ( n25469 , n24442 , n24463 );
nor ( n25470 , n9698 , n25274 );
and ( n25471 , n25469 , n25470 );
xor ( n25472 , n25469 , n25470 );
xor ( n25473 , n24446 , n24461 );
nor ( n25474 , n9707 , n25274 );
and ( n25475 , n25473 , n25474 );
xor ( n25476 , n25473 , n25474 );
xor ( n25477 , n24450 , n24459 );
nor ( n25478 , n9716 , n25274 );
and ( n25479 , n25477 , n25478 );
xor ( n25480 , n25477 , n25478 );
xor ( n25481 , n24454 , n24457 );
nor ( n25482 , n9725 , n25274 );
and ( n25483 , n25481 , n25482 );
xor ( n25484 , n25481 , n25482 );
xor ( n25485 , n24455 , n24456 );
nor ( n25486 , n9734 , n25274 );
and ( n25487 , n25485 , n25486 );
xor ( n25488 , n25485 , n25486 );
nor ( n25489 , n9752 , n24244 );
nor ( n25490 , n9743 , n25274 );
and ( n25491 , n25489 , n25490 );
and ( n25492 , n25488 , n25491 );
or ( n25493 , n25487 , n25492 );
and ( n25494 , n25484 , n25493 );
or ( n25495 , n25483 , n25494 );
and ( n25496 , n25480 , n25495 );
or ( n25497 , n25479 , n25496 );
and ( n25498 , n25476 , n25497 );
or ( n25499 , n25475 , n25498 );
and ( n25500 , n25472 , n25499 );
or ( n25501 , n25471 , n25500 );
and ( n25502 , n25468 , n25501 );
or ( n25503 , n25467 , n25502 );
and ( n25504 , n25464 , n25503 );
or ( n25505 , n25463 , n25504 );
and ( n25506 , n25460 , n25505 );
or ( n25507 , n25459 , n25506 );
and ( n25508 , n25456 , n25507 );
or ( n25509 , n25455 , n25508 );
and ( n25510 , n25452 , n25509 );
or ( n25511 , n25451 , n25510 );
and ( n25512 , n25448 , n25511 );
or ( n25513 , n25447 , n25512 );
and ( n25514 , n25444 , n25513 );
or ( n25515 , n25443 , n25514 );
and ( n25516 , n25440 , n25515 );
or ( n25517 , n25439 , n25516 );
and ( n25518 , n25436 , n25517 );
or ( n25519 , n25435 , n25518 );
and ( n25520 , n25432 , n25519 );
or ( n25521 , n25431 , n25520 );
and ( n25522 , n25428 , n25521 );
or ( n25523 , n25427 , n25522 );
and ( n25524 , n25424 , n25523 );
or ( n25525 , n25423 , n25524 );
and ( n25526 , n25420 , n25525 );
or ( n25527 , n25419 , n25526 );
and ( n25528 , n25416 , n25527 );
or ( n25529 , n25415 , n25528 );
and ( n25530 , n25412 , n25529 );
or ( n25531 , n25411 , n25530 );
and ( n25532 , n25408 , n25531 );
or ( n25533 , n25407 , n25532 );
and ( n25534 , n25404 , n25533 );
or ( n25535 , n25403 , n25534 );
and ( n25536 , n25400 , n25535 );
or ( n25537 , n25399 , n25536 );
and ( n25538 , n25396 , n25537 );
or ( n25539 , n25395 , n25538 );
and ( n25540 , n25392 , n25539 );
or ( n25541 , n25391 , n25540 );
and ( n25542 , n25388 , n25541 );
or ( n25543 , n25387 , n25542 );
and ( n25544 , n25384 , n25543 );
or ( n25545 , n25383 , n25544 );
and ( n25546 , n25380 , n25545 );
or ( n25547 , n25379 , n25546 );
and ( n25548 , n25376 , n25547 );
or ( n25549 , n25375 , n25548 );
and ( n25550 , n25372 , n25549 );
or ( n25551 , n25371 , n25550 );
and ( n25552 , n25368 , n25551 );
or ( n25553 , n25367 , n25552 );
and ( n25554 , n25364 , n25553 );
or ( n25555 , n25363 , n25554 );
and ( n25556 , n25360 , n25555 );
or ( n25557 , n25359 , n25556 );
and ( n25558 , n25356 , n25557 );
or ( n25559 , n25355 , n25558 );
and ( n25560 , n25352 , n25559 );
or ( n25561 , n25351 , n25560 );
and ( n25562 , n25348 , n25561 );
or ( n25563 , n25347 , n25562 );
and ( n25564 , n25344 , n25563 );
or ( n25565 , n25343 , n25564 );
and ( n25566 , n25340 , n25565 );
or ( n25567 , n25339 , n25566 );
and ( n25568 , n25336 , n25567 );
or ( n25569 , n25335 , n25568 );
and ( n25570 , n25332 , n25569 );
or ( n25571 , n25331 , n25570 );
and ( n25572 , n25328 , n25571 );
or ( n25573 , n25327 , n25572 );
and ( n25574 , n25324 , n25573 );
or ( n25575 , n25323 , n25574 );
and ( n25576 , n25320 , n25575 );
or ( n25577 , n25319 , n25576 );
and ( n25578 , n25316 , n25577 );
or ( n25579 , n25315 , n25578 );
and ( n25580 , n25312 , n25579 );
or ( n25581 , n25311 , n25580 );
and ( n25582 , n25308 , n25581 );
or ( n25583 , n25307 , n25582 );
and ( n25584 , n25304 , n25583 );
or ( n25585 , n25303 , n25584 );
and ( n25586 , n25300 , n25585 );
or ( n25587 , n25299 , n25586 );
and ( n25588 , n25296 , n25587 );
or ( n25589 , n25295 , n25588 );
and ( n25590 , n25292 , n25589 );
or ( n25591 , n25291 , n25590 );
and ( n25592 , n25288 , n25591 );
or ( n25593 , n25287 , n25592 );
and ( n25594 , n25284 , n25593 );
or ( n25595 , n25283 , n25594 );
and ( n25596 , n25280 , n25595 );
or ( n25597 , n25279 , n25596 );
xor ( n25598 , n25276 , n25597 );
buf ( n25599 , n478 );
not ( n25600 , n25599 );
nor ( n25601 , n601 , n25600 );
buf ( n25602 , n25601 );
nor ( n25603 , n622 , n23541 );
xor ( n25604 , n25602 , n25603 );
buf ( n25605 , n25604 );
nor ( n25606 , n646 , n22541 );
xor ( n25607 , n25605 , n25606 );
and ( n25608 , n24566 , n24567 );
buf ( n25609 , n25608 );
xor ( n25610 , n25607 , n25609 );
nor ( n25611 , n684 , n21562 );
xor ( n25612 , n25610 , n25611 );
and ( n25613 , n24569 , n24570 );
and ( n25614 , n24571 , n24573 );
or ( n25615 , n25613 , n25614 );
xor ( n25616 , n25612 , n25615 );
nor ( n25617 , n733 , n20601 );
xor ( n25618 , n25616 , n25617 );
and ( n25619 , n24574 , n24575 );
and ( n25620 , n24576 , n24579 );
or ( n25621 , n25619 , n25620 );
xor ( n25622 , n25618 , n25621 );
nor ( n25623 , n796 , n19657 );
xor ( n25624 , n25622 , n25623 );
and ( n25625 , n24580 , n24581 );
and ( n25626 , n24582 , n24585 );
or ( n25627 , n25625 , n25626 );
xor ( n25628 , n25624 , n25627 );
nor ( n25629 , n868 , n18734 );
xor ( n25630 , n25628 , n25629 );
and ( n25631 , n24586 , n24587 );
and ( n25632 , n24588 , n24591 );
or ( n25633 , n25631 , n25632 );
xor ( n25634 , n25630 , n25633 );
nor ( n25635 , n958 , n17828 );
xor ( n25636 , n25634 , n25635 );
and ( n25637 , n24592 , n24593 );
and ( n25638 , n24594 , n24597 );
or ( n25639 , n25637 , n25638 );
xor ( n25640 , n25636 , n25639 );
nor ( n25641 , n1062 , n16943 );
xor ( n25642 , n25640 , n25641 );
and ( n25643 , n24598 , n24599 );
and ( n25644 , n24600 , n24603 );
or ( n25645 , n25643 , n25644 );
xor ( n25646 , n25642 , n25645 );
nor ( n25647 , n1176 , n16077 );
xor ( n25648 , n25646 , n25647 );
and ( n25649 , n24604 , n24605 );
and ( n25650 , n24606 , n24609 );
or ( n25651 , n25649 , n25650 );
xor ( n25652 , n25648 , n25651 );
nor ( n25653 , n1303 , n15230 );
xor ( n25654 , n25652 , n25653 );
and ( n25655 , n24610 , n24611 );
and ( n25656 , n24612 , n24615 );
or ( n25657 , n25655 , n25656 );
xor ( n25658 , n25654 , n25657 );
nor ( n25659 , n1445 , n14403 );
xor ( n25660 , n25658 , n25659 );
and ( n25661 , n24616 , n24617 );
and ( n25662 , n24618 , n24621 );
or ( n25663 , n25661 , n25662 );
xor ( n25664 , n25660 , n25663 );
nor ( n25665 , n1598 , n13599 );
xor ( n25666 , n25664 , n25665 );
and ( n25667 , n24622 , n24623 );
and ( n25668 , n24624 , n24627 );
or ( n25669 , n25667 , n25668 );
xor ( n25670 , n25666 , n25669 );
nor ( n25671 , n1766 , n12808 );
xor ( n25672 , n25670 , n25671 );
and ( n25673 , n24628 , n24629 );
and ( n25674 , n24630 , n24633 );
or ( n25675 , n25673 , n25674 );
xor ( n25676 , n25672 , n25675 );
nor ( n25677 , n1945 , n12037 );
xor ( n25678 , n25676 , n25677 );
and ( n25679 , n24634 , n24635 );
and ( n25680 , n24636 , n24639 );
or ( n25681 , n25679 , n25680 );
xor ( n25682 , n25678 , n25681 );
nor ( n25683 , n2137 , n11282 );
xor ( n25684 , n25682 , n25683 );
and ( n25685 , n24640 , n24641 );
and ( n25686 , n24642 , n24645 );
or ( n25687 , n25685 , n25686 );
xor ( n25688 , n25684 , n25687 );
nor ( n25689 , n2343 , n10547 );
xor ( n25690 , n25688 , n25689 );
and ( n25691 , n24646 , n24647 );
and ( n25692 , n24648 , n24651 );
or ( n25693 , n25691 , n25692 );
xor ( n25694 , n25690 , n25693 );
nor ( n25695 , n2566 , n9829 );
xor ( n25696 , n25694 , n25695 );
and ( n25697 , n24652 , n24653 );
and ( n25698 , n24654 , n24657 );
or ( n25699 , n25697 , n25698 );
xor ( n25700 , n25696 , n25699 );
nor ( n25701 , n2797 , n8955 );
xor ( n25702 , n25700 , n25701 );
and ( n25703 , n24658 , n24659 );
and ( n25704 , n24660 , n24663 );
or ( n25705 , n25703 , n25704 );
xor ( n25706 , n25702 , n25705 );
nor ( n25707 , n3043 , n603 );
xor ( n25708 , n25706 , n25707 );
and ( n25709 , n24664 , n24665 );
and ( n25710 , n24666 , n24669 );
or ( n25711 , n25709 , n25710 );
xor ( n25712 , n25708 , n25711 );
nor ( n25713 , n3300 , n652 );
xor ( n25714 , n25712 , n25713 );
and ( n25715 , n24670 , n24671 );
and ( n25716 , n24672 , n24675 );
or ( n25717 , n25715 , n25716 );
xor ( n25718 , n25714 , n25717 );
nor ( n25719 , n3570 , n624 );
xor ( n25720 , n25718 , n25719 );
and ( n25721 , n24676 , n24677 );
and ( n25722 , n24678 , n24681 );
or ( n25723 , n25721 , n25722 );
xor ( n25724 , n25720 , n25723 );
nor ( n25725 , n3853 , n648 );
xor ( n25726 , n25724 , n25725 );
and ( n25727 , n24682 , n24683 );
and ( n25728 , n24684 , n24687 );
or ( n25729 , n25727 , n25728 );
xor ( n25730 , n25726 , n25729 );
nor ( n25731 , n4151 , n686 );
xor ( n25732 , n25730 , n25731 );
and ( n25733 , n24688 , n24689 );
and ( n25734 , n24690 , n24693 );
or ( n25735 , n25733 , n25734 );
xor ( n25736 , n25732 , n25735 );
nor ( n25737 , n4458 , n735 );
xor ( n25738 , n25736 , n25737 );
and ( n25739 , n24694 , n24695 );
and ( n25740 , n24696 , n24699 );
or ( n25741 , n25739 , n25740 );
xor ( n25742 , n25738 , n25741 );
nor ( n25743 , n4786 , n798 );
xor ( n25744 , n25742 , n25743 );
and ( n25745 , n24700 , n24701 );
and ( n25746 , n24702 , n24705 );
or ( n25747 , n25745 , n25746 );
xor ( n25748 , n25744 , n25747 );
nor ( n25749 , n5126 , n870 );
xor ( n25750 , n25748 , n25749 );
and ( n25751 , n24706 , n24707 );
and ( n25752 , n24708 , n24711 );
or ( n25753 , n25751 , n25752 );
xor ( n25754 , n25750 , n25753 );
nor ( n25755 , n5477 , n960 );
xor ( n25756 , n25754 , n25755 );
and ( n25757 , n24712 , n24713 );
and ( n25758 , n24714 , n24717 );
or ( n25759 , n25757 , n25758 );
xor ( n25760 , n25756 , n25759 );
nor ( n25761 , n5838 , n1064 );
xor ( n25762 , n25760 , n25761 );
and ( n25763 , n24718 , n24719 );
and ( n25764 , n24720 , n24723 );
or ( n25765 , n25763 , n25764 );
xor ( n25766 , n25762 , n25765 );
nor ( n25767 , n6212 , n1178 );
xor ( n25768 , n25766 , n25767 );
and ( n25769 , n24724 , n24725 );
and ( n25770 , n24726 , n24729 );
or ( n25771 , n25769 , n25770 );
xor ( n25772 , n25768 , n25771 );
nor ( n25773 , n6596 , n1305 );
xor ( n25774 , n25772 , n25773 );
and ( n25775 , n24730 , n24731 );
and ( n25776 , n24732 , n24735 );
or ( n25777 , n25775 , n25776 );
xor ( n25778 , n25774 , n25777 );
nor ( n25779 , n6997 , n1447 );
xor ( n25780 , n25778 , n25779 );
and ( n25781 , n24736 , n24737 );
and ( n25782 , n24738 , n24741 );
or ( n25783 , n25781 , n25782 );
xor ( n25784 , n25780 , n25783 );
nor ( n25785 , n7413 , n1600 );
xor ( n25786 , n25784 , n25785 );
and ( n25787 , n24742 , n24743 );
and ( n25788 , n24744 , n24747 );
or ( n25789 , n25787 , n25788 );
xor ( n25790 , n25786 , n25789 );
nor ( n25791 , n7841 , n1768 );
xor ( n25792 , n25790 , n25791 );
and ( n25793 , n24748 , n24749 );
and ( n25794 , n24750 , n24753 );
or ( n25795 , n25793 , n25794 );
xor ( n25796 , n25792 , n25795 );
nor ( n25797 , n8281 , n1947 );
xor ( n25798 , n25796 , n25797 );
and ( n25799 , n24754 , n24755 );
and ( n25800 , n24756 , n24759 );
or ( n25801 , n25799 , n25800 );
xor ( n25802 , n25798 , n25801 );
nor ( n25803 , n8737 , n2139 );
xor ( n25804 , n25802 , n25803 );
and ( n25805 , n24760 , n24761 );
and ( n25806 , n24762 , n24765 );
or ( n25807 , n25805 , n25806 );
xor ( n25808 , n25804 , n25807 );
nor ( n25809 , n9420 , n2345 );
xor ( n25810 , n25808 , n25809 );
and ( n25811 , n24766 , n24767 );
and ( n25812 , n24768 , n24771 );
or ( n25813 , n25811 , n25812 );
xor ( n25814 , n25810 , n25813 );
nor ( n25815 , n10312 , n2568 );
xor ( n25816 , n25814 , n25815 );
and ( n25817 , n24772 , n24773 );
and ( n25818 , n24774 , n24777 );
or ( n25819 , n25817 , n25818 );
xor ( n25820 , n25816 , n25819 );
nor ( n25821 , n11041 , n2799 );
xor ( n25822 , n25820 , n25821 );
and ( n25823 , n24778 , n24779 );
and ( n25824 , n24780 , n24783 );
or ( n25825 , n25823 , n25824 );
xor ( n25826 , n25822 , n25825 );
nor ( n25827 , n11790 , n3045 );
xor ( n25828 , n25826 , n25827 );
and ( n25829 , n24784 , n24785 );
and ( n25830 , n24786 , n24789 );
or ( n25831 , n25829 , n25830 );
xor ( n25832 , n25828 , n25831 );
nor ( n25833 , n12555 , n3302 );
xor ( n25834 , n25832 , n25833 );
and ( n25835 , n24790 , n24791 );
and ( n25836 , n24792 , n24795 );
or ( n25837 , n25835 , n25836 );
xor ( n25838 , n25834 , n25837 );
nor ( n25839 , n13340 , n3572 );
xor ( n25840 , n25838 , n25839 );
and ( n25841 , n24796 , n24797 );
and ( n25842 , n24798 , n24801 );
or ( n25843 , n25841 , n25842 );
xor ( n25844 , n25840 , n25843 );
nor ( n25845 , n14138 , n3855 );
xor ( n25846 , n25844 , n25845 );
and ( n25847 , n24802 , n24803 );
and ( n25848 , n24804 , n24807 );
or ( n25849 , n25847 , n25848 );
xor ( n25850 , n25846 , n25849 );
nor ( n25851 , n14959 , n4153 );
xor ( n25852 , n25850 , n25851 );
and ( n25853 , n24808 , n24809 );
and ( n25854 , n24810 , n24813 );
or ( n25855 , n25853 , n25854 );
xor ( n25856 , n25852 , n25855 );
nor ( n25857 , n15800 , n4460 );
xor ( n25858 , n25856 , n25857 );
and ( n25859 , n24814 , n24815 );
and ( n25860 , n24816 , n24819 );
or ( n25861 , n25859 , n25860 );
xor ( n25862 , n25858 , n25861 );
nor ( n25863 , n16660 , n4788 );
xor ( n25864 , n25862 , n25863 );
and ( n25865 , n24820 , n24821 );
and ( n25866 , n24822 , n24825 );
or ( n25867 , n25865 , n25866 );
xor ( n25868 , n25864 , n25867 );
nor ( n25869 , n17539 , n5128 );
xor ( n25870 , n25868 , n25869 );
and ( n25871 , n24826 , n24827 );
and ( n25872 , n24828 , n24831 );
or ( n25873 , n25871 , n25872 );
xor ( n25874 , n25870 , n25873 );
nor ( n25875 , n18439 , n5479 );
xor ( n25876 , n25874 , n25875 );
and ( n25877 , n24832 , n24833 );
and ( n25878 , n24834 , n24837 );
or ( n25879 , n25877 , n25878 );
xor ( n25880 , n25876 , n25879 );
nor ( n25881 , n19356 , n5840 );
xor ( n25882 , n25880 , n25881 );
and ( n25883 , n24838 , n24839 );
and ( n25884 , n24840 , n24843 );
or ( n25885 , n25883 , n25884 );
xor ( n25886 , n25882 , n25885 );
nor ( n25887 , n20294 , n6214 );
xor ( n25888 , n25886 , n25887 );
and ( n25889 , n24844 , n24845 );
and ( n25890 , n24846 , n24849 );
or ( n25891 , n25889 , n25890 );
xor ( n25892 , n25888 , n25891 );
nor ( n25893 , n21249 , n6598 );
xor ( n25894 , n25892 , n25893 );
and ( n25895 , n24850 , n24851 );
and ( n25896 , n24852 , n24855 );
or ( n25897 , n25895 , n25896 );
xor ( n25898 , n25894 , n25897 );
nor ( n25899 , n22222 , n6999 );
xor ( n25900 , n25898 , n25899 );
and ( n25901 , n24856 , n24857 );
and ( n25902 , n24858 , n24861 );
or ( n25903 , n25901 , n25902 );
xor ( n25904 , n25900 , n25903 );
nor ( n25905 , n23216 , n7415 );
xor ( n25906 , n25904 , n25905 );
and ( n25907 , n24862 , n24863 );
and ( n25908 , n24864 , n24867 );
or ( n25909 , n25907 , n25908 );
xor ( n25910 , n25906 , n25909 );
nor ( n25911 , n24233 , n7843 );
xor ( n25912 , n25910 , n25911 );
and ( n25913 , n24868 , n24869 );
and ( n25914 , n24870 , n24873 );
or ( n25915 , n25913 , n25914 );
xor ( n25916 , n25912 , n25915 );
nor ( n25917 , n25263 , n8283 );
xor ( n25918 , n25916 , n25917 );
and ( n25919 , n24874 , n24875 );
and ( n25920 , n24876 , n24879 );
or ( n25921 , n25919 , n25920 );
xor ( n25922 , n25918 , n25921 );
and ( n25923 , n25228 , n25229 );
and ( n25924 , n25229 , n25248 );
and ( n25925 , n25228 , n25248 );
or ( n25926 , n25923 , n25924 , n25925 );
and ( n25927 , n24893 , n25223 );
and ( n25928 , n25223 , n25249 );
and ( n25929 , n24893 , n25249 );
or ( n25930 , n25927 , n25928 , n25929 );
xor ( n25931 , n25926 , n25930 );
and ( n25932 , n24897 , n25017 );
and ( n25933 , n25017 , n25222 );
and ( n25934 , n24897 , n25222 );
or ( n25935 , n25932 , n25933 , n25934 );
and ( n25936 , n25022 , n25097 );
and ( n25937 , n25097 , n25221 );
and ( n25938 , n25022 , n25221 );
or ( n25939 , n25936 , n25937 , n25938 );
and ( n25940 , n24910 , n24978 );
and ( n25941 , n24978 , n25015 );
and ( n25942 , n24910 , n25015 );
or ( n25943 , n25940 , n25941 , n25942 );
and ( n25944 , n25026 , n25030 );
and ( n25945 , n25030 , n25096 );
and ( n25946 , n25026 , n25096 );
or ( n25947 , n25944 , n25945 , n25946 );
xor ( n25948 , n25943 , n25947 );
and ( n25949 , n24983 , n24987 );
and ( n25950 , n24987 , n25014 );
and ( n25951 , n24983 , n25014 );
or ( n25952 , n25949 , n25950 , n25951 );
and ( n25953 , n24944 , n24960 );
and ( n25954 , n24960 , n24976 );
and ( n25955 , n24944 , n24976 );
or ( n25956 , n25953 , n25954 , n25955 );
and ( n25957 , n24927 , n24931 );
and ( n25958 , n24931 , n24937 );
and ( n25959 , n24927 , n24937 );
or ( n25960 , n25957 , n25958 , n25959 );
and ( n25961 , n24948 , n24953 );
and ( n25962 , n24953 , n24959 );
and ( n25963 , n24948 , n24959 );
or ( n25964 , n25961 , n25962 , n25963 );
xor ( n25965 , n25960 , n25964 );
and ( n25966 , n24933 , n24934 );
and ( n25967 , n24934 , n24936 );
and ( n25968 , n24933 , n24936 );
or ( n25969 , n25966 , n25967 , n25968 );
and ( n25970 , n24949 , n24950 );
and ( n25971 , n24950 , n24952 );
and ( n25972 , n24949 , n24952 );
or ( n25973 , n25970 , n25971 , n25972 );
xor ( n25974 , n25969 , n25973 );
and ( n25975 , n21216 , n719 );
and ( n25976 , n22186 , n663 );
xor ( n25977 , n25975 , n25976 );
and ( n25978 , n22892 , n635 );
xor ( n25979 , n25977 , n25978 );
xor ( n25980 , n25974 , n25979 );
xor ( n25981 , n25965 , n25980 );
xor ( n25982 , n25956 , n25981 );
and ( n25983 , n24965 , n24969 );
and ( n25984 , n24969 , n24975 );
and ( n25985 , n24965 , n24975 );
or ( n25986 , n25983 , n25984 , n25985 );
and ( n25987 , n24955 , n24956 );
and ( n25988 , n24956 , n24958 );
and ( n25989 , n24955 , n24958 );
or ( n25990 , n25987 , n25988 , n25989 );
and ( n25991 , n18144 , n940 );
and ( n25992 , n19324 , n840 );
xor ( n25993 , n25991 , n25992 );
and ( n25994 , n20233 , n771 );
xor ( n25995 , n25993 , n25994 );
xor ( n25996 , n25990 , n25995 );
and ( n25997 , n15758 , n1254 );
and ( n25998 , n16637 , n1134 );
xor ( n25999 , n25997 , n25998 );
and ( n26000 , n17512 , n1034 );
xor ( n26001 , n25999 , n26000 );
xor ( n26002 , n25996 , n26001 );
xor ( n26003 , n25986 , n26002 );
and ( n26004 , n24971 , n24972 );
and ( n26005 , n24972 , n24974 );
and ( n26006 , n24971 , n24974 );
or ( n26007 , n26004 , n26005 , n26006 );
and ( n26008 , n25002 , n25003 );
and ( n26009 , n25003 , n25005 );
and ( n26010 , n25002 , n25005 );
or ( n26011 , n26008 , n26009 , n26010 );
xor ( n26012 , n26007 , n26011 );
and ( n26013 , n13322 , n1738 );
and ( n26014 , n14118 , n1551 );
xor ( n26015 , n26013 , n26014 );
and ( n26016 , n14938 , n1424 );
xor ( n26017 , n26015 , n26016 );
xor ( n26018 , n26012 , n26017 );
xor ( n26019 , n26003 , n26018 );
xor ( n26020 , n25982 , n26019 );
xor ( n26021 , n25952 , n26020 );
and ( n26022 , n24992 , n24996 );
and ( n26023 , n24996 , n25013 );
and ( n26024 , n24992 , n25013 );
or ( n26025 , n26022 , n26023 , n26024 );
and ( n26026 , n25065 , n25080 );
and ( n26027 , n25080 , n25094 );
and ( n26028 , n25065 , n25094 );
or ( n26029 , n26026 , n26027 , n26028 );
xor ( n26030 , n26025 , n26029 );
and ( n26031 , n25001 , n25006 );
and ( n26032 , n25006 , n25012 );
and ( n26033 , n25001 , n25012 );
or ( n26034 , n26031 , n26032 , n26033 );
and ( n26035 , n25069 , n25073 );
and ( n26036 , n25073 , n25079 );
and ( n26037 , n25069 , n25079 );
or ( n26038 , n26035 , n26036 , n26037 );
xor ( n26039 , n26034 , n26038 );
and ( n26040 , n25008 , n25009 );
and ( n26041 , n25009 , n25011 );
and ( n26042 , n25008 , n25011 );
or ( n26043 , n26040 , n26041 , n26042 );
and ( n26044 , n11015 , n2298 );
and ( n26045 , n11769 , n2100 );
xor ( n26046 , n26044 , n26045 );
and ( n26047 , n12320 , n1882 );
xor ( n26048 , n26046 , n26047 );
xor ( n26049 , n26043 , n26048 );
and ( n26050 , n8718 , n2981 );
and ( n26051 , n9400 , n2739 );
xor ( n26052 , n26050 , n26051 );
and ( n26053 , n10291 , n2544 );
xor ( n26054 , n26052 , n26053 );
xor ( n26055 , n26049 , n26054 );
xor ( n26056 , n26039 , n26055 );
xor ( n26057 , n26030 , n26056 );
xor ( n26058 , n26021 , n26057 );
xor ( n26059 , n25948 , n26058 );
xor ( n26060 , n25939 , n26059 );
and ( n26061 , n25102 , n25149 );
and ( n26062 , n25149 , n25220 );
and ( n26063 , n25102 , n25220 );
or ( n26064 , n26061 , n26062 , n26063 );
and ( n26065 , n25035 , n25060 );
and ( n26066 , n25060 , n25095 );
and ( n26067 , n25035 , n25095 );
or ( n26068 , n26065 , n26066 , n26067 );
and ( n26069 , n25106 , n25110 );
and ( n26070 , n25110 , n25148 );
and ( n26071 , n25106 , n25148 );
or ( n26072 , n26069 , n26070 , n26071 );
xor ( n26073 , n26068 , n26072 );
and ( n26074 , n25039 , n25043 );
and ( n26075 , n25043 , n25059 );
and ( n26076 , n25039 , n25059 );
or ( n26077 , n26074 , n26075 , n26076 );
and ( n26078 , n25119 , n25124 );
and ( n26079 , n25124 , n25130 );
and ( n26080 , n25119 , n25130 );
or ( n26081 , n26078 , n26079 , n26080 );
and ( n26082 , n25048 , n25052 );
and ( n26083 , n25052 , n25058 );
and ( n26084 , n25048 , n25058 );
or ( n26085 , n26082 , n26083 , n26084 );
xor ( n26086 , n26081 , n26085 );
and ( n26087 , n25054 , n25055 );
and ( n26088 , n25055 , n25057 );
and ( n26089 , n25054 , n25057 );
or ( n26090 , n26087 , n26088 , n26089 );
and ( n26091 , n25126 , n25127 );
and ( n26092 , n25127 , n25129 );
and ( n26093 , n25126 , n25129 );
or ( n26094 , n26091 , n26092 , n26093 );
xor ( n26095 , n26090 , n26094 );
and ( n26096 , n4132 , n6971 );
and ( n26097 , n4438 , n6504 );
xor ( n26098 , n26096 , n26097 );
and ( n26099 , n4766 , n6132 );
xor ( n26100 , n26098 , n26099 );
xor ( n26101 , n26095 , n26100 );
xor ( n26102 , n26086 , n26101 );
xor ( n26103 , n26077 , n26102 );
and ( n26104 , n25085 , n25090 );
and ( n26105 , n25090 , n25093 );
and ( n26106 , n25085 , n25093 );
or ( n26107 , n26104 , n26105 , n26106 );
and ( n26108 , n25075 , n25076 );
and ( n26109 , n25076 , n25078 );
and ( n26110 , n25075 , n25078 );
or ( n26111 , n26108 , n26109 , n26110 );
and ( n26112 , n25086 , n25087 );
and ( n26113 , n25087 , n25089 );
and ( n26114 , n25086 , n25089 );
or ( n26115 , n26112 , n26113 , n26114 );
xor ( n26116 , n26111 , n26115 );
and ( n26117 , n7385 , n3749 );
and ( n26118 , n7808 , n3495 );
xor ( n26119 , n26117 , n26118 );
and ( n26120 , n8079 , n3271 );
xor ( n26121 , n26119 , n26120 );
xor ( n26122 , n26116 , n26121 );
xor ( n26123 , n26107 , n26122 );
and ( n26124 , n4959 , n5408 );
and ( n26125 , n5459 , n5103 );
and ( n26126 , n26124 , n26125 );
and ( n26127 , n26125 , n25092 );
and ( n26128 , n26124 , n25092 );
or ( n26129 , n26126 , n26127 , n26128 );
and ( n26130 , n6187 , n4730 );
and ( n26131 , n6569 , n4403 );
xor ( n26132 , n26130 , n26131 );
and ( n26133 , n6816 , n4102 );
xor ( n26134 , n26132 , n26133 );
xor ( n26135 , n26129 , n26134 );
and ( n26136 , n4959 , n5765 );
buf ( n26137 , n5459 );
xor ( n26138 , n26136 , n26137 );
and ( n26139 , n5819 , n5103 );
xor ( n26140 , n26138 , n26139 );
xor ( n26141 , n26135 , n26140 );
xor ( n26142 , n26123 , n26141 );
xor ( n26143 , n26103 , n26142 );
xor ( n26144 , n26073 , n26143 );
xor ( n26145 , n26064 , n26144 );
and ( n26146 , n25154 , n25192 );
and ( n26147 , n25192 , n25219 );
and ( n26148 , n25154 , n25219 );
or ( n26149 , n26146 , n26147 , n26148 );
and ( n26150 , n25197 , n25201 );
and ( n26151 , n25201 , n25218 );
and ( n26152 , n25197 , n25218 );
or ( n26153 , n26150 , n26151 , n26152 );
and ( n26154 , n25115 , n25131 );
and ( n26155 , n25131 , n25147 );
and ( n26156 , n25115 , n25147 );
or ( n26157 , n26154 , n26155 , n26156 );
xor ( n26158 , n26153 , n26157 );
and ( n26159 , n25136 , n25140 );
and ( n26160 , n25140 , n25146 );
and ( n26161 , n25136 , n25146 );
or ( n26162 , n26159 , n26160 , n26161 );
and ( n26163 , n25120 , n25121 );
and ( n26164 , n25121 , n25123 );
and ( n26165 , n25120 , n25123 );
or ( n26166 , n26163 , n26164 , n26165 );
and ( n26167 , n3182 , n8243 );
and ( n26168 , n3545 , n7662 );
xor ( n26169 , n26167 , n26168 );
and ( n26170 , n3801 , n7310 );
xor ( n26171 , n26169 , n26170 );
xor ( n26172 , n26166 , n26171 );
and ( n26173 , n2462 , n10239 );
and ( n26174 , n2779 , n9348 );
xor ( n26175 , n26173 , n26174 );
and ( n26176 , n3024 , n8669 );
xor ( n26177 , n26175 , n26176 );
xor ( n26178 , n26172 , n26177 );
xor ( n26179 , n26162 , n26178 );
and ( n26180 , n25142 , n25143 );
and ( n26181 , n25143 , n25145 );
and ( n26182 , n25142 , n25145 );
or ( n26183 , n26180 , n26181 , n26182 );
and ( n26184 , n25213 , n25214 );
and ( n26185 , n25214 , n25216 );
and ( n26186 , n25213 , n25216 );
or ( n26187 , n26184 , n26185 , n26186 );
xor ( n26188 , n26183 , n26187 );
and ( n26189 , n1933 , n12531 );
and ( n26190 , n2120 , n11718 );
xor ( n26191 , n26189 , n26190 );
and ( n26192 , n2324 , n10977 );
xor ( n26193 , n26191 , n26192 );
xor ( n26194 , n26188 , n26193 );
xor ( n26195 , n26179 , n26194 );
xor ( n26196 , n26158 , n26195 );
xor ( n26197 , n26149 , n26196 );
and ( n26198 , n25158 , n25175 );
and ( n26199 , n25175 , n25191 );
and ( n26200 , n25158 , n25191 );
or ( n26201 , n26198 , n26199 , n26200 );
and ( n26202 , n25162 , n25168 );
and ( n26203 , n25168 , n25174 );
and ( n26204 , n25162 , n25174 );
or ( n26205 , n26202 , n26203 , n26204 );
and ( n26206 , n25164 , n25165 );
and ( n26207 , n25165 , n25167 );
and ( n26208 , n25164 , n25167 );
or ( n26209 , n26206 , n26207 , n26208 );
and ( n26210 , n632 , n23075 );
and ( n26211 , n671 , n22065 );
xor ( n26212 , n26210 , n26211 );
and ( n26213 , n715 , n20976 );
xor ( n26214 , n26212 , n26213 );
xor ( n26215 , n26209 , n26214 );
buf ( n26216 , n414 );
and ( n26217 , n599 , n26216 );
and ( n26218 , n608 , n25163 );
xor ( n26219 , n26217 , n26218 );
and ( n26220 , n611 , n24137 );
xor ( n26221 , n26219 , n26220 );
xor ( n26222 , n26215 , n26221 );
xor ( n26223 , n26205 , n26222 );
and ( n26224 , n25170 , n25171 );
and ( n26225 , n25171 , n25173 );
and ( n26226 , n25170 , n25173 );
or ( n26227 , n26224 , n26225 , n26226 );
and ( n26228 , n25186 , n25187 );
and ( n26229 , n25187 , n25189 );
and ( n26230 , n25186 , n25189 );
or ( n26231 , n26228 , n26229 , n26230 );
xor ( n26232 , n26227 , n26231 );
and ( n26233 , n783 , n20156 );
and ( n26234 , n856 , n19222 );
xor ( n26235 , n26233 , n26234 );
and ( n26236 , n925 , n18407 );
xor ( n26237 , n26235 , n26236 );
xor ( n26238 , n26232 , n26237 );
xor ( n26239 , n26223 , n26238 );
xor ( n26240 , n26201 , n26239 );
and ( n26241 , n25180 , n25184 );
and ( n26242 , n25184 , n25190 );
and ( n26243 , n25180 , n25190 );
or ( n26244 , n26241 , n26242 , n26243 );
and ( n26245 , n25206 , n25211 );
and ( n26246 , n25211 , n25217 );
and ( n26247 , n25206 , n25217 );
or ( n26248 , n26245 , n26246 , n26247 );
xor ( n26249 , n26244 , n26248 );
and ( n26250 , n25207 , n25208 );
and ( n26251 , n25208 , n25210 );
and ( n26252 , n25207 , n25210 );
or ( n26253 , n26250 , n26251 , n26252 );
and ( n26254 , n1383 , n14838 );
and ( n26255 , n1580 , n14044 );
xor ( n26256 , n26254 , n26255 );
and ( n26257 , n1694 , n13256 );
xor ( n26258 , n26256 , n26257 );
xor ( n26259 , n26253 , n26258 );
and ( n26260 , n1047 , n17422 );
and ( n26261 , n1164 , n16550 );
xor ( n26262 , n26260 , n26261 );
and ( n26263 , n1287 , n15691 );
xor ( n26264 , n26262 , n26263 );
xor ( n26265 , n26259 , n26264 );
xor ( n26266 , n26249 , n26265 );
xor ( n26267 , n26240 , n26266 );
xor ( n26268 , n26197 , n26267 );
xor ( n26269 , n26145 , n26268 );
xor ( n26270 , n26060 , n26269 );
xor ( n26271 , n25935 , n26270 );
and ( n26272 , n24901 , n24905 );
and ( n26273 , n24905 , n25016 );
and ( n26274 , n24901 , n25016 );
or ( n26275 , n26272 , n26273 , n26274 );
and ( n26276 , n25231 , n25247 );
xor ( n26277 , n26275 , n26276 );
and ( n26278 , n25235 , n25236 );
and ( n26279 , n25236 , n25246 );
and ( n26280 , n25235 , n25246 );
or ( n26281 , n26278 , n26279 , n26280 );
and ( n26282 , n24914 , n24939 );
and ( n26283 , n24939 , n24977 );
and ( n26284 , n24914 , n24977 );
or ( n26285 , n26282 , n26283 , n26284 );
and ( n26286 , n25241 , n25245 );
xor ( n26287 , n26285 , n26286 );
and ( n26288 , n24918 , n24922 );
and ( n26289 , n24922 , n24938 );
and ( n26290 , n24918 , n24938 );
or ( n26291 , n26288 , n26289 , n26290 );
and ( n26292 , n25242 , n25244 );
and ( n26293 , n24214 , n606 );
and ( n26294 , n25243 , n615 );
xor ( n26295 , n26293 , n26294 );
buf ( n26296 , n414 );
and ( n26297 , n26296 , n612 );
xor ( n26298 , n26295 , n26297 );
xor ( n26299 , n26292 , n26298 );
xor ( n26300 , n26291 , n26299 );
xor ( n26301 , n26287 , n26300 );
xor ( n26302 , n26281 , n26301 );
xor ( n26303 , n26277 , n26302 );
xor ( n26304 , n26271 , n26303 );
xor ( n26305 , n25931 , n26304 );
and ( n26306 , n24884 , n24888 );
and ( n26307 , n24888 , n25250 );
and ( n26308 , n24884 , n25250 );
or ( n26309 , n26306 , n26307 , n26308 );
xor ( n26310 , n26305 , n26309 );
and ( n26311 , n25251 , n25255 );
and ( n26312 , n25256 , n25259 );
or ( n26313 , n26311 , n26312 );
xor ( n26314 , n26310 , n26313 );
buf ( n26315 , n26314 );
buf ( n26316 , n26315 );
not ( n26317 , n26316 );
nor ( n26318 , n26317 , n8739 );
xor ( n26319 , n25922 , n26318 );
and ( n26320 , n24880 , n25264 );
and ( n26321 , n25265 , n25268 );
or ( n26322 , n26320 , n26321 );
xor ( n26323 , n26319 , n26322 );
buf ( n26324 , n26323 );
buf ( n26325 , n26324 );
not ( n26326 , n26325 );
buf ( n26327 , n555 );
not ( n26328 , n26327 );
nor ( n26329 , n26326 , n26328 );
xor ( n26330 , n25598 , n26329 );
xor ( n26331 , n25280 , n25595 );
nor ( n26332 , n25272 , n26328 );
and ( n26333 , n26331 , n26332 );
xor ( n26334 , n26331 , n26332 );
xor ( n26335 , n25284 , n25593 );
nor ( n26336 , n24242 , n26328 );
and ( n26337 , n26335 , n26336 );
xor ( n26338 , n26335 , n26336 );
xor ( n26339 , n25288 , n25591 );
nor ( n26340 , n23225 , n26328 );
and ( n26341 , n26339 , n26340 );
xor ( n26342 , n26339 , n26340 );
xor ( n26343 , n25292 , n25589 );
nor ( n26344 , n22231 , n26328 );
and ( n26345 , n26343 , n26344 );
xor ( n26346 , n26343 , n26344 );
xor ( n26347 , n25296 , n25587 );
nor ( n26348 , n21258 , n26328 );
and ( n26349 , n26347 , n26348 );
xor ( n26350 , n26347 , n26348 );
xor ( n26351 , n25300 , n25585 );
nor ( n26352 , n20303 , n26328 );
and ( n26353 , n26351 , n26352 );
xor ( n26354 , n26351 , n26352 );
xor ( n26355 , n25304 , n25583 );
nor ( n26356 , n19365 , n26328 );
and ( n26357 , n26355 , n26356 );
xor ( n26358 , n26355 , n26356 );
xor ( n26359 , n25308 , n25581 );
nor ( n26360 , n18448 , n26328 );
and ( n26361 , n26359 , n26360 );
xor ( n26362 , n26359 , n26360 );
xor ( n26363 , n25312 , n25579 );
nor ( n26364 , n17548 , n26328 );
and ( n26365 , n26363 , n26364 );
xor ( n26366 , n26363 , n26364 );
xor ( n26367 , n25316 , n25577 );
nor ( n26368 , n16669 , n26328 );
and ( n26369 , n26367 , n26368 );
xor ( n26370 , n26367 , n26368 );
xor ( n26371 , n25320 , n25575 );
nor ( n26372 , n15809 , n26328 );
and ( n26373 , n26371 , n26372 );
xor ( n26374 , n26371 , n26372 );
xor ( n26375 , n25324 , n25573 );
nor ( n26376 , n14968 , n26328 );
and ( n26377 , n26375 , n26376 );
xor ( n26378 , n26375 , n26376 );
xor ( n26379 , n25328 , n25571 );
nor ( n26380 , n14147 , n26328 );
and ( n26381 , n26379 , n26380 );
xor ( n26382 , n26379 , n26380 );
xor ( n26383 , n25332 , n25569 );
nor ( n26384 , n13349 , n26328 );
and ( n26385 , n26383 , n26384 );
xor ( n26386 , n26383 , n26384 );
xor ( n26387 , n25336 , n25567 );
nor ( n26388 , n12564 , n26328 );
and ( n26389 , n26387 , n26388 );
xor ( n26390 , n26387 , n26388 );
xor ( n26391 , n25340 , n25565 );
nor ( n26392 , n11799 , n26328 );
and ( n26393 , n26391 , n26392 );
xor ( n26394 , n26391 , n26392 );
xor ( n26395 , n25344 , n25563 );
nor ( n26396 , n11050 , n26328 );
and ( n26397 , n26395 , n26396 );
xor ( n26398 , n26395 , n26396 );
xor ( n26399 , n25348 , n25561 );
nor ( n26400 , n10321 , n26328 );
and ( n26401 , n26399 , n26400 );
xor ( n26402 , n26399 , n26400 );
xor ( n26403 , n25352 , n25559 );
nor ( n26404 , n9429 , n26328 );
and ( n26405 , n26403 , n26404 );
xor ( n26406 , n26403 , n26404 );
xor ( n26407 , n25356 , n25557 );
nor ( n26408 , n8949 , n26328 );
and ( n26409 , n26407 , n26408 );
xor ( n26410 , n26407 , n26408 );
xor ( n26411 , n25360 , n25555 );
nor ( n26412 , n9437 , n26328 );
and ( n26413 , n26411 , n26412 );
xor ( n26414 , n26411 , n26412 );
xor ( n26415 , n25364 , n25553 );
nor ( n26416 , n9446 , n26328 );
and ( n26417 , n26415 , n26416 );
xor ( n26418 , n26415 , n26416 );
xor ( n26419 , n25368 , n25551 );
nor ( n26420 , n9455 , n26328 );
and ( n26421 , n26419 , n26420 );
xor ( n26422 , n26419 , n26420 );
xor ( n26423 , n25372 , n25549 );
nor ( n26424 , n9464 , n26328 );
and ( n26425 , n26423 , n26424 );
xor ( n26426 , n26423 , n26424 );
xor ( n26427 , n25376 , n25547 );
nor ( n26428 , n9473 , n26328 );
and ( n26429 , n26427 , n26428 );
xor ( n26430 , n26427 , n26428 );
xor ( n26431 , n25380 , n25545 );
nor ( n26432 , n9482 , n26328 );
and ( n26433 , n26431 , n26432 );
xor ( n26434 , n26431 , n26432 );
xor ( n26435 , n25384 , n25543 );
nor ( n26436 , n9491 , n26328 );
and ( n26437 , n26435 , n26436 );
xor ( n26438 , n26435 , n26436 );
xor ( n26439 , n25388 , n25541 );
nor ( n26440 , n9500 , n26328 );
and ( n26441 , n26439 , n26440 );
xor ( n26442 , n26439 , n26440 );
xor ( n26443 , n25392 , n25539 );
nor ( n26444 , n9509 , n26328 );
and ( n26445 , n26443 , n26444 );
xor ( n26446 , n26443 , n26444 );
xor ( n26447 , n25396 , n25537 );
nor ( n26448 , n9518 , n26328 );
and ( n26449 , n26447 , n26448 );
xor ( n26450 , n26447 , n26448 );
xor ( n26451 , n25400 , n25535 );
nor ( n26452 , n9527 , n26328 );
and ( n26453 , n26451 , n26452 );
xor ( n26454 , n26451 , n26452 );
xor ( n26455 , n25404 , n25533 );
nor ( n26456 , n9536 , n26328 );
and ( n26457 , n26455 , n26456 );
xor ( n26458 , n26455 , n26456 );
xor ( n26459 , n25408 , n25531 );
nor ( n26460 , n9545 , n26328 );
and ( n26461 , n26459 , n26460 );
xor ( n26462 , n26459 , n26460 );
xor ( n26463 , n25412 , n25529 );
nor ( n26464 , n9554 , n26328 );
and ( n26465 , n26463 , n26464 );
xor ( n26466 , n26463 , n26464 );
xor ( n26467 , n25416 , n25527 );
nor ( n26468 , n9563 , n26328 );
and ( n26469 , n26467 , n26468 );
xor ( n26470 , n26467 , n26468 );
xor ( n26471 , n25420 , n25525 );
nor ( n26472 , n9572 , n26328 );
and ( n26473 , n26471 , n26472 );
xor ( n26474 , n26471 , n26472 );
xor ( n26475 , n25424 , n25523 );
nor ( n26476 , n9581 , n26328 );
and ( n26477 , n26475 , n26476 );
xor ( n26478 , n26475 , n26476 );
xor ( n26479 , n25428 , n25521 );
nor ( n26480 , n9590 , n26328 );
and ( n26481 , n26479 , n26480 );
xor ( n26482 , n26479 , n26480 );
xor ( n26483 , n25432 , n25519 );
nor ( n26484 , n9599 , n26328 );
and ( n26485 , n26483 , n26484 );
xor ( n26486 , n26483 , n26484 );
xor ( n26487 , n25436 , n25517 );
nor ( n26488 , n9608 , n26328 );
and ( n26489 , n26487 , n26488 );
xor ( n26490 , n26487 , n26488 );
xor ( n26491 , n25440 , n25515 );
nor ( n26492 , n9617 , n26328 );
and ( n26493 , n26491 , n26492 );
xor ( n26494 , n26491 , n26492 );
xor ( n26495 , n25444 , n25513 );
nor ( n26496 , n9626 , n26328 );
and ( n26497 , n26495 , n26496 );
xor ( n26498 , n26495 , n26496 );
xor ( n26499 , n25448 , n25511 );
nor ( n26500 , n9635 , n26328 );
and ( n26501 , n26499 , n26500 );
xor ( n26502 , n26499 , n26500 );
xor ( n26503 , n25452 , n25509 );
nor ( n26504 , n9644 , n26328 );
and ( n26505 , n26503 , n26504 );
xor ( n26506 , n26503 , n26504 );
xor ( n26507 , n25456 , n25507 );
nor ( n26508 , n9653 , n26328 );
and ( n26509 , n26507 , n26508 );
xor ( n26510 , n26507 , n26508 );
xor ( n26511 , n25460 , n25505 );
nor ( n26512 , n9662 , n26328 );
and ( n26513 , n26511 , n26512 );
xor ( n26514 , n26511 , n26512 );
xor ( n26515 , n25464 , n25503 );
nor ( n26516 , n9671 , n26328 );
and ( n26517 , n26515 , n26516 );
xor ( n26518 , n26515 , n26516 );
xor ( n26519 , n25468 , n25501 );
nor ( n26520 , n9680 , n26328 );
and ( n26521 , n26519 , n26520 );
xor ( n26522 , n26519 , n26520 );
xor ( n26523 , n25472 , n25499 );
nor ( n26524 , n9689 , n26328 );
and ( n26525 , n26523 , n26524 );
xor ( n26526 , n26523 , n26524 );
xor ( n26527 , n25476 , n25497 );
nor ( n26528 , n9698 , n26328 );
and ( n26529 , n26527 , n26528 );
xor ( n26530 , n26527 , n26528 );
xor ( n26531 , n25480 , n25495 );
nor ( n26532 , n9707 , n26328 );
and ( n26533 , n26531 , n26532 );
xor ( n26534 , n26531 , n26532 );
xor ( n26535 , n25484 , n25493 );
nor ( n26536 , n9716 , n26328 );
and ( n26537 , n26535 , n26536 );
xor ( n26538 , n26535 , n26536 );
xor ( n26539 , n25488 , n25491 );
nor ( n26540 , n9725 , n26328 );
and ( n26541 , n26539 , n26540 );
xor ( n26542 , n26539 , n26540 );
xor ( n26543 , n25489 , n25490 );
nor ( n26544 , n9734 , n26328 );
and ( n26545 , n26543 , n26544 );
xor ( n26546 , n26543 , n26544 );
nor ( n26547 , n9752 , n25274 );
nor ( n26548 , n9743 , n26328 );
and ( n26549 , n26547 , n26548 );
and ( n26550 , n26546 , n26549 );
or ( n26551 , n26545 , n26550 );
and ( n26552 , n26542 , n26551 );
or ( n26553 , n26541 , n26552 );
and ( n26554 , n26538 , n26553 );
or ( n26555 , n26537 , n26554 );
and ( n26556 , n26534 , n26555 );
or ( n26557 , n26533 , n26556 );
and ( n26558 , n26530 , n26557 );
or ( n26559 , n26529 , n26558 );
and ( n26560 , n26526 , n26559 );
or ( n26561 , n26525 , n26560 );
and ( n26562 , n26522 , n26561 );
or ( n26563 , n26521 , n26562 );
and ( n26564 , n26518 , n26563 );
or ( n26565 , n26517 , n26564 );
and ( n26566 , n26514 , n26565 );
or ( n26567 , n26513 , n26566 );
and ( n26568 , n26510 , n26567 );
or ( n26569 , n26509 , n26568 );
and ( n26570 , n26506 , n26569 );
or ( n26571 , n26505 , n26570 );
and ( n26572 , n26502 , n26571 );
or ( n26573 , n26501 , n26572 );
and ( n26574 , n26498 , n26573 );
or ( n26575 , n26497 , n26574 );
and ( n26576 , n26494 , n26575 );
or ( n26577 , n26493 , n26576 );
and ( n26578 , n26490 , n26577 );
or ( n26579 , n26489 , n26578 );
and ( n26580 , n26486 , n26579 );
or ( n26581 , n26485 , n26580 );
and ( n26582 , n26482 , n26581 );
or ( n26583 , n26481 , n26582 );
and ( n26584 , n26478 , n26583 );
or ( n26585 , n26477 , n26584 );
and ( n26586 , n26474 , n26585 );
or ( n26587 , n26473 , n26586 );
and ( n26588 , n26470 , n26587 );
or ( n26589 , n26469 , n26588 );
and ( n26590 , n26466 , n26589 );
or ( n26591 , n26465 , n26590 );
and ( n26592 , n26462 , n26591 );
or ( n26593 , n26461 , n26592 );
and ( n26594 , n26458 , n26593 );
or ( n26595 , n26457 , n26594 );
and ( n26596 , n26454 , n26595 );
or ( n26597 , n26453 , n26596 );
and ( n26598 , n26450 , n26597 );
or ( n26599 , n26449 , n26598 );
and ( n26600 , n26446 , n26599 );
or ( n26601 , n26445 , n26600 );
and ( n26602 , n26442 , n26601 );
or ( n26603 , n26441 , n26602 );
and ( n26604 , n26438 , n26603 );
or ( n26605 , n26437 , n26604 );
and ( n26606 , n26434 , n26605 );
or ( n26607 , n26433 , n26606 );
and ( n26608 , n26430 , n26607 );
or ( n26609 , n26429 , n26608 );
and ( n26610 , n26426 , n26609 );
or ( n26611 , n26425 , n26610 );
and ( n26612 , n26422 , n26611 );
or ( n26613 , n26421 , n26612 );
and ( n26614 , n26418 , n26613 );
or ( n26615 , n26417 , n26614 );
and ( n26616 , n26414 , n26615 );
or ( n26617 , n26413 , n26616 );
and ( n26618 , n26410 , n26617 );
or ( n26619 , n26409 , n26618 );
and ( n26620 , n26406 , n26619 );
or ( n26621 , n26405 , n26620 );
and ( n26622 , n26402 , n26621 );
or ( n26623 , n26401 , n26622 );
and ( n26624 , n26398 , n26623 );
or ( n26625 , n26397 , n26624 );
and ( n26626 , n26394 , n26625 );
or ( n26627 , n26393 , n26626 );
and ( n26628 , n26390 , n26627 );
or ( n26629 , n26389 , n26628 );
and ( n26630 , n26386 , n26629 );
or ( n26631 , n26385 , n26630 );
and ( n26632 , n26382 , n26631 );
or ( n26633 , n26381 , n26632 );
and ( n26634 , n26378 , n26633 );
or ( n26635 , n26377 , n26634 );
and ( n26636 , n26374 , n26635 );
or ( n26637 , n26373 , n26636 );
and ( n26638 , n26370 , n26637 );
or ( n26639 , n26369 , n26638 );
and ( n26640 , n26366 , n26639 );
or ( n26641 , n26365 , n26640 );
and ( n26642 , n26362 , n26641 );
or ( n26643 , n26361 , n26642 );
and ( n26644 , n26358 , n26643 );
or ( n26645 , n26357 , n26644 );
and ( n26646 , n26354 , n26645 );
or ( n26647 , n26353 , n26646 );
and ( n26648 , n26350 , n26647 );
or ( n26649 , n26349 , n26648 );
and ( n26650 , n26346 , n26649 );
or ( n26651 , n26345 , n26650 );
and ( n26652 , n26342 , n26651 );
or ( n26653 , n26341 , n26652 );
and ( n26654 , n26338 , n26653 );
or ( n26655 , n26337 , n26654 );
and ( n26656 , n26334 , n26655 );
or ( n26657 , n26333 , n26656 );
xor ( n26658 , n26330 , n26657 );
buf ( n26659 , n477 );
not ( n26660 , n26659 );
nor ( n26661 , n601 , n26660 );
buf ( n26662 , n26661 );
nor ( n26663 , n622 , n24564 );
xor ( n26664 , n26662 , n26663 );
buf ( n26665 , n26664 );
nor ( n26666 , n646 , n23541 );
xor ( n26667 , n26665 , n26666 );
and ( n26668 , n25602 , n25603 );
buf ( n26669 , n26668 );
xor ( n26670 , n26667 , n26669 );
nor ( n26671 , n684 , n22541 );
xor ( n26672 , n26670 , n26671 );
and ( n26673 , n25605 , n25606 );
and ( n26674 , n25607 , n25609 );
or ( n26675 , n26673 , n26674 );
xor ( n26676 , n26672 , n26675 );
nor ( n26677 , n733 , n21562 );
xor ( n26678 , n26676 , n26677 );
and ( n26679 , n25610 , n25611 );
and ( n26680 , n25612 , n25615 );
or ( n26681 , n26679 , n26680 );
xor ( n26682 , n26678 , n26681 );
nor ( n26683 , n796 , n20601 );
xor ( n26684 , n26682 , n26683 );
and ( n26685 , n25616 , n25617 );
and ( n26686 , n25618 , n25621 );
or ( n26687 , n26685 , n26686 );
xor ( n26688 , n26684 , n26687 );
nor ( n26689 , n868 , n19657 );
xor ( n26690 , n26688 , n26689 );
and ( n26691 , n25622 , n25623 );
and ( n26692 , n25624 , n25627 );
or ( n26693 , n26691 , n26692 );
xor ( n26694 , n26690 , n26693 );
nor ( n26695 , n958 , n18734 );
xor ( n26696 , n26694 , n26695 );
and ( n26697 , n25628 , n25629 );
and ( n26698 , n25630 , n25633 );
or ( n26699 , n26697 , n26698 );
xor ( n26700 , n26696 , n26699 );
nor ( n26701 , n1062 , n17828 );
xor ( n26702 , n26700 , n26701 );
and ( n26703 , n25634 , n25635 );
and ( n26704 , n25636 , n25639 );
or ( n26705 , n26703 , n26704 );
xor ( n26706 , n26702 , n26705 );
nor ( n26707 , n1176 , n16943 );
xor ( n26708 , n26706 , n26707 );
and ( n26709 , n25640 , n25641 );
and ( n26710 , n25642 , n25645 );
or ( n26711 , n26709 , n26710 );
xor ( n26712 , n26708 , n26711 );
nor ( n26713 , n1303 , n16077 );
xor ( n26714 , n26712 , n26713 );
and ( n26715 , n25646 , n25647 );
and ( n26716 , n25648 , n25651 );
or ( n26717 , n26715 , n26716 );
xor ( n26718 , n26714 , n26717 );
nor ( n26719 , n1445 , n15230 );
xor ( n26720 , n26718 , n26719 );
and ( n26721 , n25652 , n25653 );
and ( n26722 , n25654 , n25657 );
or ( n26723 , n26721 , n26722 );
xor ( n26724 , n26720 , n26723 );
nor ( n26725 , n1598 , n14403 );
xor ( n26726 , n26724 , n26725 );
and ( n26727 , n25658 , n25659 );
and ( n26728 , n25660 , n25663 );
or ( n26729 , n26727 , n26728 );
xor ( n26730 , n26726 , n26729 );
nor ( n26731 , n1766 , n13599 );
xor ( n26732 , n26730 , n26731 );
and ( n26733 , n25664 , n25665 );
and ( n26734 , n25666 , n25669 );
or ( n26735 , n26733 , n26734 );
xor ( n26736 , n26732 , n26735 );
nor ( n26737 , n1945 , n12808 );
xor ( n26738 , n26736 , n26737 );
and ( n26739 , n25670 , n25671 );
and ( n26740 , n25672 , n25675 );
or ( n26741 , n26739 , n26740 );
xor ( n26742 , n26738 , n26741 );
nor ( n26743 , n2137 , n12037 );
xor ( n26744 , n26742 , n26743 );
and ( n26745 , n25676 , n25677 );
and ( n26746 , n25678 , n25681 );
or ( n26747 , n26745 , n26746 );
xor ( n26748 , n26744 , n26747 );
nor ( n26749 , n2343 , n11282 );
xor ( n26750 , n26748 , n26749 );
and ( n26751 , n25682 , n25683 );
and ( n26752 , n25684 , n25687 );
or ( n26753 , n26751 , n26752 );
xor ( n26754 , n26750 , n26753 );
nor ( n26755 , n2566 , n10547 );
xor ( n26756 , n26754 , n26755 );
and ( n26757 , n25688 , n25689 );
and ( n26758 , n25690 , n25693 );
or ( n26759 , n26757 , n26758 );
xor ( n26760 , n26756 , n26759 );
nor ( n26761 , n2797 , n9829 );
xor ( n26762 , n26760 , n26761 );
and ( n26763 , n25694 , n25695 );
and ( n26764 , n25696 , n25699 );
or ( n26765 , n26763 , n26764 );
xor ( n26766 , n26762 , n26765 );
nor ( n26767 , n3043 , n8955 );
xor ( n26768 , n26766 , n26767 );
and ( n26769 , n25700 , n25701 );
and ( n26770 , n25702 , n25705 );
or ( n26771 , n26769 , n26770 );
xor ( n26772 , n26768 , n26771 );
nor ( n26773 , n3300 , n603 );
xor ( n26774 , n26772 , n26773 );
and ( n26775 , n25706 , n25707 );
and ( n26776 , n25708 , n25711 );
or ( n26777 , n26775 , n26776 );
xor ( n26778 , n26774 , n26777 );
nor ( n26779 , n3570 , n652 );
xor ( n26780 , n26778 , n26779 );
and ( n26781 , n25712 , n25713 );
and ( n26782 , n25714 , n25717 );
or ( n26783 , n26781 , n26782 );
xor ( n26784 , n26780 , n26783 );
nor ( n26785 , n3853 , n624 );
xor ( n26786 , n26784 , n26785 );
and ( n26787 , n25718 , n25719 );
and ( n26788 , n25720 , n25723 );
or ( n26789 , n26787 , n26788 );
xor ( n26790 , n26786 , n26789 );
nor ( n26791 , n4151 , n648 );
xor ( n26792 , n26790 , n26791 );
and ( n26793 , n25724 , n25725 );
and ( n26794 , n25726 , n25729 );
or ( n26795 , n26793 , n26794 );
xor ( n26796 , n26792 , n26795 );
nor ( n26797 , n4458 , n686 );
xor ( n26798 , n26796 , n26797 );
and ( n26799 , n25730 , n25731 );
and ( n26800 , n25732 , n25735 );
or ( n26801 , n26799 , n26800 );
xor ( n26802 , n26798 , n26801 );
nor ( n26803 , n4786 , n735 );
xor ( n26804 , n26802 , n26803 );
and ( n26805 , n25736 , n25737 );
and ( n26806 , n25738 , n25741 );
or ( n26807 , n26805 , n26806 );
xor ( n26808 , n26804 , n26807 );
nor ( n26809 , n5126 , n798 );
xor ( n26810 , n26808 , n26809 );
and ( n26811 , n25742 , n25743 );
and ( n26812 , n25744 , n25747 );
or ( n26813 , n26811 , n26812 );
xor ( n26814 , n26810 , n26813 );
nor ( n26815 , n5477 , n870 );
xor ( n26816 , n26814 , n26815 );
and ( n26817 , n25748 , n25749 );
and ( n26818 , n25750 , n25753 );
or ( n26819 , n26817 , n26818 );
xor ( n26820 , n26816 , n26819 );
nor ( n26821 , n5838 , n960 );
xor ( n26822 , n26820 , n26821 );
and ( n26823 , n25754 , n25755 );
and ( n26824 , n25756 , n25759 );
or ( n26825 , n26823 , n26824 );
xor ( n26826 , n26822 , n26825 );
nor ( n26827 , n6212 , n1064 );
xor ( n26828 , n26826 , n26827 );
and ( n26829 , n25760 , n25761 );
and ( n26830 , n25762 , n25765 );
or ( n26831 , n26829 , n26830 );
xor ( n26832 , n26828 , n26831 );
nor ( n26833 , n6596 , n1178 );
xor ( n26834 , n26832 , n26833 );
and ( n26835 , n25766 , n25767 );
and ( n26836 , n25768 , n25771 );
or ( n26837 , n26835 , n26836 );
xor ( n26838 , n26834 , n26837 );
nor ( n26839 , n6997 , n1305 );
xor ( n26840 , n26838 , n26839 );
and ( n26841 , n25772 , n25773 );
and ( n26842 , n25774 , n25777 );
or ( n26843 , n26841 , n26842 );
xor ( n26844 , n26840 , n26843 );
nor ( n26845 , n7413 , n1447 );
xor ( n26846 , n26844 , n26845 );
and ( n26847 , n25778 , n25779 );
and ( n26848 , n25780 , n25783 );
or ( n26849 , n26847 , n26848 );
xor ( n26850 , n26846 , n26849 );
nor ( n26851 , n7841 , n1600 );
xor ( n26852 , n26850 , n26851 );
and ( n26853 , n25784 , n25785 );
and ( n26854 , n25786 , n25789 );
or ( n26855 , n26853 , n26854 );
xor ( n26856 , n26852 , n26855 );
nor ( n26857 , n8281 , n1768 );
xor ( n26858 , n26856 , n26857 );
and ( n26859 , n25790 , n25791 );
and ( n26860 , n25792 , n25795 );
or ( n26861 , n26859 , n26860 );
xor ( n26862 , n26858 , n26861 );
nor ( n26863 , n8737 , n1947 );
xor ( n26864 , n26862 , n26863 );
and ( n26865 , n25796 , n25797 );
and ( n26866 , n25798 , n25801 );
or ( n26867 , n26865 , n26866 );
xor ( n26868 , n26864 , n26867 );
nor ( n26869 , n9420 , n2139 );
xor ( n26870 , n26868 , n26869 );
and ( n26871 , n25802 , n25803 );
and ( n26872 , n25804 , n25807 );
or ( n26873 , n26871 , n26872 );
xor ( n26874 , n26870 , n26873 );
nor ( n26875 , n10312 , n2345 );
xor ( n26876 , n26874 , n26875 );
and ( n26877 , n25808 , n25809 );
and ( n26878 , n25810 , n25813 );
or ( n26879 , n26877 , n26878 );
xor ( n26880 , n26876 , n26879 );
nor ( n26881 , n11041 , n2568 );
xor ( n26882 , n26880 , n26881 );
and ( n26883 , n25814 , n25815 );
and ( n26884 , n25816 , n25819 );
or ( n26885 , n26883 , n26884 );
xor ( n26886 , n26882 , n26885 );
nor ( n26887 , n11790 , n2799 );
xor ( n26888 , n26886 , n26887 );
and ( n26889 , n25820 , n25821 );
and ( n26890 , n25822 , n25825 );
or ( n26891 , n26889 , n26890 );
xor ( n26892 , n26888 , n26891 );
nor ( n26893 , n12555 , n3045 );
xor ( n26894 , n26892 , n26893 );
and ( n26895 , n25826 , n25827 );
and ( n26896 , n25828 , n25831 );
or ( n26897 , n26895 , n26896 );
xor ( n26898 , n26894 , n26897 );
nor ( n26899 , n13340 , n3302 );
xor ( n26900 , n26898 , n26899 );
and ( n26901 , n25832 , n25833 );
and ( n26902 , n25834 , n25837 );
or ( n26903 , n26901 , n26902 );
xor ( n26904 , n26900 , n26903 );
nor ( n26905 , n14138 , n3572 );
xor ( n26906 , n26904 , n26905 );
and ( n26907 , n25838 , n25839 );
and ( n26908 , n25840 , n25843 );
or ( n26909 , n26907 , n26908 );
xor ( n26910 , n26906 , n26909 );
nor ( n26911 , n14959 , n3855 );
xor ( n26912 , n26910 , n26911 );
and ( n26913 , n25844 , n25845 );
and ( n26914 , n25846 , n25849 );
or ( n26915 , n26913 , n26914 );
xor ( n26916 , n26912 , n26915 );
nor ( n26917 , n15800 , n4153 );
xor ( n26918 , n26916 , n26917 );
and ( n26919 , n25850 , n25851 );
and ( n26920 , n25852 , n25855 );
or ( n26921 , n26919 , n26920 );
xor ( n26922 , n26918 , n26921 );
nor ( n26923 , n16660 , n4460 );
xor ( n26924 , n26922 , n26923 );
and ( n26925 , n25856 , n25857 );
and ( n26926 , n25858 , n25861 );
or ( n26927 , n26925 , n26926 );
xor ( n26928 , n26924 , n26927 );
nor ( n26929 , n17539 , n4788 );
xor ( n26930 , n26928 , n26929 );
and ( n26931 , n25862 , n25863 );
and ( n26932 , n25864 , n25867 );
or ( n26933 , n26931 , n26932 );
xor ( n26934 , n26930 , n26933 );
nor ( n26935 , n18439 , n5128 );
xor ( n26936 , n26934 , n26935 );
and ( n26937 , n25868 , n25869 );
and ( n26938 , n25870 , n25873 );
or ( n26939 , n26937 , n26938 );
xor ( n26940 , n26936 , n26939 );
nor ( n26941 , n19356 , n5479 );
xor ( n26942 , n26940 , n26941 );
and ( n26943 , n25874 , n25875 );
and ( n26944 , n25876 , n25879 );
or ( n26945 , n26943 , n26944 );
xor ( n26946 , n26942 , n26945 );
nor ( n26947 , n20294 , n5840 );
xor ( n26948 , n26946 , n26947 );
and ( n26949 , n25880 , n25881 );
and ( n26950 , n25882 , n25885 );
or ( n26951 , n26949 , n26950 );
xor ( n26952 , n26948 , n26951 );
nor ( n26953 , n21249 , n6214 );
xor ( n26954 , n26952 , n26953 );
and ( n26955 , n25886 , n25887 );
and ( n26956 , n25888 , n25891 );
or ( n26957 , n26955 , n26956 );
xor ( n26958 , n26954 , n26957 );
nor ( n26959 , n22222 , n6598 );
xor ( n26960 , n26958 , n26959 );
and ( n26961 , n25892 , n25893 );
and ( n26962 , n25894 , n25897 );
or ( n26963 , n26961 , n26962 );
xor ( n26964 , n26960 , n26963 );
nor ( n26965 , n23216 , n6999 );
xor ( n26966 , n26964 , n26965 );
and ( n26967 , n25898 , n25899 );
and ( n26968 , n25900 , n25903 );
or ( n26969 , n26967 , n26968 );
xor ( n26970 , n26966 , n26969 );
nor ( n26971 , n24233 , n7415 );
xor ( n26972 , n26970 , n26971 );
and ( n26973 , n25904 , n25905 );
and ( n26974 , n25906 , n25909 );
or ( n26975 , n26973 , n26974 );
xor ( n26976 , n26972 , n26975 );
nor ( n26977 , n25263 , n7843 );
xor ( n26978 , n26976 , n26977 );
and ( n26979 , n25910 , n25911 );
and ( n26980 , n25912 , n25915 );
or ( n26981 , n26979 , n26980 );
xor ( n26982 , n26978 , n26981 );
nor ( n26983 , n26317 , n8283 );
xor ( n26984 , n26982 , n26983 );
and ( n26985 , n25916 , n25917 );
and ( n26986 , n25918 , n25921 );
or ( n26987 , n26985 , n26986 );
xor ( n26988 , n26984 , n26987 );
and ( n26989 , n26275 , n26276 );
and ( n26990 , n26276 , n26302 );
and ( n26991 , n26275 , n26302 );
or ( n26992 , n26989 , n26990 , n26991 );
and ( n26993 , n25935 , n26270 );
and ( n26994 , n26270 , n26303 );
and ( n26995 , n25935 , n26303 );
or ( n26996 , n26993 , n26994 , n26995 );
xor ( n26997 , n26992 , n26996 );
and ( n26998 , n25939 , n26059 );
and ( n26999 , n26059 , n26269 );
and ( n27000 , n25939 , n26269 );
or ( n27001 , n26998 , n26999 , n27000 );
and ( n27002 , n26064 , n26144 );
and ( n27003 , n26144 , n26268 );
and ( n27004 , n26064 , n26268 );
or ( n27005 , n27002 , n27003 , n27004 );
and ( n27006 , n25952 , n26020 );
and ( n27007 , n26020 , n26057 );
and ( n27008 , n25952 , n26057 );
or ( n27009 , n27006 , n27007 , n27008 );
and ( n27010 , n26068 , n26072 );
and ( n27011 , n26072 , n26143 );
and ( n27012 , n26068 , n26143 );
or ( n27013 , n27010 , n27011 , n27012 );
xor ( n27014 , n27009 , n27013 );
and ( n27015 , n26025 , n26029 );
and ( n27016 , n26029 , n26056 );
and ( n27017 , n26025 , n26056 );
or ( n27018 , n27015 , n27016 , n27017 );
and ( n27019 , n25986 , n26002 );
and ( n27020 , n26002 , n26018 );
and ( n27021 , n25986 , n26018 );
or ( n27022 , n27019 , n27020 , n27021 );
and ( n27023 , n25969 , n25973 );
and ( n27024 , n25973 , n25979 );
and ( n27025 , n25969 , n25979 );
or ( n27026 , n27023 , n27024 , n27025 );
and ( n27027 , n25990 , n25995 );
and ( n27028 , n25995 , n26001 );
and ( n27029 , n25990 , n26001 );
or ( n27030 , n27027 , n27028 , n27029 );
xor ( n27031 , n27026 , n27030 );
and ( n27032 , n25975 , n25976 );
and ( n27033 , n25976 , n25978 );
and ( n27034 , n25975 , n25978 );
or ( n27035 , n27032 , n27033 , n27034 );
and ( n27036 , n25991 , n25992 );
and ( n27037 , n25992 , n25994 );
and ( n27038 , n25991 , n25994 );
or ( n27039 , n27036 , n27037 , n27038 );
xor ( n27040 , n27035 , n27039 );
and ( n27041 , n21216 , n771 );
and ( n27042 , n22186 , n719 );
xor ( n27043 , n27041 , n27042 );
and ( n27044 , n22892 , n663 );
xor ( n27045 , n27043 , n27044 );
xor ( n27046 , n27040 , n27045 );
xor ( n27047 , n27031 , n27046 );
xor ( n27048 , n27022 , n27047 );
and ( n27049 , n26007 , n26011 );
and ( n27050 , n26011 , n26017 );
and ( n27051 , n26007 , n26017 );
or ( n27052 , n27049 , n27050 , n27051 );
and ( n27053 , n25997 , n25998 );
and ( n27054 , n25998 , n26000 );
and ( n27055 , n25997 , n26000 );
or ( n27056 , n27053 , n27054 , n27055 );
and ( n27057 , n18144 , n1034 );
and ( n27058 , n19324 , n940 );
xor ( n27059 , n27057 , n27058 );
and ( n27060 , n20233 , n840 );
xor ( n27061 , n27059 , n27060 );
xor ( n27062 , n27056 , n27061 );
and ( n27063 , n15758 , n1424 );
and ( n27064 , n16637 , n1254 );
xor ( n27065 , n27063 , n27064 );
and ( n27066 , n17512 , n1134 );
xor ( n27067 , n27065 , n27066 );
xor ( n27068 , n27062 , n27067 );
xor ( n27069 , n27052 , n27068 );
and ( n27070 , n26013 , n26014 );
and ( n27071 , n26014 , n26016 );
and ( n27072 , n26013 , n26016 );
or ( n27073 , n27070 , n27071 , n27072 );
and ( n27074 , n26044 , n26045 );
and ( n27075 , n26045 , n26047 );
and ( n27076 , n26044 , n26047 );
or ( n27077 , n27074 , n27075 , n27076 );
xor ( n27078 , n27073 , n27077 );
and ( n27079 , n13322 , n1882 );
and ( n27080 , n14118 , n1738 );
xor ( n27081 , n27079 , n27080 );
and ( n27082 , n14938 , n1551 );
xor ( n27083 , n27081 , n27082 );
xor ( n27084 , n27078 , n27083 );
xor ( n27085 , n27069 , n27084 );
xor ( n27086 , n27048 , n27085 );
xor ( n27087 , n27018 , n27086 );
and ( n27088 , n26034 , n26038 );
and ( n27089 , n26038 , n26055 );
and ( n27090 , n26034 , n26055 );
or ( n27091 , n27088 , n27089 , n27090 );
and ( n27092 , n26107 , n26122 );
and ( n27093 , n26122 , n26141 );
and ( n27094 , n26107 , n26141 );
or ( n27095 , n27092 , n27093 , n27094 );
xor ( n27096 , n27091 , n27095 );
and ( n27097 , n26043 , n26048 );
and ( n27098 , n26048 , n26054 );
and ( n27099 , n26043 , n26054 );
or ( n27100 , n27097 , n27098 , n27099 );
and ( n27101 , n26111 , n26115 );
and ( n27102 , n26115 , n26121 );
and ( n27103 , n26111 , n26121 );
or ( n27104 , n27101 , n27102 , n27103 );
xor ( n27105 , n27100 , n27104 );
and ( n27106 , n26050 , n26051 );
and ( n27107 , n26051 , n26053 );
and ( n27108 , n26050 , n26053 );
or ( n27109 , n27106 , n27107 , n27108 );
and ( n27110 , n11015 , n2544 );
and ( n27111 , n11769 , n2298 );
xor ( n27112 , n27110 , n27111 );
and ( n27113 , n12320 , n2100 );
xor ( n27114 , n27112 , n27113 );
xor ( n27115 , n27109 , n27114 );
and ( n27116 , n8718 , n3271 );
and ( n27117 , n9400 , n2981 );
xor ( n27118 , n27116 , n27117 );
and ( n27119 , n10291 , n2739 );
xor ( n27120 , n27118 , n27119 );
xor ( n27121 , n27115 , n27120 );
xor ( n27122 , n27105 , n27121 );
xor ( n27123 , n27096 , n27122 );
xor ( n27124 , n27087 , n27123 );
xor ( n27125 , n27014 , n27124 );
xor ( n27126 , n27005 , n27125 );
and ( n27127 , n26149 , n26196 );
and ( n27128 , n26196 , n26267 );
and ( n27129 , n26149 , n26267 );
or ( n27130 , n27127 , n27128 , n27129 );
and ( n27131 , n26077 , n26102 );
and ( n27132 , n26102 , n26142 );
and ( n27133 , n26077 , n26142 );
or ( n27134 , n27131 , n27132 , n27133 );
and ( n27135 , n26153 , n26157 );
and ( n27136 , n26157 , n26195 );
and ( n27137 , n26153 , n26195 );
or ( n27138 , n27135 , n27136 , n27137 );
xor ( n27139 , n27134 , n27138 );
and ( n27140 , n26081 , n26085 );
and ( n27141 , n26085 , n26101 );
and ( n27142 , n26081 , n26101 );
or ( n27143 , n27140 , n27141 , n27142 );
and ( n27144 , n26166 , n26171 );
and ( n27145 , n26171 , n26177 );
and ( n27146 , n26166 , n26177 );
or ( n27147 , n27144 , n27145 , n27146 );
and ( n27148 , n26090 , n26094 );
and ( n27149 , n26094 , n26100 );
and ( n27150 , n26090 , n26100 );
or ( n27151 , n27148 , n27149 , n27150 );
xor ( n27152 , n27147 , n27151 );
and ( n27153 , n26096 , n26097 );
and ( n27154 , n26097 , n26099 );
and ( n27155 , n26096 , n26099 );
or ( n27156 , n27153 , n27154 , n27155 );
and ( n27157 , n26167 , n26168 );
and ( n27158 , n26168 , n26170 );
and ( n27159 , n26167 , n26170 );
or ( n27160 , n27157 , n27158 , n27159 );
xor ( n27161 , n27156 , n27160 );
and ( n27162 , n4132 , n7310 );
and ( n27163 , n4438 , n6971 );
xor ( n27164 , n27162 , n27163 );
and ( n27165 , n4766 , n6504 );
xor ( n27166 , n27164 , n27165 );
xor ( n27167 , n27161 , n27166 );
xor ( n27168 , n27152 , n27167 );
xor ( n27169 , n27143 , n27168 );
and ( n27170 , n26129 , n26134 );
and ( n27171 , n26134 , n26140 );
and ( n27172 , n26129 , n26140 );
or ( n27173 , n27170 , n27171 , n27172 );
and ( n27174 , n26117 , n26118 );
and ( n27175 , n26118 , n26120 );
and ( n27176 , n26117 , n26120 );
or ( n27177 , n27174 , n27175 , n27176 );
and ( n27178 , n26130 , n26131 );
and ( n27179 , n26131 , n26133 );
and ( n27180 , n26130 , n26133 );
or ( n27181 , n27178 , n27179 , n27180 );
xor ( n27182 , n27177 , n27181 );
and ( n27183 , n7385 , n4102 );
and ( n27184 , n7808 , n3749 );
xor ( n27185 , n27183 , n27184 );
and ( n27186 , n8079 , n3495 );
xor ( n27187 , n27185 , n27186 );
xor ( n27188 , n27182 , n27187 );
xor ( n27189 , n27173 , n27188 );
and ( n27190 , n26136 , n26137 );
and ( n27191 , n26137 , n26139 );
and ( n27192 , n26136 , n26139 );
or ( n27193 , n27190 , n27191 , n27192 );
and ( n27194 , n6187 , n5103 );
and ( n27195 , n6569 , n4730 );
xor ( n27196 , n27194 , n27195 );
and ( n27197 , n6816 , n4403 );
xor ( n27198 , n27196 , n27197 );
xor ( n27199 , n27193 , n27198 );
and ( n27200 , n4959 , n6132 );
and ( n27201 , n5459 , n5765 );
xor ( n27202 , n27200 , n27201 );
and ( n27203 , n5819 , n5408 );
xor ( n27204 , n27202 , n27203 );
xor ( n27205 , n27199 , n27204 );
xor ( n27206 , n27189 , n27205 );
xor ( n27207 , n27169 , n27206 );
xor ( n27208 , n27139 , n27207 );
xor ( n27209 , n27130 , n27208 );
and ( n27210 , n26201 , n26239 );
and ( n27211 , n26239 , n26266 );
and ( n27212 , n26201 , n26266 );
or ( n27213 , n27210 , n27211 , n27212 );
and ( n27214 , n26244 , n26248 );
and ( n27215 , n26248 , n26265 );
and ( n27216 , n26244 , n26265 );
or ( n27217 , n27214 , n27215 , n27216 );
and ( n27218 , n26162 , n26178 );
and ( n27219 , n26178 , n26194 );
and ( n27220 , n26162 , n26194 );
or ( n27221 , n27218 , n27219 , n27220 );
xor ( n27222 , n27217 , n27221 );
and ( n27223 , n26183 , n26187 );
and ( n27224 , n26187 , n26193 );
and ( n27225 , n26183 , n26193 );
or ( n27226 , n27223 , n27224 , n27225 );
and ( n27227 , n26173 , n26174 );
and ( n27228 , n26174 , n26176 );
and ( n27229 , n26173 , n26176 );
or ( n27230 , n27227 , n27228 , n27229 );
and ( n27231 , n3182 , n8669 );
and ( n27232 , n3545 , n8243 );
xor ( n27233 , n27231 , n27232 );
and ( n27234 , n3801 , n7662 );
xor ( n27235 , n27233 , n27234 );
xor ( n27236 , n27230 , n27235 );
and ( n27237 , n2462 , n10977 );
and ( n27238 , n2779 , n10239 );
xor ( n27239 , n27237 , n27238 );
and ( n27240 , n3024 , n9348 );
xor ( n27241 , n27239 , n27240 );
xor ( n27242 , n27236 , n27241 );
xor ( n27243 , n27226 , n27242 );
and ( n27244 , n26189 , n26190 );
and ( n27245 , n26190 , n26192 );
and ( n27246 , n26189 , n26192 );
or ( n27247 , n27244 , n27245 , n27246 );
and ( n27248 , n26254 , n26255 );
and ( n27249 , n26255 , n26257 );
and ( n27250 , n26254 , n26257 );
or ( n27251 , n27248 , n27249 , n27250 );
xor ( n27252 , n27247 , n27251 );
and ( n27253 , n1933 , n13256 );
and ( n27254 , n2120 , n12531 );
xor ( n27255 , n27253 , n27254 );
and ( n27256 , n2324 , n11718 );
xor ( n27257 , n27255 , n27256 );
xor ( n27258 , n27252 , n27257 );
xor ( n27259 , n27243 , n27258 );
xor ( n27260 , n27222 , n27259 );
xor ( n27261 , n27213 , n27260 );
and ( n27262 , n26205 , n26222 );
and ( n27263 , n26222 , n26238 );
and ( n27264 , n26205 , n26238 );
or ( n27265 , n27262 , n27263 , n27264 );
and ( n27266 , n26209 , n26214 );
and ( n27267 , n26214 , n26221 );
and ( n27268 , n26209 , n26221 );
or ( n27269 , n27266 , n27267 , n27268 );
and ( n27270 , n26233 , n26234 );
and ( n27271 , n26234 , n26236 );
and ( n27272 , n26233 , n26236 );
or ( n27273 , n27270 , n27271 , n27272 );
and ( n27274 , n26210 , n26211 );
and ( n27275 , n26211 , n26213 );
and ( n27276 , n26210 , n26213 );
or ( n27277 , n27274 , n27275 , n27276 );
xor ( n27278 , n27273 , n27277 );
and ( n27279 , n783 , n20976 );
and ( n27280 , n856 , n20156 );
xor ( n27281 , n27279 , n27280 );
and ( n27282 , n925 , n19222 );
xor ( n27283 , n27281 , n27282 );
xor ( n27284 , n27278 , n27283 );
xor ( n27285 , n27269 , n27284 );
and ( n27286 , n26217 , n26218 );
and ( n27287 , n26218 , n26220 );
and ( n27288 , n26217 , n26220 );
or ( n27289 , n27286 , n27287 , n27288 );
and ( n27290 , n632 , n24137 );
and ( n27291 , n671 , n23075 );
xor ( n27292 , n27290 , n27291 );
and ( n27293 , n715 , n22065 );
xor ( n27294 , n27292 , n27293 );
xor ( n27295 , n27289 , n27294 );
buf ( n27296 , n413 );
and ( n27297 , n599 , n27296 );
and ( n27298 , n608 , n26216 );
xor ( n27299 , n27297 , n27298 );
and ( n27300 , n611 , n25163 );
xor ( n27301 , n27299 , n27300 );
xor ( n27302 , n27295 , n27301 );
xor ( n27303 , n27285 , n27302 );
xor ( n27304 , n27265 , n27303 );
and ( n27305 , n26227 , n26231 );
and ( n27306 , n26231 , n26237 );
and ( n27307 , n26227 , n26237 );
or ( n27308 , n27305 , n27306 , n27307 );
and ( n27309 , n26253 , n26258 );
and ( n27310 , n26258 , n26264 );
and ( n27311 , n26253 , n26264 );
or ( n27312 , n27309 , n27310 , n27311 );
xor ( n27313 , n27308 , n27312 );
and ( n27314 , n26260 , n26261 );
and ( n27315 , n26261 , n26263 );
and ( n27316 , n26260 , n26263 );
or ( n27317 , n27314 , n27315 , n27316 );
and ( n27318 , n1383 , n15691 );
and ( n27319 , n1580 , n14838 );
xor ( n27320 , n27318 , n27319 );
and ( n27321 , n1694 , n14044 );
xor ( n27322 , n27320 , n27321 );
xor ( n27323 , n27317 , n27322 );
and ( n27324 , n1047 , n18407 );
and ( n27325 , n1164 , n17422 );
xor ( n27326 , n27324 , n27325 );
and ( n27327 , n1287 , n16550 );
xor ( n27328 , n27326 , n27327 );
xor ( n27329 , n27323 , n27328 );
xor ( n27330 , n27313 , n27329 );
xor ( n27331 , n27304 , n27330 );
xor ( n27332 , n27261 , n27331 );
xor ( n27333 , n27209 , n27332 );
xor ( n27334 , n27126 , n27333 );
xor ( n27335 , n27001 , n27334 );
and ( n27336 , n25943 , n25947 );
and ( n27337 , n25947 , n26058 );
and ( n27338 , n25943 , n26058 );
or ( n27339 , n27336 , n27337 , n27338 );
and ( n27340 , n26281 , n26301 );
xor ( n27341 , n27339 , n27340 );
and ( n27342 , n26285 , n26286 );
and ( n27343 , n26286 , n26300 );
and ( n27344 , n26285 , n26300 );
or ( n27345 , n27342 , n27343 , n27344 );
and ( n27346 , n25956 , n25981 );
and ( n27347 , n25981 , n26019 );
and ( n27348 , n25956 , n26019 );
or ( n27349 , n27346 , n27347 , n27348 );
and ( n27350 , n26291 , n26299 );
xor ( n27351 , n27349 , n27350 );
and ( n27352 , n25960 , n25964 );
and ( n27353 , n25964 , n25980 );
and ( n27354 , n25960 , n25980 );
or ( n27355 , n27352 , n27353 , n27354 );
and ( n27356 , n26292 , n26298 );
and ( n27357 , n26293 , n26294 );
and ( n27358 , n26294 , n26297 );
and ( n27359 , n26293 , n26297 );
or ( n27360 , n27357 , n27358 , n27359 );
buf ( n27361 , n413 );
and ( n27362 , n27361 , n612 );
xor ( n27363 , n27360 , n27362 );
and ( n27364 , n24214 , n635 );
and ( n27365 , n25243 , n606 );
xor ( n27366 , n27364 , n27365 );
and ( n27367 , n26296 , n615 );
xor ( n27368 , n27366 , n27367 );
xor ( n27369 , n27363 , n27368 );
xor ( n27370 , n27356 , n27369 );
xor ( n27371 , n27355 , n27370 );
xor ( n27372 , n27351 , n27371 );
xor ( n27373 , n27345 , n27372 );
xor ( n27374 , n27341 , n27373 );
xor ( n27375 , n27335 , n27374 );
xor ( n27376 , n26997 , n27375 );
and ( n27377 , n25926 , n25930 );
and ( n27378 , n25930 , n26304 );
and ( n27379 , n25926 , n26304 );
or ( n27380 , n27377 , n27378 , n27379 );
xor ( n27381 , n27376 , n27380 );
and ( n27382 , n26305 , n26309 );
and ( n27383 , n26310 , n26313 );
or ( n27384 , n27382 , n27383 );
xor ( n27385 , n27381 , n27384 );
buf ( n27386 , n27385 );
buf ( n27387 , n27386 );
not ( n27388 , n27387 );
nor ( n27389 , n27388 , n8739 );
xor ( n27390 , n26988 , n27389 );
and ( n27391 , n25922 , n26318 );
and ( n27392 , n26319 , n26322 );
or ( n27393 , n27391 , n27392 );
xor ( n27394 , n27390 , n27393 );
buf ( n27395 , n27394 );
buf ( n27396 , n27395 );
not ( n27397 , n27396 );
buf ( n27398 , n556 );
not ( n27399 , n27398 );
nor ( n27400 , n27397 , n27399 );
xor ( n27401 , n26658 , n27400 );
xor ( n27402 , n26334 , n26655 );
nor ( n27403 , n26326 , n27399 );
and ( n27404 , n27402 , n27403 );
xor ( n27405 , n27402 , n27403 );
xor ( n27406 , n26338 , n26653 );
nor ( n27407 , n25272 , n27399 );
and ( n27408 , n27406 , n27407 );
xor ( n27409 , n27406 , n27407 );
xor ( n27410 , n26342 , n26651 );
nor ( n27411 , n24242 , n27399 );
and ( n27412 , n27410 , n27411 );
xor ( n27413 , n27410 , n27411 );
xor ( n27414 , n26346 , n26649 );
nor ( n27415 , n23225 , n27399 );
and ( n27416 , n27414 , n27415 );
xor ( n27417 , n27414 , n27415 );
xor ( n27418 , n26350 , n26647 );
nor ( n27419 , n22231 , n27399 );
and ( n27420 , n27418 , n27419 );
xor ( n27421 , n27418 , n27419 );
xor ( n27422 , n26354 , n26645 );
nor ( n27423 , n21258 , n27399 );
and ( n27424 , n27422 , n27423 );
xor ( n27425 , n27422 , n27423 );
xor ( n27426 , n26358 , n26643 );
nor ( n27427 , n20303 , n27399 );
and ( n27428 , n27426 , n27427 );
xor ( n27429 , n27426 , n27427 );
xor ( n27430 , n26362 , n26641 );
nor ( n27431 , n19365 , n27399 );
and ( n27432 , n27430 , n27431 );
xor ( n27433 , n27430 , n27431 );
xor ( n27434 , n26366 , n26639 );
nor ( n27435 , n18448 , n27399 );
and ( n27436 , n27434 , n27435 );
xor ( n27437 , n27434 , n27435 );
xor ( n27438 , n26370 , n26637 );
nor ( n27439 , n17548 , n27399 );
and ( n27440 , n27438 , n27439 );
xor ( n27441 , n27438 , n27439 );
xor ( n27442 , n26374 , n26635 );
nor ( n27443 , n16669 , n27399 );
and ( n27444 , n27442 , n27443 );
xor ( n27445 , n27442 , n27443 );
xor ( n27446 , n26378 , n26633 );
nor ( n27447 , n15809 , n27399 );
and ( n27448 , n27446 , n27447 );
xor ( n27449 , n27446 , n27447 );
xor ( n27450 , n26382 , n26631 );
nor ( n27451 , n14968 , n27399 );
and ( n27452 , n27450 , n27451 );
xor ( n27453 , n27450 , n27451 );
xor ( n27454 , n26386 , n26629 );
nor ( n27455 , n14147 , n27399 );
and ( n27456 , n27454 , n27455 );
xor ( n27457 , n27454 , n27455 );
xor ( n27458 , n26390 , n26627 );
nor ( n27459 , n13349 , n27399 );
and ( n27460 , n27458 , n27459 );
xor ( n27461 , n27458 , n27459 );
xor ( n27462 , n26394 , n26625 );
nor ( n27463 , n12564 , n27399 );
and ( n27464 , n27462 , n27463 );
xor ( n27465 , n27462 , n27463 );
xor ( n27466 , n26398 , n26623 );
nor ( n27467 , n11799 , n27399 );
and ( n27468 , n27466 , n27467 );
xor ( n27469 , n27466 , n27467 );
xor ( n27470 , n26402 , n26621 );
nor ( n27471 , n11050 , n27399 );
and ( n27472 , n27470 , n27471 );
xor ( n27473 , n27470 , n27471 );
xor ( n27474 , n26406 , n26619 );
nor ( n27475 , n10321 , n27399 );
and ( n27476 , n27474 , n27475 );
xor ( n27477 , n27474 , n27475 );
xor ( n27478 , n26410 , n26617 );
nor ( n27479 , n9429 , n27399 );
and ( n27480 , n27478 , n27479 );
xor ( n27481 , n27478 , n27479 );
xor ( n27482 , n26414 , n26615 );
nor ( n27483 , n8949 , n27399 );
and ( n27484 , n27482 , n27483 );
xor ( n27485 , n27482 , n27483 );
xor ( n27486 , n26418 , n26613 );
nor ( n27487 , n9437 , n27399 );
and ( n27488 , n27486 , n27487 );
xor ( n27489 , n27486 , n27487 );
xor ( n27490 , n26422 , n26611 );
nor ( n27491 , n9446 , n27399 );
and ( n27492 , n27490 , n27491 );
xor ( n27493 , n27490 , n27491 );
xor ( n27494 , n26426 , n26609 );
nor ( n27495 , n9455 , n27399 );
and ( n27496 , n27494 , n27495 );
xor ( n27497 , n27494 , n27495 );
xor ( n27498 , n26430 , n26607 );
nor ( n27499 , n9464 , n27399 );
and ( n27500 , n27498 , n27499 );
xor ( n27501 , n27498 , n27499 );
xor ( n27502 , n26434 , n26605 );
nor ( n27503 , n9473 , n27399 );
and ( n27504 , n27502 , n27503 );
xor ( n27505 , n27502 , n27503 );
xor ( n27506 , n26438 , n26603 );
nor ( n27507 , n9482 , n27399 );
and ( n27508 , n27506 , n27507 );
xor ( n27509 , n27506 , n27507 );
xor ( n27510 , n26442 , n26601 );
nor ( n27511 , n9491 , n27399 );
and ( n27512 , n27510 , n27511 );
xor ( n27513 , n27510 , n27511 );
xor ( n27514 , n26446 , n26599 );
nor ( n27515 , n9500 , n27399 );
and ( n27516 , n27514 , n27515 );
xor ( n27517 , n27514 , n27515 );
xor ( n27518 , n26450 , n26597 );
nor ( n27519 , n9509 , n27399 );
and ( n27520 , n27518 , n27519 );
xor ( n27521 , n27518 , n27519 );
xor ( n27522 , n26454 , n26595 );
nor ( n27523 , n9518 , n27399 );
and ( n27524 , n27522 , n27523 );
xor ( n27525 , n27522 , n27523 );
xor ( n27526 , n26458 , n26593 );
nor ( n27527 , n9527 , n27399 );
and ( n27528 , n27526 , n27527 );
xor ( n27529 , n27526 , n27527 );
xor ( n27530 , n26462 , n26591 );
nor ( n27531 , n9536 , n27399 );
and ( n27532 , n27530 , n27531 );
xor ( n27533 , n27530 , n27531 );
xor ( n27534 , n26466 , n26589 );
nor ( n27535 , n9545 , n27399 );
and ( n27536 , n27534 , n27535 );
xor ( n27537 , n27534 , n27535 );
xor ( n27538 , n26470 , n26587 );
nor ( n27539 , n9554 , n27399 );
and ( n27540 , n27538 , n27539 );
xor ( n27541 , n27538 , n27539 );
xor ( n27542 , n26474 , n26585 );
nor ( n27543 , n9563 , n27399 );
and ( n27544 , n27542 , n27543 );
xor ( n27545 , n27542 , n27543 );
xor ( n27546 , n26478 , n26583 );
nor ( n27547 , n9572 , n27399 );
and ( n27548 , n27546 , n27547 );
xor ( n27549 , n27546 , n27547 );
xor ( n27550 , n26482 , n26581 );
nor ( n27551 , n9581 , n27399 );
and ( n27552 , n27550 , n27551 );
xor ( n27553 , n27550 , n27551 );
xor ( n27554 , n26486 , n26579 );
nor ( n27555 , n9590 , n27399 );
and ( n27556 , n27554 , n27555 );
xor ( n27557 , n27554 , n27555 );
xor ( n27558 , n26490 , n26577 );
nor ( n27559 , n9599 , n27399 );
and ( n27560 , n27558 , n27559 );
xor ( n27561 , n27558 , n27559 );
xor ( n27562 , n26494 , n26575 );
nor ( n27563 , n9608 , n27399 );
and ( n27564 , n27562 , n27563 );
xor ( n27565 , n27562 , n27563 );
xor ( n27566 , n26498 , n26573 );
nor ( n27567 , n9617 , n27399 );
and ( n27568 , n27566 , n27567 );
xor ( n27569 , n27566 , n27567 );
xor ( n27570 , n26502 , n26571 );
nor ( n27571 , n9626 , n27399 );
and ( n27572 , n27570 , n27571 );
xor ( n27573 , n27570 , n27571 );
xor ( n27574 , n26506 , n26569 );
nor ( n27575 , n9635 , n27399 );
and ( n27576 , n27574 , n27575 );
xor ( n27577 , n27574 , n27575 );
xor ( n27578 , n26510 , n26567 );
nor ( n27579 , n9644 , n27399 );
and ( n27580 , n27578 , n27579 );
xor ( n27581 , n27578 , n27579 );
xor ( n27582 , n26514 , n26565 );
nor ( n27583 , n9653 , n27399 );
and ( n27584 , n27582 , n27583 );
xor ( n27585 , n27582 , n27583 );
xor ( n27586 , n26518 , n26563 );
nor ( n27587 , n9662 , n27399 );
and ( n27588 , n27586 , n27587 );
xor ( n27589 , n27586 , n27587 );
xor ( n27590 , n26522 , n26561 );
nor ( n27591 , n9671 , n27399 );
and ( n27592 , n27590 , n27591 );
xor ( n27593 , n27590 , n27591 );
xor ( n27594 , n26526 , n26559 );
nor ( n27595 , n9680 , n27399 );
and ( n27596 , n27594 , n27595 );
xor ( n27597 , n27594 , n27595 );
xor ( n27598 , n26530 , n26557 );
nor ( n27599 , n9689 , n27399 );
and ( n27600 , n27598 , n27599 );
xor ( n27601 , n27598 , n27599 );
xor ( n27602 , n26534 , n26555 );
nor ( n27603 , n9698 , n27399 );
and ( n27604 , n27602 , n27603 );
xor ( n27605 , n27602 , n27603 );
xor ( n27606 , n26538 , n26553 );
nor ( n27607 , n9707 , n27399 );
and ( n27608 , n27606 , n27607 );
xor ( n27609 , n27606 , n27607 );
xor ( n27610 , n26542 , n26551 );
nor ( n27611 , n9716 , n27399 );
and ( n27612 , n27610 , n27611 );
xor ( n27613 , n27610 , n27611 );
xor ( n27614 , n26546 , n26549 );
nor ( n27615 , n9725 , n27399 );
and ( n27616 , n27614 , n27615 );
xor ( n27617 , n27614 , n27615 );
xor ( n27618 , n26547 , n26548 );
nor ( n27619 , n9734 , n27399 );
and ( n27620 , n27618 , n27619 );
xor ( n27621 , n27618 , n27619 );
nor ( n27622 , n9752 , n26328 );
nor ( n27623 , n9743 , n27399 );
and ( n27624 , n27622 , n27623 );
and ( n27625 , n27621 , n27624 );
or ( n27626 , n27620 , n27625 );
and ( n27627 , n27617 , n27626 );
or ( n27628 , n27616 , n27627 );
and ( n27629 , n27613 , n27628 );
or ( n27630 , n27612 , n27629 );
and ( n27631 , n27609 , n27630 );
or ( n27632 , n27608 , n27631 );
and ( n27633 , n27605 , n27632 );
or ( n27634 , n27604 , n27633 );
and ( n27635 , n27601 , n27634 );
or ( n27636 , n27600 , n27635 );
and ( n27637 , n27597 , n27636 );
or ( n27638 , n27596 , n27637 );
and ( n27639 , n27593 , n27638 );
or ( n27640 , n27592 , n27639 );
and ( n27641 , n27589 , n27640 );
or ( n27642 , n27588 , n27641 );
and ( n27643 , n27585 , n27642 );
or ( n27644 , n27584 , n27643 );
and ( n27645 , n27581 , n27644 );
or ( n27646 , n27580 , n27645 );
and ( n27647 , n27577 , n27646 );
or ( n27648 , n27576 , n27647 );
and ( n27649 , n27573 , n27648 );
or ( n27650 , n27572 , n27649 );
and ( n27651 , n27569 , n27650 );
or ( n27652 , n27568 , n27651 );
and ( n27653 , n27565 , n27652 );
or ( n27654 , n27564 , n27653 );
and ( n27655 , n27561 , n27654 );
or ( n27656 , n27560 , n27655 );
and ( n27657 , n27557 , n27656 );
or ( n27658 , n27556 , n27657 );
and ( n27659 , n27553 , n27658 );
or ( n27660 , n27552 , n27659 );
and ( n27661 , n27549 , n27660 );
or ( n27662 , n27548 , n27661 );
and ( n27663 , n27545 , n27662 );
or ( n27664 , n27544 , n27663 );
and ( n27665 , n27541 , n27664 );
or ( n27666 , n27540 , n27665 );
and ( n27667 , n27537 , n27666 );
or ( n27668 , n27536 , n27667 );
and ( n27669 , n27533 , n27668 );
or ( n27670 , n27532 , n27669 );
and ( n27671 , n27529 , n27670 );
or ( n27672 , n27528 , n27671 );
and ( n27673 , n27525 , n27672 );
or ( n27674 , n27524 , n27673 );
and ( n27675 , n27521 , n27674 );
or ( n27676 , n27520 , n27675 );
and ( n27677 , n27517 , n27676 );
or ( n27678 , n27516 , n27677 );
and ( n27679 , n27513 , n27678 );
or ( n27680 , n27512 , n27679 );
and ( n27681 , n27509 , n27680 );
or ( n27682 , n27508 , n27681 );
and ( n27683 , n27505 , n27682 );
or ( n27684 , n27504 , n27683 );
and ( n27685 , n27501 , n27684 );
or ( n27686 , n27500 , n27685 );
and ( n27687 , n27497 , n27686 );
or ( n27688 , n27496 , n27687 );
and ( n27689 , n27493 , n27688 );
or ( n27690 , n27492 , n27689 );
and ( n27691 , n27489 , n27690 );
or ( n27692 , n27488 , n27691 );
and ( n27693 , n27485 , n27692 );
or ( n27694 , n27484 , n27693 );
and ( n27695 , n27481 , n27694 );
or ( n27696 , n27480 , n27695 );
and ( n27697 , n27477 , n27696 );
or ( n27698 , n27476 , n27697 );
and ( n27699 , n27473 , n27698 );
or ( n27700 , n27472 , n27699 );
and ( n27701 , n27469 , n27700 );
or ( n27702 , n27468 , n27701 );
and ( n27703 , n27465 , n27702 );
or ( n27704 , n27464 , n27703 );
and ( n27705 , n27461 , n27704 );
or ( n27706 , n27460 , n27705 );
and ( n27707 , n27457 , n27706 );
or ( n27708 , n27456 , n27707 );
and ( n27709 , n27453 , n27708 );
or ( n27710 , n27452 , n27709 );
and ( n27711 , n27449 , n27710 );
or ( n27712 , n27448 , n27711 );
and ( n27713 , n27445 , n27712 );
or ( n27714 , n27444 , n27713 );
and ( n27715 , n27441 , n27714 );
or ( n27716 , n27440 , n27715 );
and ( n27717 , n27437 , n27716 );
or ( n27718 , n27436 , n27717 );
and ( n27719 , n27433 , n27718 );
or ( n27720 , n27432 , n27719 );
and ( n27721 , n27429 , n27720 );
or ( n27722 , n27428 , n27721 );
and ( n27723 , n27425 , n27722 );
or ( n27724 , n27424 , n27723 );
and ( n27725 , n27421 , n27724 );
or ( n27726 , n27420 , n27725 );
and ( n27727 , n27417 , n27726 );
or ( n27728 , n27416 , n27727 );
and ( n27729 , n27413 , n27728 );
or ( n27730 , n27412 , n27729 );
and ( n27731 , n27409 , n27730 );
or ( n27732 , n27408 , n27731 );
and ( n27733 , n27405 , n27732 );
or ( n27734 , n27404 , n27733 );
xor ( n27735 , n27401 , n27734 );
buf ( n27736 , n476 );
not ( n27737 , n27736 );
nor ( n27738 , n601 , n27737 );
buf ( n27739 , n27738 );
nor ( n27740 , n622 , n25600 );
xor ( n27741 , n27739 , n27740 );
buf ( n27742 , n27741 );
nor ( n27743 , n646 , n24564 );
xor ( n27744 , n27742 , n27743 );
and ( n27745 , n26662 , n26663 );
buf ( n27746 , n27745 );
xor ( n27747 , n27744 , n27746 );
nor ( n27748 , n684 , n23541 );
xor ( n27749 , n27747 , n27748 );
and ( n27750 , n26665 , n26666 );
and ( n27751 , n26667 , n26669 );
or ( n27752 , n27750 , n27751 );
xor ( n27753 , n27749 , n27752 );
nor ( n27754 , n733 , n22541 );
xor ( n27755 , n27753 , n27754 );
and ( n27756 , n26670 , n26671 );
and ( n27757 , n26672 , n26675 );
or ( n27758 , n27756 , n27757 );
xor ( n27759 , n27755 , n27758 );
nor ( n27760 , n796 , n21562 );
xor ( n27761 , n27759 , n27760 );
and ( n27762 , n26676 , n26677 );
and ( n27763 , n26678 , n26681 );
or ( n27764 , n27762 , n27763 );
xor ( n27765 , n27761 , n27764 );
nor ( n27766 , n868 , n20601 );
xor ( n27767 , n27765 , n27766 );
and ( n27768 , n26682 , n26683 );
and ( n27769 , n26684 , n26687 );
or ( n27770 , n27768 , n27769 );
xor ( n27771 , n27767 , n27770 );
nor ( n27772 , n958 , n19657 );
xor ( n27773 , n27771 , n27772 );
and ( n27774 , n26688 , n26689 );
and ( n27775 , n26690 , n26693 );
or ( n27776 , n27774 , n27775 );
xor ( n27777 , n27773 , n27776 );
nor ( n27778 , n1062 , n18734 );
xor ( n27779 , n27777 , n27778 );
and ( n27780 , n26694 , n26695 );
and ( n27781 , n26696 , n26699 );
or ( n27782 , n27780 , n27781 );
xor ( n27783 , n27779 , n27782 );
nor ( n27784 , n1176 , n17828 );
xor ( n27785 , n27783 , n27784 );
and ( n27786 , n26700 , n26701 );
and ( n27787 , n26702 , n26705 );
or ( n27788 , n27786 , n27787 );
xor ( n27789 , n27785 , n27788 );
nor ( n27790 , n1303 , n16943 );
xor ( n27791 , n27789 , n27790 );
and ( n27792 , n26706 , n26707 );
and ( n27793 , n26708 , n26711 );
or ( n27794 , n27792 , n27793 );
xor ( n27795 , n27791 , n27794 );
nor ( n27796 , n1445 , n16077 );
xor ( n27797 , n27795 , n27796 );
and ( n27798 , n26712 , n26713 );
and ( n27799 , n26714 , n26717 );
or ( n27800 , n27798 , n27799 );
xor ( n27801 , n27797 , n27800 );
nor ( n27802 , n1598 , n15230 );
xor ( n27803 , n27801 , n27802 );
and ( n27804 , n26718 , n26719 );
and ( n27805 , n26720 , n26723 );
or ( n27806 , n27804 , n27805 );
xor ( n27807 , n27803 , n27806 );
nor ( n27808 , n1766 , n14403 );
xor ( n27809 , n27807 , n27808 );
and ( n27810 , n26724 , n26725 );
and ( n27811 , n26726 , n26729 );
or ( n27812 , n27810 , n27811 );
xor ( n27813 , n27809 , n27812 );
nor ( n27814 , n1945 , n13599 );
xor ( n27815 , n27813 , n27814 );
and ( n27816 , n26730 , n26731 );
and ( n27817 , n26732 , n26735 );
or ( n27818 , n27816 , n27817 );
xor ( n27819 , n27815 , n27818 );
nor ( n27820 , n2137 , n12808 );
xor ( n27821 , n27819 , n27820 );
and ( n27822 , n26736 , n26737 );
and ( n27823 , n26738 , n26741 );
or ( n27824 , n27822 , n27823 );
xor ( n27825 , n27821 , n27824 );
nor ( n27826 , n2343 , n12037 );
xor ( n27827 , n27825 , n27826 );
and ( n27828 , n26742 , n26743 );
and ( n27829 , n26744 , n26747 );
or ( n27830 , n27828 , n27829 );
xor ( n27831 , n27827 , n27830 );
nor ( n27832 , n2566 , n11282 );
xor ( n27833 , n27831 , n27832 );
and ( n27834 , n26748 , n26749 );
and ( n27835 , n26750 , n26753 );
or ( n27836 , n27834 , n27835 );
xor ( n27837 , n27833 , n27836 );
nor ( n27838 , n2797 , n10547 );
xor ( n27839 , n27837 , n27838 );
and ( n27840 , n26754 , n26755 );
and ( n27841 , n26756 , n26759 );
or ( n27842 , n27840 , n27841 );
xor ( n27843 , n27839 , n27842 );
nor ( n27844 , n3043 , n9829 );
xor ( n27845 , n27843 , n27844 );
and ( n27846 , n26760 , n26761 );
and ( n27847 , n26762 , n26765 );
or ( n27848 , n27846 , n27847 );
xor ( n27849 , n27845 , n27848 );
nor ( n27850 , n3300 , n8955 );
xor ( n27851 , n27849 , n27850 );
and ( n27852 , n26766 , n26767 );
and ( n27853 , n26768 , n26771 );
or ( n27854 , n27852 , n27853 );
xor ( n27855 , n27851 , n27854 );
nor ( n27856 , n3570 , n603 );
xor ( n27857 , n27855 , n27856 );
and ( n27858 , n26772 , n26773 );
and ( n27859 , n26774 , n26777 );
or ( n27860 , n27858 , n27859 );
xor ( n27861 , n27857 , n27860 );
nor ( n27862 , n3853 , n652 );
xor ( n27863 , n27861 , n27862 );
and ( n27864 , n26778 , n26779 );
and ( n27865 , n26780 , n26783 );
or ( n27866 , n27864 , n27865 );
xor ( n27867 , n27863 , n27866 );
nor ( n27868 , n4151 , n624 );
xor ( n27869 , n27867 , n27868 );
and ( n27870 , n26784 , n26785 );
and ( n27871 , n26786 , n26789 );
or ( n27872 , n27870 , n27871 );
xor ( n27873 , n27869 , n27872 );
nor ( n27874 , n4458 , n648 );
xor ( n27875 , n27873 , n27874 );
and ( n27876 , n26790 , n26791 );
and ( n27877 , n26792 , n26795 );
or ( n27878 , n27876 , n27877 );
xor ( n27879 , n27875 , n27878 );
nor ( n27880 , n4786 , n686 );
xor ( n27881 , n27879 , n27880 );
and ( n27882 , n26796 , n26797 );
and ( n27883 , n26798 , n26801 );
or ( n27884 , n27882 , n27883 );
xor ( n27885 , n27881 , n27884 );
nor ( n27886 , n5126 , n735 );
xor ( n27887 , n27885 , n27886 );
and ( n27888 , n26802 , n26803 );
and ( n27889 , n26804 , n26807 );
or ( n27890 , n27888 , n27889 );
xor ( n27891 , n27887 , n27890 );
nor ( n27892 , n5477 , n798 );
xor ( n27893 , n27891 , n27892 );
and ( n27894 , n26808 , n26809 );
and ( n27895 , n26810 , n26813 );
or ( n27896 , n27894 , n27895 );
xor ( n27897 , n27893 , n27896 );
nor ( n27898 , n5838 , n870 );
xor ( n27899 , n27897 , n27898 );
and ( n27900 , n26814 , n26815 );
and ( n27901 , n26816 , n26819 );
or ( n27902 , n27900 , n27901 );
xor ( n27903 , n27899 , n27902 );
nor ( n27904 , n6212 , n960 );
xor ( n27905 , n27903 , n27904 );
and ( n27906 , n26820 , n26821 );
and ( n27907 , n26822 , n26825 );
or ( n27908 , n27906 , n27907 );
xor ( n27909 , n27905 , n27908 );
nor ( n27910 , n6596 , n1064 );
xor ( n27911 , n27909 , n27910 );
and ( n27912 , n26826 , n26827 );
and ( n27913 , n26828 , n26831 );
or ( n27914 , n27912 , n27913 );
xor ( n27915 , n27911 , n27914 );
nor ( n27916 , n6997 , n1178 );
xor ( n27917 , n27915 , n27916 );
and ( n27918 , n26832 , n26833 );
and ( n27919 , n26834 , n26837 );
or ( n27920 , n27918 , n27919 );
xor ( n27921 , n27917 , n27920 );
nor ( n27922 , n7413 , n1305 );
xor ( n27923 , n27921 , n27922 );
and ( n27924 , n26838 , n26839 );
and ( n27925 , n26840 , n26843 );
or ( n27926 , n27924 , n27925 );
xor ( n27927 , n27923 , n27926 );
nor ( n27928 , n7841 , n1447 );
xor ( n27929 , n27927 , n27928 );
and ( n27930 , n26844 , n26845 );
and ( n27931 , n26846 , n26849 );
or ( n27932 , n27930 , n27931 );
xor ( n27933 , n27929 , n27932 );
nor ( n27934 , n8281 , n1600 );
xor ( n27935 , n27933 , n27934 );
and ( n27936 , n26850 , n26851 );
and ( n27937 , n26852 , n26855 );
or ( n27938 , n27936 , n27937 );
xor ( n27939 , n27935 , n27938 );
nor ( n27940 , n8737 , n1768 );
xor ( n27941 , n27939 , n27940 );
and ( n27942 , n26856 , n26857 );
and ( n27943 , n26858 , n26861 );
or ( n27944 , n27942 , n27943 );
xor ( n27945 , n27941 , n27944 );
nor ( n27946 , n9420 , n1947 );
xor ( n27947 , n27945 , n27946 );
and ( n27948 , n26862 , n26863 );
and ( n27949 , n26864 , n26867 );
or ( n27950 , n27948 , n27949 );
xor ( n27951 , n27947 , n27950 );
nor ( n27952 , n10312 , n2139 );
xor ( n27953 , n27951 , n27952 );
and ( n27954 , n26868 , n26869 );
and ( n27955 , n26870 , n26873 );
or ( n27956 , n27954 , n27955 );
xor ( n27957 , n27953 , n27956 );
nor ( n27958 , n11041 , n2345 );
xor ( n27959 , n27957 , n27958 );
and ( n27960 , n26874 , n26875 );
and ( n27961 , n26876 , n26879 );
or ( n27962 , n27960 , n27961 );
xor ( n27963 , n27959 , n27962 );
nor ( n27964 , n11790 , n2568 );
xor ( n27965 , n27963 , n27964 );
and ( n27966 , n26880 , n26881 );
and ( n27967 , n26882 , n26885 );
or ( n27968 , n27966 , n27967 );
xor ( n27969 , n27965 , n27968 );
nor ( n27970 , n12555 , n2799 );
xor ( n27971 , n27969 , n27970 );
and ( n27972 , n26886 , n26887 );
and ( n27973 , n26888 , n26891 );
or ( n27974 , n27972 , n27973 );
xor ( n27975 , n27971 , n27974 );
nor ( n27976 , n13340 , n3045 );
xor ( n27977 , n27975 , n27976 );
and ( n27978 , n26892 , n26893 );
and ( n27979 , n26894 , n26897 );
or ( n27980 , n27978 , n27979 );
xor ( n27981 , n27977 , n27980 );
nor ( n27982 , n14138 , n3302 );
xor ( n27983 , n27981 , n27982 );
and ( n27984 , n26898 , n26899 );
and ( n27985 , n26900 , n26903 );
or ( n27986 , n27984 , n27985 );
xor ( n27987 , n27983 , n27986 );
nor ( n27988 , n14959 , n3572 );
xor ( n27989 , n27987 , n27988 );
and ( n27990 , n26904 , n26905 );
and ( n27991 , n26906 , n26909 );
or ( n27992 , n27990 , n27991 );
xor ( n27993 , n27989 , n27992 );
nor ( n27994 , n15800 , n3855 );
xor ( n27995 , n27993 , n27994 );
and ( n27996 , n26910 , n26911 );
and ( n27997 , n26912 , n26915 );
or ( n27998 , n27996 , n27997 );
xor ( n27999 , n27995 , n27998 );
nor ( n28000 , n16660 , n4153 );
xor ( n28001 , n27999 , n28000 );
and ( n28002 , n26916 , n26917 );
and ( n28003 , n26918 , n26921 );
or ( n28004 , n28002 , n28003 );
xor ( n28005 , n28001 , n28004 );
nor ( n28006 , n17539 , n4460 );
xor ( n28007 , n28005 , n28006 );
and ( n28008 , n26922 , n26923 );
and ( n28009 , n26924 , n26927 );
or ( n28010 , n28008 , n28009 );
xor ( n28011 , n28007 , n28010 );
nor ( n28012 , n18439 , n4788 );
xor ( n28013 , n28011 , n28012 );
and ( n28014 , n26928 , n26929 );
and ( n28015 , n26930 , n26933 );
or ( n28016 , n28014 , n28015 );
xor ( n28017 , n28013 , n28016 );
nor ( n28018 , n19356 , n5128 );
xor ( n28019 , n28017 , n28018 );
and ( n28020 , n26934 , n26935 );
and ( n28021 , n26936 , n26939 );
or ( n28022 , n28020 , n28021 );
xor ( n28023 , n28019 , n28022 );
nor ( n28024 , n20294 , n5479 );
xor ( n28025 , n28023 , n28024 );
and ( n28026 , n26940 , n26941 );
and ( n28027 , n26942 , n26945 );
or ( n28028 , n28026 , n28027 );
xor ( n28029 , n28025 , n28028 );
nor ( n28030 , n21249 , n5840 );
xor ( n28031 , n28029 , n28030 );
and ( n28032 , n26946 , n26947 );
and ( n28033 , n26948 , n26951 );
or ( n28034 , n28032 , n28033 );
xor ( n28035 , n28031 , n28034 );
nor ( n28036 , n22222 , n6214 );
xor ( n28037 , n28035 , n28036 );
and ( n28038 , n26952 , n26953 );
and ( n28039 , n26954 , n26957 );
or ( n28040 , n28038 , n28039 );
xor ( n28041 , n28037 , n28040 );
nor ( n28042 , n23216 , n6598 );
xor ( n28043 , n28041 , n28042 );
and ( n28044 , n26958 , n26959 );
and ( n28045 , n26960 , n26963 );
or ( n28046 , n28044 , n28045 );
xor ( n28047 , n28043 , n28046 );
nor ( n28048 , n24233 , n6999 );
xor ( n28049 , n28047 , n28048 );
and ( n28050 , n26964 , n26965 );
and ( n28051 , n26966 , n26969 );
or ( n28052 , n28050 , n28051 );
xor ( n28053 , n28049 , n28052 );
nor ( n28054 , n25263 , n7415 );
xor ( n28055 , n28053 , n28054 );
and ( n28056 , n26970 , n26971 );
and ( n28057 , n26972 , n26975 );
or ( n28058 , n28056 , n28057 );
xor ( n28059 , n28055 , n28058 );
nor ( n28060 , n26317 , n7843 );
xor ( n28061 , n28059 , n28060 );
and ( n28062 , n26976 , n26977 );
and ( n28063 , n26978 , n26981 );
or ( n28064 , n28062 , n28063 );
xor ( n28065 , n28061 , n28064 );
nor ( n28066 , n27388 , n8283 );
xor ( n28067 , n28065 , n28066 );
and ( n28068 , n26982 , n26983 );
and ( n28069 , n26984 , n26987 );
or ( n28070 , n28068 , n28069 );
xor ( n28071 , n28067 , n28070 );
and ( n28072 , n27339 , n27340 );
and ( n28073 , n27340 , n27373 );
and ( n28074 , n27339 , n27373 );
or ( n28075 , n28072 , n28073 , n28074 );
and ( n28076 , n27001 , n27334 );
and ( n28077 , n27334 , n27374 );
and ( n28078 , n27001 , n27374 );
or ( n28079 , n28076 , n28077 , n28078 );
xor ( n28080 , n28075 , n28079 );
and ( n28081 , n27005 , n27125 );
and ( n28082 , n27125 , n27333 );
and ( n28083 , n27005 , n27333 );
or ( n28084 , n28081 , n28082 , n28083 );
and ( n28085 , n27130 , n27208 );
and ( n28086 , n27208 , n27332 );
and ( n28087 , n27130 , n27332 );
or ( n28088 , n28085 , n28086 , n28087 );
and ( n28089 , n27018 , n27086 );
and ( n28090 , n27086 , n27123 );
and ( n28091 , n27018 , n27123 );
or ( n28092 , n28089 , n28090 , n28091 );
and ( n28093 , n27134 , n27138 );
and ( n28094 , n27138 , n27207 );
and ( n28095 , n27134 , n27207 );
or ( n28096 , n28093 , n28094 , n28095 );
xor ( n28097 , n28092 , n28096 );
and ( n28098 , n27091 , n27095 );
and ( n28099 , n27095 , n27122 );
and ( n28100 , n27091 , n27122 );
or ( n28101 , n28098 , n28099 , n28100 );
and ( n28102 , n27052 , n27068 );
and ( n28103 , n27068 , n27084 );
and ( n28104 , n27052 , n27084 );
or ( n28105 , n28102 , n28103 , n28104 );
and ( n28106 , n27035 , n27039 );
and ( n28107 , n27039 , n27045 );
and ( n28108 , n27035 , n27045 );
or ( n28109 , n28106 , n28107 , n28108 );
and ( n28110 , n27056 , n27061 );
and ( n28111 , n27061 , n27067 );
and ( n28112 , n27056 , n27067 );
or ( n28113 , n28110 , n28111 , n28112 );
xor ( n28114 , n28109 , n28113 );
and ( n28115 , n27041 , n27042 );
and ( n28116 , n27042 , n27044 );
and ( n28117 , n27041 , n27044 );
or ( n28118 , n28115 , n28116 , n28117 );
and ( n28119 , n27057 , n27058 );
and ( n28120 , n27058 , n27060 );
and ( n28121 , n27057 , n27060 );
or ( n28122 , n28119 , n28120 , n28121 );
xor ( n28123 , n28118 , n28122 );
and ( n28124 , n21216 , n840 );
and ( n28125 , n22186 , n771 );
xor ( n28126 , n28124 , n28125 );
and ( n28127 , n22892 , n719 );
xor ( n28128 , n28126 , n28127 );
xor ( n28129 , n28123 , n28128 );
xor ( n28130 , n28114 , n28129 );
xor ( n28131 , n28105 , n28130 );
and ( n28132 , n27073 , n27077 );
and ( n28133 , n27077 , n27083 );
and ( n28134 , n27073 , n27083 );
or ( n28135 , n28132 , n28133 , n28134 );
and ( n28136 , n27063 , n27064 );
and ( n28137 , n27064 , n27066 );
and ( n28138 , n27063 , n27066 );
or ( n28139 , n28136 , n28137 , n28138 );
and ( n28140 , n18144 , n1134 );
and ( n28141 , n19324 , n1034 );
xor ( n28142 , n28140 , n28141 );
and ( n28143 , n20233 , n940 );
xor ( n28144 , n28142 , n28143 );
xor ( n28145 , n28139 , n28144 );
and ( n28146 , n15758 , n1551 );
and ( n28147 , n16637 , n1424 );
xor ( n28148 , n28146 , n28147 );
and ( n28149 , n17512 , n1254 );
xor ( n28150 , n28148 , n28149 );
xor ( n28151 , n28145 , n28150 );
xor ( n28152 , n28135 , n28151 );
and ( n28153 , n27079 , n27080 );
and ( n28154 , n27080 , n27082 );
and ( n28155 , n27079 , n27082 );
or ( n28156 , n28153 , n28154 , n28155 );
and ( n28157 , n27110 , n27111 );
and ( n28158 , n27111 , n27113 );
and ( n28159 , n27110 , n27113 );
or ( n28160 , n28157 , n28158 , n28159 );
xor ( n28161 , n28156 , n28160 );
and ( n28162 , n13322 , n2100 );
and ( n28163 , n14118 , n1882 );
xor ( n28164 , n28162 , n28163 );
and ( n28165 , n14938 , n1738 );
xor ( n28166 , n28164 , n28165 );
xor ( n28167 , n28161 , n28166 );
xor ( n28168 , n28152 , n28167 );
xor ( n28169 , n28131 , n28168 );
xor ( n28170 , n28101 , n28169 );
and ( n28171 , n27100 , n27104 );
and ( n28172 , n27104 , n27121 );
and ( n28173 , n27100 , n27121 );
or ( n28174 , n28171 , n28172 , n28173 );
and ( n28175 , n27173 , n27188 );
and ( n28176 , n27188 , n27205 );
and ( n28177 , n27173 , n27205 );
or ( n28178 , n28175 , n28176 , n28177 );
xor ( n28179 , n28174 , n28178 );
and ( n28180 , n27109 , n27114 );
and ( n28181 , n27114 , n27120 );
and ( n28182 , n27109 , n27120 );
or ( n28183 , n28180 , n28181 , n28182 );
and ( n28184 , n27177 , n27181 );
and ( n28185 , n27181 , n27187 );
and ( n28186 , n27177 , n27187 );
or ( n28187 , n28184 , n28185 , n28186 );
xor ( n28188 , n28183 , n28187 );
and ( n28189 , n27116 , n27117 );
and ( n28190 , n27117 , n27119 );
and ( n28191 , n27116 , n27119 );
or ( n28192 , n28189 , n28190 , n28191 );
and ( n28193 , n11015 , n2739 );
and ( n28194 , n11769 , n2544 );
xor ( n28195 , n28193 , n28194 );
and ( n28196 , n12320 , n2298 );
xor ( n28197 , n28195 , n28196 );
xor ( n28198 , n28192 , n28197 );
and ( n28199 , n8718 , n3495 );
and ( n28200 , n9400 , n3271 );
xor ( n28201 , n28199 , n28200 );
and ( n28202 , n10291 , n2981 );
xor ( n28203 , n28201 , n28202 );
xor ( n28204 , n28198 , n28203 );
xor ( n28205 , n28188 , n28204 );
xor ( n28206 , n28179 , n28205 );
xor ( n28207 , n28170 , n28206 );
xor ( n28208 , n28097 , n28207 );
xor ( n28209 , n28088 , n28208 );
and ( n28210 , n27213 , n27260 );
and ( n28211 , n27260 , n27331 );
and ( n28212 , n27213 , n27331 );
or ( n28213 , n28210 , n28211 , n28212 );
and ( n28214 , n27143 , n27168 );
and ( n28215 , n27168 , n27206 );
and ( n28216 , n27143 , n27206 );
or ( n28217 , n28214 , n28215 , n28216 );
and ( n28218 , n27217 , n27221 );
and ( n28219 , n27221 , n27259 );
and ( n28220 , n27217 , n27259 );
or ( n28221 , n28218 , n28219 , n28220 );
xor ( n28222 , n28217 , n28221 );
and ( n28223 , n27147 , n27151 );
and ( n28224 , n27151 , n27167 );
and ( n28225 , n27147 , n27167 );
or ( n28226 , n28223 , n28224 , n28225 );
and ( n28227 , n27193 , n27198 );
and ( n28228 , n27198 , n27204 );
and ( n28229 , n27193 , n27204 );
or ( n28230 , n28227 , n28228 , n28229 );
and ( n28231 , n27183 , n27184 );
and ( n28232 , n27184 , n27186 );
and ( n28233 , n27183 , n27186 );
or ( n28234 , n28231 , n28232 , n28233 );
and ( n28235 , n27194 , n27195 );
and ( n28236 , n27195 , n27197 );
and ( n28237 , n27194 , n27197 );
or ( n28238 , n28235 , n28236 , n28237 );
xor ( n28239 , n28234 , n28238 );
and ( n28240 , n7385 , n4403 );
and ( n28241 , n7808 , n4102 );
xor ( n28242 , n28240 , n28241 );
and ( n28243 , n8079 , n3749 );
xor ( n28244 , n28242 , n28243 );
xor ( n28245 , n28239 , n28244 );
xor ( n28246 , n28230 , n28245 );
and ( n28247 , n27200 , n27201 );
and ( n28248 , n27201 , n27203 );
and ( n28249 , n27200 , n27203 );
or ( n28250 , n28247 , n28248 , n28249 );
and ( n28251 , n6187 , n5408 );
and ( n28252 , n6569 , n5103 );
xor ( n28253 , n28251 , n28252 );
and ( n28254 , n6816 , n4730 );
xor ( n28255 , n28253 , n28254 );
xor ( n28256 , n28250 , n28255 );
and ( n28257 , n4959 , n6504 );
and ( n28258 , n5459 , n6132 );
xor ( n28259 , n28257 , n28258 );
buf ( n28260 , n5819 );
xor ( n28261 , n28259 , n28260 );
xor ( n28262 , n28256 , n28261 );
xor ( n28263 , n28246 , n28262 );
xor ( n28264 , n28226 , n28263 );
and ( n28265 , n27156 , n27160 );
and ( n28266 , n27160 , n27166 );
and ( n28267 , n27156 , n27166 );
or ( n28268 , n28265 , n28266 , n28267 );
and ( n28269 , n27230 , n27235 );
and ( n28270 , n27235 , n27241 );
and ( n28271 , n27230 , n27241 );
or ( n28272 , n28269 , n28270 , n28271 );
xor ( n28273 , n28268 , n28272 );
and ( n28274 , n27162 , n27163 );
and ( n28275 , n27163 , n27165 );
and ( n28276 , n27162 , n27165 );
or ( n28277 , n28274 , n28275 , n28276 );
and ( n28278 , n27231 , n27232 );
and ( n28279 , n27232 , n27234 );
and ( n28280 , n27231 , n27234 );
or ( n28281 , n28278 , n28279 , n28280 );
xor ( n28282 , n28277 , n28281 );
and ( n28283 , n4132 , n7662 );
and ( n28284 , n4438 , n7310 );
xor ( n28285 , n28283 , n28284 );
and ( n28286 , n4766 , n6971 );
xor ( n28287 , n28285 , n28286 );
xor ( n28288 , n28282 , n28287 );
xor ( n28289 , n28273 , n28288 );
xor ( n28290 , n28264 , n28289 );
xor ( n28291 , n28222 , n28290 );
xor ( n28292 , n28213 , n28291 );
and ( n28293 , n27265 , n27303 );
and ( n28294 , n27303 , n27330 );
and ( n28295 , n27265 , n27330 );
or ( n28296 , n28293 , n28294 , n28295 );
and ( n28297 , n27308 , n27312 );
and ( n28298 , n27312 , n27329 );
and ( n28299 , n27308 , n27329 );
or ( n28300 , n28297 , n28298 , n28299 );
and ( n28301 , n27226 , n27242 );
and ( n28302 , n27242 , n27258 );
and ( n28303 , n27226 , n27258 );
or ( n28304 , n28301 , n28302 , n28303 );
xor ( n28305 , n28300 , n28304 );
and ( n28306 , n27247 , n27251 );
and ( n28307 , n27251 , n27257 );
and ( n28308 , n27247 , n27257 );
or ( n28309 , n28306 , n28307 , n28308 );
and ( n28310 , n27237 , n27238 );
and ( n28311 , n27238 , n27240 );
and ( n28312 , n27237 , n27240 );
or ( n28313 , n28310 , n28311 , n28312 );
and ( n28314 , n3182 , n9348 );
and ( n28315 , n3545 , n8669 );
xor ( n28316 , n28314 , n28315 );
and ( n28317 , n3801 , n8243 );
xor ( n28318 , n28316 , n28317 );
xor ( n28319 , n28313 , n28318 );
and ( n28320 , n2462 , n11718 );
and ( n28321 , n2779 , n10977 );
xor ( n28322 , n28320 , n28321 );
and ( n28323 , n3024 , n10239 );
xor ( n28324 , n28322 , n28323 );
xor ( n28325 , n28319 , n28324 );
xor ( n28326 , n28309 , n28325 );
and ( n28327 , n27253 , n27254 );
and ( n28328 , n27254 , n27256 );
and ( n28329 , n27253 , n27256 );
or ( n28330 , n28327 , n28328 , n28329 );
and ( n28331 , n27318 , n27319 );
and ( n28332 , n27319 , n27321 );
and ( n28333 , n27318 , n27321 );
or ( n28334 , n28331 , n28332 , n28333 );
xor ( n28335 , n28330 , n28334 );
and ( n28336 , n1933 , n14044 );
and ( n28337 , n2120 , n13256 );
xor ( n28338 , n28336 , n28337 );
and ( n28339 , n2324 , n12531 );
xor ( n28340 , n28338 , n28339 );
xor ( n28341 , n28335 , n28340 );
xor ( n28342 , n28326 , n28341 );
xor ( n28343 , n28305 , n28342 );
xor ( n28344 , n28296 , n28343 );
and ( n28345 , n27269 , n27284 );
and ( n28346 , n27284 , n27302 );
and ( n28347 , n27269 , n27302 );
or ( n28348 , n28345 , n28346 , n28347 );
and ( n28349 , n27317 , n27322 );
and ( n28350 , n27322 , n27328 );
and ( n28351 , n27317 , n27328 );
or ( n28352 , n28349 , n28350 , n28351 );
and ( n28353 , n27273 , n27277 );
and ( n28354 , n27277 , n27283 );
and ( n28355 , n27273 , n27283 );
or ( n28356 , n28353 , n28354 , n28355 );
xor ( n28357 , n28352 , n28356 );
and ( n28358 , n27324 , n27325 );
and ( n28359 , n27325 , n27327 );
and ( n28360 , n27324 , n27327 );
or ( n28361 , n28358 , n28359 , n28360 );
and ( n28362 , n1383 , n16550 );
and ( n28363 , n1580 , n15691 );
xor ( n28364 , n28362 , n28363 );
and ( n28365 , n1694 , n14838 );
xor ( n28366 , n28364 , n28365 );
xor ( n28367 , n28361 , n28366 );
and ( n28368 , n1047 , n19222 );
and ( n28369 , n1164 , n18407 );
xor ( n28370 , n28368 , n28369 );
and ( n28371 , n1287 , n17422 );
xor ( n28372 , n28370 , n28371 );
xor ( n28373 , n28367 , n28372 );
xor ( n28374 , n28357 , n28373 );
xor ( n28375 , n28348 , n28374 );
and ( n28376 , n27289 , n27294 );
and ( n28377 , n27294 , n27301 );
and ( n28378 , n27289 , n27301 );
or ( n28379 , n28376 , n28377 , n28378 );
and ( n28380 , n27279 , n27280 );
and ( n28381 , n27280 , n27282 );
and ( n28382 , n27279 , n27282 );
or ( n28383 , n28380 , n28381 , n28382 );
and ( n28384 , n27290 , n27291 );
and ( n28385 , n27291 , n27293 );
and ( n28386 , n27290 , n27293 );
or ( n28387 , n28384 , n28385 , n28386 );
xor ( n28388 , n28383 , n28387 );
and ( n28389 , n783 , n22065 );
and ( n28390 , n856 , n20976 );
xor ( n28391 , n28389 , n28390 );
and ( n28392 , n925 , n20156 );
xor ( n28393 , n28391 , n28392 );
xor ( n28394 , n28388 , n28393 );
xor ( n28395 , n28379 , n28394 );
and ( n28396 , n27297 , n27298 );
and ( n28397 , n27298 , n27300 );
and ( n28398 , n27297 , n27300 );
or ( n28399 , n28396 , n28397 , n28398 );
and ( n28400 , n632 , n25163 );
and ( n28401 , n671 , n24137 );
xor ( n28402 , n28400 , n28401 );
and ( n28403 , n715 , n23075 );
xor ( n28404 , n28402 , n28403 );
xor ( n28405 , n28399 , n28404 );
buf ( n28406 , n412 );
and ( n28407 , n599 , n28406 );
and ( n28408 , n608 , n27296 );
xor ( n28409 , n28407 , n28408 );
and ( n28410 , n611 , n26216 );
xor ( n28411 , n28409 , n28410 );
xor ( n28412 , n28405 , n28411 );
xor ( n28413 , n28395 , n28412 );
xor ( n28414 , n28375 , n28413 );
xor ( n28415 , n28344 , n28414 );
xor ( n28416 , n28292 , n28415 );
xor ( n28417 , n28209 , n28416 );
xor ( n28418 , n28084 , n28417 );
and ( n28419 , n27009 , n27013 );
and ( n28420 , n27013 , n27124 );
and ( n28421 , n27009 , n27124 );
or ( n28422 , n28419 , n28420 , n28421 );
and ( n28423 , n27345 , n27372 );
xor ( n28424 , n28422 , n28423 );
and ( n28425 , n27349 , n27350 );
and ( n28426 , n27350 , n27371 );
and ( n28427 , n27349 , n27371 );
or ( n28428 , n28425 , n28426 , n28427 );
and ( n28429 , n27022 , n27047 );
and ( n28430 , n27047 , n27085 );
and ( n28431 , n27022 , n27085 );
or ( n28432 , n28429 , n28430 , n28431 );
and ( n28433 , n27355 , n27370 );
xor ( n28434 , n28432 , n28433 );
and ( n28435 , n27026 , n27030 );
and ( n28436 , n27030 , n27046 );
and ( n28437 , n27026 , n27046 );
or ( n28438 , n28435 , n28436 , n28437 );
and ( n28439 , n27356 , n27369 );
xor ( n28440 , n28438 , n28439 );
and ( n28441 , n27360 , n27362 );
and ( n28442 , n27362 , n27368 );
and ( n28443 , n27360 , n27368 );
or ( n28444 , n28441 , n28442 , n28443 );
and ( n28445 , n27364 , n27365 );
and ( n28446 , n27365 , n27367 );
and ( n28447 , n27364 , n27367 );
or ( n28448 , n28445 , n28446 , n28447 );
and ( n28449 , n24214 , n663 );
and ( n28450 , n25243 , n635 );
xor ( n28451 , n28449 , n28450 );
and ( n28452 , n26296 , n606 );
xor ( n28453 , n28451 , n28452 );
xor ( n28454 , n28448 , n28453 );
and ( n28455 , n27361 , n615 );
buf ( n28456 , n412 );
and ( n28457 , n28456 , n612 );
xor ( n28458 , n28455 , n28457 );
xor ( n28459 , n28454 , n28458 );
xor ( n28460 , n28444 , n28459 );
xor ( n28461 , n28440 , n28460 );
xor ( n28462 , n28434 , n28461 );
xor ( n28463 , n28428 , n28462 );
xor ( n28464 , n28424 , n28463 );
xor ( n28465 , n28418 , n28464 );
xor ( n28466 , n28080 , n28465 );
and ( n28467 , n26992 , n26996 );
and ( n28468 , n26996 , n27375 );
and ( n28469 , n26992 , n27375 );
or ( n28470 , n28467 , n28468 , n28469 );
xor ( n28471 , n28466 , n28470 );
and ( n28472 , n27376 , n27380 );
and ( n28473 , n27381 , n27384 );
or ( n28474 , n28472 , n28473 );
xor ( n28475 , n28471 , n28474 );
buf ( n28476 , n28475 );
buf ( n28477 , n28476 );
not ( n28478 , n28477 );
nor ( n28479 , n28478 , n8739 );
xor ( n28480 , n28071 , n28479 );
and ( n28481 , n26988 , n27389 );
and ( n28482 , n27390 , n27393 );
or ( n28483 , n28481 , n28482 );
xor ( n28484 , n28480 , n28483 );
buf ( n28485 , n28484 );
buf ( n28486 , n28485 );
not ( n28487 , n28486 );
buf ( n28488 , n557 );
not ( n28489 , n28488 );
nor ( n28490 , n28487 , n28489 );
xor ( n28491 , n27735 , n28490 );
xor ( n28492 , n27405 , n27732 );
nor ( n28493 , n27397 , n28489 );
and ( n28494 , n28492 , n28493 );
xor ( n28495 , n28492 , n28493 );
xor ( n28496 , n27409 , n27730 );
nor ( n28497 , n26326 , n28489 );
and ( n28498 , n28496 , n28497 );
xor ( n28499 , n28496 , n28497 );
xor ( n28500 , n27413 , n27728 );
nor ( n28501 , n25272 , n28489 );
and ( n28502 , n28500 , n28501 );
xor ( n28503 , n28500 , n28501 );
xor ( n28504 , n27417 , n27726 );
nor ( n28505 , n24242 , n28489 );
and ( n28506 , n28504 , n28505 );
xor ( n28507 , n28504 , n28505 );
xor ( n28508 , n27421 , n27724 );
nor ( n28509 , n23225 , n28489 );
and ( n28510 , n28508 , n28509 );
xor ( n28511 , n28508 , n28509 );
xor ( n28512 , n27425 , n27722 );
nor ( n28513 , n22231 , n28489 );
and ( n28514 , n28512 , n28513 );
xor ( n28515 , n28512 , n28513 );
xor ( n28516 , n27429 , n27720 );
nor ( n28517 , n21258 , n28489 );
and ( n28518 , n28516 , n28517 );
xor ( n28519 , n28516 , n28517 );
xor ( n28520 , n27433 , n27718 );
nor ( n28521 , n20303 , n28489 );
and ( n28522 , n28520 , n28521 );
xor ( n28523 , n28520 , n28521 );
xor ( n28524 , n27437 , n27716 );
nor ( n28525 , n19365 , n28489 );
and ( n28526 , n28524 , n28525 );
xor ( n28527 , n28524 , n28525 );
xor ( n28528 , n27441 , n27714 );
nor ( n28529 , n18448 , n28489 );
and ( n28530 , n28528 , n28529 );
xor ( n28531 , n28528 , n28529 );
xor ( n28532 , n27445 , n27712 );
nor ( n28533 , n17548 , n28489 );
and ( n28534 , n28532 , n28533 );
xor ( n28535 , n28532 , n28533 );
xor ( n28536 , n27449 , n27710 );
nor ( n28537 , n16669 , n28489 );
and ( n28538 , n28536 , n28537 );
xor ( n28539 , n28536 , n28537 );
xor ( n28540 , n27453 , n27708 );
nor ( n28541 , n15809 , n28489 );
and ( n28542 , n28540 , n28541 );
xor ( n28543 , n28540 , n28541 );
xor ( n28544 , n27457 , n27706 );
nor ( n28545 , n14968 , n28489 );
and ( n28546 , n28544 , n28545 );
xor ( n28547 , n28544 , n28545 );
xor ( n28548 , n27461 , n27704 );
nor ( n28549 , n14147 , n28489 );
and ( n28550 , n28548 , n28549 );
xor ( n28551 , n28548 , n28549 );
xor ( n28552 , n27465 , n27702 );
nor ( n28553 , n13349 , n28489 );
and ( n28554 , n28552 , n28553 );
xor ( n28555 , n28552 , n28553 );
xor ( n28556 , n27469 , n27700 );
nor ( n28557 , n12564 , n28489 );
and ( n28558 , n28556 , n28557 );
xor ( n28559 , n28556 , n28557 );
xor ( n28560 , n27473 , n27698 );
nor ( n28561 , n11799 , n28489 );
and ( n28562 , n28560 , n28561 );
xor ( n28563 , n28560 , n28561 );
xor ( n28564 , n27477 , n27696 );
nor ( n28565 , n11050 , n28489 );
and ( n28566 , n28564 , n28565 );
xor ( n28567 , n28564 , n28565 );
xor ( n28568 , n27481 , n27694 );
nor ( n28569 , n10321 , n28489 );
and ( n28570 , n28568 , n28569 );
xor ( n28571 , n28568 , n28569 );
xor ( n28572 , n27485 , n27692 );
nor ( n28573 , n9429 , n28489 );
and ( n28574 , n28572 , n28573 );
xor ( n28575 , n28572 , n28573 );
xor ( n28576 , n27489 , n27690 );
nor ( n28577 , n8949 , n28489 );
and ( n28578 , n28576 , n28577 );
xor ( n28579 , n28576 , n28577 );
xor ( n28580 , n27493 , n27688 );
nor ( n28581 , n9437 , n28489 );
and ( n28582 , n28580 , n28581 );
xor ( n28583 , n28580 , n28581 );
xor ( n28584 , n27497 , n27686 );
nor ( n28585 , n9446 , n28489 );
and ( n28586 , n28584 , n28585 );
xor ( n28587 , n28584 , n28585 );
xor ( n28588 , n27501 , n27684 );
nor ( n28589 , n9455 , n28489 );
and ( n28590 , n28588 , n28589 );
xor ( n28591 , n28588 , n28589 );
xor ( n28592 , n27505 , n27682 );
nor ( n28593 , n9464 , n28489 );
and ( n28594 , n28592 , n28593 );
xor ( n28595 , n28592 , n28593 );
xor ( n28596 , n27509 , n27680 );
nor ( n28597 , n9473 , n28489 );
and ( n28598 , n28596 , n28597 );
xor ( n28599 , n28596 , n28597 );
xor ( n28600 , n27513 , n27678 );
nor ( n28601 , n9482 , n28489 );
and ( n28602 , n28600 , n28601 );
xor ( n28603 , n28600 , n28601 );
xor ( n28604 , n27517 , n27676 );
nor ( n28605 , n9491 , n28489 );
and ( n28606 , n28604 , n28605 );
xor ( n28607 , n28604 , n28605 );
xor ( n28608 , n27521 , n27674 );
nor ( n28609 , n9500 , n28489 );
and ( n28610 , n28608 , n28609 );
xor ( n28611 , n28608 , n28609 );
xor ( n28612 , n27525 , n27672 );
nor ( n28613 , n9509 , n28489 );
and ( n28614 , n28612 , n28613 );
xor ( n28615 , n28612 , n28613 );
xor ( n28616 , n27529 , n27670 );
nor ( n28617 , n9518 , n28489 );
and ( n28618 , n28616 , n28617 );
xor ( n28619 , n28616 , n28617 );
xor ( n28620 , n27533 , n27668 );
nor ( n28621 , n9527 , n28489 );
and ( n28622 , n28620 , n28621 );
xor ( n28623 , n28620 , n28621 );
xor ( n28624 , n27537 , n27666 );
nor ( n28625 , n9536 , n28489 );
and ( n28626 , n28624 , n28625 );
xor ( n28627 , n28624 , n28625 );
xor ( n28628 , n27541 , n27664 );
nor ( n28629 , n9545 , n28489 );
and ( n28630 , n28628 , n28629 );
xor ( n28631 , n28628 , n28629 );
xor ( n28632 , n27545 , n27662 );
nor ( n28633 , n9554 , n28489 );
and ( n28634 , n28632 , n28633 );
xor ( n28635 , n28632 , n28633 );
xor ( n28636 , n27549 , n27660 );
nor ( n28637 , n9563 , n28489 );
and ( n28638 , n28636 , n28637 );
xor ( n28639 , n28636 , n28637 );
xor ( n28640 , n27553 , n27658 );
nor ( n28641 , n9572 , n28489 );
and ( n28642 , n28640 , n28641 );
xor ( n28643 , n28640 , n28641 );
xor ( n28644 , n27557 , n27656 );
nor ( n28645 , n9581 , n28489 );
and ( n28646 , n28644 , n28645 );
xor ( n28647 , n28644 , n28645 );
xor ( n28648 , n27561 , n27654 );
nor ( n28649 , n9590 , n28489 );
and ( n28650 , n28648 , n28649 );
xor ( n28651 , n28648 , n28649 );
xor ( n28652 , n27565 , n27652 );
nor ( n28653 , n9599 , n28489 );
and ( n28654 , n28652 , n28653 );
xor ( n28655 , n28652 , n28653 );
xor ( n28656 , n27569 , n27650 );
nor ( n28657 , n9608 , n28489 );
and ( n28658 , n28656 , n28657 );
xor ( n28659 , n28656 , n28657 );
xor ( n28660 , n27573 , n27648 );
nor ( n28661 , n9617 , n28489 );
and ( n28662 , n28660 , n28661 );
xor ( n28663 , n28660 , n28661 );
xor ( n28664 , n27577 , n27646 );
nor ( n28665 , n9626 , n28489 );
and ( n28666 , n28664 , n28665 );
xor ( n28667 , n28664 , n28665 );
xor ( n28668 , n27581 , n27644 );
nor ( n28669 , n9635 , n28489 );
and ( n28670 , n28668 , n28669 );
xor ( n28671 , n28668 , n28669 );
xor ( n28672 , n27585 , n27642 );
nor ( n28673 , n9644 , n28489 );
and ( n28674 , n28672 , n28673 );
xor ( n28675 , n28672 , n28673 );
xor ( n28676 , n27589 , n27640 );
nor ( n28677 , n9653 , n28489 );
and ( n28678 , n28676 , n28677 );
xor ( n28679 , n28676 , n28677 );
xor ( n28680 , n27593 , n27638 );
nor ( n28681 , n9662 , n28489 );
and ( n28682 , n28680 , n28681 );
xor ( n28683 , n28680 , n28681 );
xor ( n28684 , n27597 , n27636 );
nor ( n28685 , n9671 , n28489 );
and ( n28686 , n28684 , n28685 );
xor ( n28687 , n28684 , n28685 );
xor ( n28688 , n27601 , n27634 );
nor ( n28689 , n9680 , n28489 );
and ( n28690 , n28688 , n28689 );
xor ( n28691 , n28688 , n28689 );
xor ( n28692 , n27605 , n27632 );
nor ( n28693 , n9689 , n28489 );
and ( n28694 , n28692 , n28693 );
xor ( n28695 , n28692 , n28693 );
xor ( n28696 , n27609 , n27630 );
nor ( n28697 , n9698 , n28489 );
and ( n28698 , n28696 , n28697 );
xor ( n28699 , n28696 , n28697 );
xor ( n28700 , n27613 , n27628 );
nor ( n28701 , n9707 , n28489 );
and ( n28702 , n28700 , n28701 );
xor ( n28703 , n28700 , n28701 );
xor ( n28704 , n27617 , n27626 );
nor ( n28705 , n9716 , n28489 );
and ( n28706 , n28704 , n28705 );
xor ( n28707 , n28704 , n28705 );
xor ( n28708 , n27621 , n27624 );
nor ( n28709 , n9725 , n28489 );
and ( n28710 , n28708 , n28709 );
xor ( n28711 , n28708 , n28709 );
xor ( n28712 , n27622 , n27623 );
nor ( n28713 , n9734 , n28489 );
and ( n28714 , n28712 , n28713 );
xor ( n28715 , n28712 , n28713 );
nor ( n28716 , n9752 , n27399 );
nor ( n28717 , n9743 , n28489 );
and ( n28718 , n28716 , n28717 );
and ( n28719 , n28715 , n28718 );
or ( n28720 , n28714 , n28719 );
and ( n28721 , n28711 , n28720 );
or ( n28722 , n28710 , n28721 );
and ( n28723 , n28707 , n28722 );
or ( n28724 , n28706 , n28723 );
and ( n28725 , n28703 , n28724 );
or ( n28726 , n28702 , n28725 );
and ( n28727 , n28699 , n28726 );
or ( n28728 , n28698 , n28727 );
and ( n28729 , n28695 , n28728 );
or ( n28730 , n28694 , n28729 );
and ( n28731 , n28691 , n28730 );
or ( n28732 , n28690 , n28731 );
and ( n28733 , n28687 , n28732 );
or ( n28734 , n28686 , n28733 );
and ( n28735 , n28683 , n28734 );
or ( n28736 , n28682 , n28735 );
and ( n28737 , n28679 , n28736 );
or ( n28738 , n28678 , n28737 );
and ( n28739 , n28675 , n28738 );
or ( n28740 , n28674 , n28739 );
and ( n28741 , n28671 , n28740 );
or ( n28742 , n28670 , n28741 );
and ( n28743 , n28667 , n28742 );
or ( n28744 , n28666 , n28743 );
and ( n28745 , n28663 , n28744 );
or ( n28746 , n28662 , n28745 );
and ( n28747 , n28659 , n28746 );
or ( n28748 , n28658 , n28747 );
and ( n28749 , n28655 , n28748 );
or ( n28750 , n28654 , n28749 );
and ( n28751 , n28651 , n28750 );
or ( n28752 , n28650 , n28751 );
and ( n28753 , n28647 , n28752 );
or ( n28754 , n28646 , n28753 );
and ( n28755 , n28643 , n28754 );
or ( n28756 , n28642 , n28755 );
and ( n28757 , n28639 , n28756 );
or ( n28758 , n28638 , n28757 );
and ( n28759 , n28635 , n28758 );
or ( n28760 , n28634 , n28759 );
and ( n28761 , n28631 , n28760 );
or ( n28762 , n28630 , n28761 );
and ( n28763 , n28627 , n28762 );
or ( n28764 , n28626 , n28763 );
and ( n28765 , n28623 , n28764 );
or ( n28766 , n28622 , n28765 );
and ( n28767 , n28619 , n28766 );
or ( n28768 , n28618 , n28767 );
and ( n28769 , n28615 , n28768 );
or ( n28770 , n28614 , n28769 );
and ( n28771 , n28611 , n28770 );
or ( n28772 , n28610 , n28771 );
and ( n28773 , n28607 , n28772 );
or ( n28774 , n28606 , n28773 );
and ( n28775 , n28603 , n28774 );
or ( n28776 , n28602 , n28775 );
and ( n28777 , n28599 , n28776 );
or ( n28778 , n28598 , n28777 );
and ( n28779 , n28595 , n28778 );
or ( n28780 , n28594 , n28779 );
and ( n28781 , n28591 , n28780 );
or ( n28782 , n28590 , n28781 );
and ( n28783 , n28587 , n28782 );
or ( n28784 , n28586 , n28783 );
and ( n28785 , n28583 , n28784 );
or ( n28786 , n28582 , n28785 );
and ( n28787 , n28579 , n28786 );
or ( n28788 , n28578 , n28787 );
and ( n28789 , n28575 , n28788 );
or ( n28790 , n28574 , n28789 );
and ( n28791 , n28571 , n28790 );
or ( n28792 , n28570 , n28791 );
and ( n28793 , n28567 , n28792 );
or ( n28794 , n28566 , n28793 );
and ( n28795 , n28563 , n28794 );
or ( n28796 , n28562 , n28795 );
and ( n28797 , n28559 , n28796 );
or ( n28798 , n28558 , n28797 );
and ( n28799 , n28555 , n28798 );
or ( n28800 , n28554 , n28799 );
and ( n28801 , n28551 , n28800 );
or ( n28802 , n28550 , n28801 );
and ( n28803 , n28547 , n28802 );
or ( n28804 , n28546 , n28803 );
and ( n28805 , n28543 , n28804 );
or ( n28806 , n28542 , n28805 );
and ( n28807 , n28539 , n28806 );
or ( n28808 , n28538 , n28807 );
and ( n28809 , n28535 , n28808 );
or ( n28810 , n28534 , n28809 );
and ( n28811 , n28531 , n28810 );
or ( n28812 , n28530 , n28811 );
and ( n28813 , n28527 , n28812 );
or ( n28814 , n28526 , n28813 );
and ( n28815 , n28523 , n28814 );
or ( n28816 , n28522 , n28815 );
and ( n28817 , n28519 , n28816 );
or ( n28818 , n28518 , n28817 );
and ( n28819 , n28515 , n28818 );
or ( n28820 , n28514 , n28819 );
and ( n28821 , n28511 , n28820 );
or ( n28822 , n28510 , n28821 );
and ( n28823 , n28507 , n28822 );
or ( n28824 , n28506 , n28823 );
and ( n28825 , n28503 , n28824 );
or ( n28826 , n28502 , n28825 );
and ( n28827 , n28499 , n28826 );
or ( n28828 , n28498 , n28827 );
and ( n28829 , n28495 , n28828 );
or ( n28830 , n28494 , n28829 );
xor ( n28831 , n28491 , n28830 );
buf ( n28832 , n475 );
not ( n28833 , n28832 );
nor ( n28834 , n601 , n28833 );
buf ( n28835 , n28834 );
nor ( n28836 , n622 , n26660 );
xor ( n28837 , n28835 , n28836 );
buf ( n28838 , n28837 );
nor ( n28839 , n646 , n25600 );
xor ( n28840 , n28838 , n28839 );
and ( n28841 , n27739 , n27740 );
buf ( n28842 , n28841 );
xor ( n28843 , n28840 , n28842 );
nor ( n28844 , n684 , n24564 );
xor ( n28845 , n28843 , n28844 );
and ( n28846 , n27742 , n27743 );
and ( n28847 , n27744 , n27746 );
or ( n28848 , n28846 , n28847 );
xor ( n28849 , n28845 , n28848 );
nor ( n28850 , n733 , n23541 );
xor ( n28851 , n28849 , n28850 );
and ( n28852 , n27747 , n27748 );
and ( n28853 , n27749 , n27752 );
or ( n28854 , n28852 , n28853 );
xor ( n28855 , n28851 , n28854 );
nor ( n28856 , n796 , n22541 );
xor ( n28857 , n28855 , n28856 );
and ( n28858 , n27753 , n27754 );
and ( n28859 , n27755 , n27758 );
or ( n28860 , n28858 , n28859 );
xor ( n28861 , n28857 , n28860 );
nor ( n28862 , n868 , n21562 );
xor ( n28863 , n28861 , n28862 );
and ( n28864 , n27759 , n27760 );
and ( n28865 , n27761 , n27764 );
or ( n28866 , n28864 , n28865 );
xor ( n28867 , n28863 , n28866 );
nor ( n28868 , n958 , n20601 );
xor ( n28869 , n28867 , n28868 );
and ( n28870 , n27765 , n27766 );
and ( n28871 , n27767 , n27770 );
or ( n28872 , n28870 , n28871 );
xor ( n28873 , n28869 , n28872 );
nor ( n28874 , n1062 , n19657 );
xor ( n28875 , n28873 , n28874 );
and ( n28876 , n27771 , n27772 );
and ( n28877 , n27773 , n27776 );
or ( n28878 , n28876 , n28877 );
xor ( n28879 , n28875 , n28878 );
nor ( n28880 , n1176 , n18734 );
xor ( n28881 , n28879 , n28880 );
and ( n28882 , n27777 , n27778 );
and ( n28883 , n27779 , n27782 );
or ( n28884 , n28882 , n28883 );
xor ( n28885 , n28881 , n28884 );
nor ( n28886 , n1303 , n17828 );
xor ( n28887 , n28885 , n28886 );
and ( n28888 , n27783 , n27784 );
and ( n28889 , n27785 , n27788 );
or ( n28890 , n28888 , n28889 );
xor ( n28891 , n28887 , n28890 );
nor ( n28892 , n1445 , n16943 );
xor ( n28893 , n28891 , n28892 );
and ( n28894 , n27789 , n27790 );
and ( n28895 , n27791 , n27794 );
or ( n28896 , n28894 , n28895 );
xor ( n28897 , n28893 , n28896 );
nor ( n28898 , n1598 , n16077 );
xor ( n28899 , n28897 , n28898 );
and ( n28900 , n27795 , n27796 );
and ( n28901 , n27797 , n27800 );
or ( n28902 , n28900 , n28901 );
xor ( n28903 , n28899 , n28902 );
nor ( n28904 , n1766 , n15230 );
xor ( n28905 , n28903 , n28904 );
and ( n28906 , n27801 , n27802 );
and ( n28907 , n27803 , n27806 );
or ( n28908 , n28906 , n28907 );
xor ( n28909 , n28905 , n28908 );
nor ( n28910 , n1945 , n14403 );
xor ( n28911 , n28909 , n28910 );
and ( n28912 , n27807 , n27808 );
and ( n28913 , n27809 , n27812 );
or ( n28914 , n28912 , n28913 );
xor ( n28915 , n28911 , n28914 );
nor ( n28916 , n2137 , n13599 );
xor ( n28917 , n28915 , n28916 );
and ( n28918 , n27813 , n27814 );
and ( n28919 , n27815 , n27818 );
or ( n28920 , n28918 , n28919 );
xor ( n28921 , n28917 , n28920 );
nor ( n28922 , n2343 , n12808 );
xor ( n28923 , n28921 , n28922 );
and ( n28924 , n27819 , n27820 );
and ( n28925 , n27821 , n27824 );
or ( n28926 , n28924 , n28925 );
xor ( n28927 , n28923 , n28926 );
nor ( n28928 , n2566 , n12037 );
xor ( n28929 , n28927 , n28928 );
and ( n28930 , n27825 , n27826 );
and ( n28931 , n27827 , n27830 );
or ( n28932 , n28930 , n28931 );
xor ( n28933 , n28929 , n28932 );
nor ( n28934 , n2797 , n11282 );
xor ( n28935 , n28933 , n28934 );
and ( n28936 , n27831 , n27832 );
and ( n28937 , n27833 , n27836 );
or ( n28938 , n28936 , n28937 );
xor ( n28939 , n28935 , n28938 );
nor ( n28940 , n3043 , n10547 );
xor ( n28941 , n28939 , n28940 );
and ( n28942 , n27837 , n27838 );
and ( n28943 , n27839 , n27842 );
or ( n28944 , n28942 , n28943 );
xor ( n28945 , n28941 , n28944 );
nor ( n28946 , n3300 , n9829 );
xor ( n28947 , n28945 , n28946 );
and ( n28948 , n27843 , n27844 );
and ( n28949 , n27845 , n27848 );
or ( n28950 , n28948 , n28949 );
xor ( n28951 , n28947 , n28950 );
nor ( n28952 , n3570 , n8955 );
xor ( n28953 , n28951 , n28952 );
and ( n28954 , n27849 , n27850 );
and ( n28955 , n27851 , n27854 );
or ( n28956 , n28954 , n28955 );
xor ( n28957 , n28953 , n28956 );
nor ( n28958 , n3853 , n603 );
xor ( n28959 , n28957 , n28958 );
and ( n28960 , n27855 , n27856 );
and ( n28961 , n27857 , n27860 );
or ( n28962 , n28960 , n28961 );
xor ( n28963 , n28959 , n28962 );
nor ( n28964 , n4151 , n652 );
xor ( n28965 , n28963 , n28964 );
and ( n28966 , n27861 , n27862 );
and ( n28967 , n27863 , n27866 );
or ( n28968 , n28966 , n28967 );
xor ( n28969 , n28965 , n28968 );
nor ( n28970 , n4458 , n624 );
xor ( n28971 , n28969 , n28970 );
and ( n28972 , n27867 , n27868 );
and ( n28973 , n27869 , n27872 );
or ( n28974 , n28972 , n28973 );
xor ( n28975 , n28971 , n28974 );
nor ( n28976 , n4786 , n648 );
xor ( n28977 , n28975 , n28976 );
and ( n28978 , n27873 , n27874 );
and ( n28979 , n27875 , n27878 );
or ( n28980 , n28978 , n28979 );
xor ( n28981 , n28977 , n28980 );
nor ( n28982 , n5126 , n686 );
xor ( n28983 , n28981 , n28982 );
and ( n28984 , n27879 , n27880 );
and ( n28985 , n27881 , n27884 );
or ( n28986 , n28984 , n28985 );
xor ( n28987 , n28983 , n28986 );
nor ( n28988 , n5477 , n735 );
xor ( n28989 , n28987 , n28988 );
and ( n28990 , n27885 , n27886 );
and ( n28991 , n27887 , n27890 );
or ( n28992 , n28990 , n28991 );
xor ( n28993 , n28989 , n28992 );
nor ( n28994 , n5838 , n798 );
xor ( n28995 , n28993 , n28994 );
and ( n28996 , n27891 , n27892 );
and ( n28997 , n27893 , n27896 );
or ( n28998 , n28996 , n28997 );
xor ( n28999 , n28995 , n28998 );
nor ( n29000 , n6212 , n870 );
xor ( n29001 , n28999 , n29000 );
and ( n29002 , n27897 , n27898 );
and ( n29003 , n27899 , n27902 );
or ( n29004 , n29002 , n29003 );
xor ( n29005 , n29001 , n29004 );
nor ( n29006 , n6596 , n960 );
xor ( n29007 , n29005 , n29006 );
and ( n29008 , n27903 , n27904 );
and ( n29009 , n27905 , n27908 );
or ( n29010 , n29008 , n29009 );
xor ( n29011 , n29007 , n29010 );
nor ( n29012 , n6997 , n1064 );
xor ( n29013 , n29011 , n29012 );
and ( n29014 , n27909 , n27910 );
and ( n29015 , n27911 , n27914 );
or ( n29016 , n29014 , n29015 );
xor ( n29017 , n29013 , n29016 );
nor ( n29018 , n7413 , n1178 );
xor ( n29019 , n29017 , n29018 );
and ( n29020 , n27915 , n27916 );
and ( n29021 , n27917 , n27920 );
or ( n29022 , n29020 , n29021 );
xor ( n29023 , n29019 , n29022 );
nor ( n29024 , n7841 , n1305 );
xor ( n29025 , n29023 , n29024 );
and ( n29026 , n27921 , n27922 );
and ( n29027 , n27923 , n27926 );
or ( n29028 , n29026 , n29027 );
xor ( n29029 , n29025 , n29028 );
nor ( n29030 , n8281 , n1447 );
xor ( n29031 , n29029 , n29030 );
and ( n29032 , n27927 , n27928 );
and ( n29033 , n27929 , n27932 );
or ( n29034 , n29032 , n29033 );
xor ( n29035 , n29031 , n29034 );
nor ( n29036 , n8737 , n1600 );
xor ( n29037 , n29035 , n29036 );
and ( n29038 , n27933 , n27934 );
and ( n29039 , n27935 , n27938 );
or ( n29040 , n29038 , n29039 );
xor ( n29041 , n29037 , n29040 );
nor ( n29042 , n9420 , n1768 );
xor ( n29043 , n29041 , n29042 );
and ( n29044 , n27939 , n27940 );
and ( n29045 , n27941 , n27944 );
or ( n29046 , n29044 , n29045 );
xor ( n29047 , n29043 , n29046 );
nor ( n29048 , n10312 , n1947 );
xor ( n29049 , n29047 , n29048 );
and ( n29050 , n27945 , n27946 );
and ( n29051 , n27947 , n27950 );
or ( n29052 , n29050 , n29051 );
xor ( n29053 , n29049 , n29052 );
nor ( n29054 , n11041 , n2139 );
xor ( n29055 , n29053 , n29054 );
and ( n29056 , n27951 , n27952 );
and ( n29057 , n27953 , n27956 );
or ( n29058 , n29056 , n29057 );
xor ( n29059 , n29055 , n29058 );
nor ( n29060 , n11790 , n2345 );
xor ( n29061 , n29059 , n29060 );
and ( n29062 , n27957 , n27958 );
and ( n29063 , n27959 , n27962 );
or ( n29064 , n29062 , n29063 );
xor ( n29065 , n29061 , n29064 );
nor ( n29066 , n12555 , n2568 );
xor ( n29067 , n29065 , n29066 );
and ( n29068 , n27963 , n27964 );
and ( n29069 , n27965 , n27968 );
or ( n29070 , n29068 , n29069 );
xor ( n29071 , n29067 , n29070 );
nor ( n29072 , n13340 , n2799 );
xor ( n29073 , n29071 , n29072 );
and ( n29074 , n27969 , n27970 );
and ( n29075 , n27971 , n27974 );
or ( n29076 , n29074 , n29075 );
xor ( n29077 , n29073 , n29076 );
nor ( n29078 , n14138 , n3045 );
xor ( n29079 , n29077 , n29078 );
and ( n29080 , n27975 , n27976 );
and ( n29081 , n27977 , n27980 );
or ( n29082 , n29080 , n29081 );
xor ( n29083 , n29079 , n29082 );
nor ( n29084 , n14959 , n3302 );
xor ( n29085 , n29083 , n29084 );
and ( n29086 , n27981 , n27982 );
and ( n29087 , n27983 , n27986 );
or ( n29088 , n29086 , n29087 );
xor ( n29089 , n29085 , n29088 );
nor ( n29090 , n15800 , n3572 );
xor ( n29091 , n29089 , n29090 );
and ( n29092 , n27987 , n27988 );
and ( n29093 , n27989 , n27992 );
or ( n29094 , n29092 , n29093 );
xor ( n29095 , n29091 , n29094 );
nor ( n29096 , n16660 , n3855 );
xor ( n29097 , n29095 , n29096 );
and ( n29098 , n27993 , n27994 );
and ( n29099 , n27995 , n27998 );
or ( n29100 , n29098 , n29099 );
xor ( n29101 , n29097 , n29100 );
nor ( n29102 , n17539 , n4153 );
xor ( n29103 , n29101 , n29102 );
and ( n29104 , n27999 , n28000 );
and ( n29105 , n28001 , n28004 );
or ( n29106 , n29104 , n29105 );
xor ( n29107 , n29103 , n29106 );
nor ( n29108 , n18439 , n4460 );
xor ( n29109 , n29107 , n29108 );
and ( n29110 , n28005 , n28006 );
and ( n29111 , n28007 , n28010 );
or ( n29112 , n29110 , n29111 );
xor ( n29113 , n29109 , n29112 );
nor ( n29114 , n19356 , n4788 );
xor ( n29115 , n29113 , n29114 );
and ( n29116 , n28011 , n28012 );
and ( n29117 , n28013 , n28016 );
or ( n29118 , n29116 , n29117 );
xor ( n29119 , n29115 , n29118 );
nor ( n29120 , n20294 , n5128 );
xor ( n29121 , n29119 , n29120 );
and ( n29122 , n28017 , n28018 );
and ( n29123 , n28019 , n28022 );
or ( n29124 , n29122 , n29123 );
xor ( n29125 , n29121 , n29124 );
nor ( n29126 , n21249 , n5479 );
xor ( n29127 , n29125 , n29126 );
and ( n29128 , n28023 , n28024 );
and ( n29129 , n28025 , n28028 );
or ( n29130 , n29128 , n29129 );
xor ( n29131 , n29127 , n29130 );
nor ( n29132 , n22222 , n5840 );
xor ( n29133 , n29131 , n29132 );
and ( n29134 , n28029 , n28030 );
and ( n29135 , n28031 , n28034 );
or ( n29136 , n29134 , n29135 );
xor ( n29137 , n29133 , n29136 );
nor ( n29138 , n23216 , n6214 );
xor ( n29139 , n29137 , n29138 );
and ( n29140 , n28035 , n28036 );
and ( n29141 , n28037 , n28040 );
or ( n29142 , n29140 , n29141 );
xor ( n29143 , n29139 , n29142 );
nor ( n29144 , n24233 , n6598 );
xor ( n29145 , n29143 , n29144 );
and ( n29146 , n28041 , n28042 );
and ( n29147 , n28043 , n28046 );
or ( n29148 , n29146 , n29147 );
xor ( n29149 , n29145 , n29148 );
nor ( n29150 , n25263 , n6999 );
xor ( n29151 , n29149 , n29150 );
and ( n29152 , n28047 , n28048 );
and ( n29153 , n28049 , n28052 );
or ( n29154 , n29152 , n29153 );
xor ( n29155 , n29151 , n29154 );
nor ( n29156 , n26317 , n7415 );
xor ( n29157 , n29155 , n29156 );
and ( n29158 , n28053 , n28054 );
and ( n29159 , n28055 , n28058 );
or ( n29160 , n29158 , n29159 );
xor ( n29161 , n29157 , n29160 );
nor ( n29162 , n27388 , n7843 );
xor ( n29163 , n29161 , n29162 );
and ( n29164 , n28059 , n28060 );
and ( n29165 , n28061 , n28064 );
or ( n29166 , n29164 , n29165 );
xor ( n29167 , n29163 , n29166 );
nor ( n29168 , n28478 , n8283 );
xor ( n29169 , n29167 , n29168 );
and ( n29170 , n28065 , n28066 );
and ( n29171 , n28067 , n28070 );
or ( n29172 , n29170 , n29171 );
xor ( n29173 , n29169 , n29172 );
and ( n29174 , n28422 , n28423 );
and ( n29175 , n28423 , n28463 );
and ( n29176 , n28422 , n28463 );
or ( n29177 , n29174 , n29175 , n29176 );
and ( n29178 , n28084 , n28417 );
and ( n29179 , n28417 , n28464 );
and ( n29180 , n28084 , n28464 );
or ( n29181 , n29178 , n29179 , n29180 );
xor ( n29182 , n29177 , n29181 );
and ( n29183 , n28088 , n28208 );
and ( n29184 , n28208 , n28416 );
and ( n29185 , n28088 , n28416 );
or ( n29186 , n29183 , n29184 , n29185 );
and ( n29187 , n28213 , n28291 );
and ( n29188 , n28291 , n28415 );
and ( n29189 , n28213 , n28415 );
or ( n29190 , n29187 , n29188 , n29189 );
and ( n29191 , n28101 , n28169 );
and ( n29192 , n28169 , n28206 );
and ( n29193 , n28101 , n28206 );
or ( n29194 , n29191 , n29192 , n29193 );
and ( n29195 , n28217 , n28221 );
and ( n29196 , n28221 , n28290 );
and ( n29197 , n28217 , n28290 );
or ( n29198 , n29195 , n29196 , n29197 );
xor ( n29199 , n29194 , n29198 );
and ( n29200 , n28174 , n28178 );
and ( n29201 , n28178 , n28205 );
and ( n29202 , n28174 , n28205 );
or ( n29203 , n29200 , n29201 , n29202 );
and ( n29204 , n28135 , n28151 );
and ( n29205 , n28151 , n28167 );
and ( n29206 , n28135 , n28167 );
or ( n29207 , n29204 , n29205 , n29206 );
and ( n29208 , n28118 , n28122 );
and ( n29209 , n28122 , n28128 );
and ( n29210 , n28118 , n28128 );
or ( n29211 , n29208 , n29209 , n29210 );
and ( n29212 , n28139 , n28144 );
and ( n29213 , n28144 , n28150 );
and ( n29214 , n28139 , n28150 );
or ( n29215 , n29212 , n29213 , n29214 );
xor ( n29216 , n29211 , n29215 );
and ( n29217 , n28124 , n28125 );
and ( n29218 , n28125 , n28127 );
and ( n29219 , n28124 , n28127 );
or ( n29220 , n29217 , n29218 , n29219 );
and ( n29221 , n28140 , n28141 );
and ( n29222 , n28141 , n28143 );
and ( n29223 , n28140 , n28143 );
or ( n29224 , n29221 , n29222 , n29223 );
xor ( n29225 , n29220 , n29224 );
and ( n29226 , n21216 , n940 );
and ( n29227 , n22186 , n840 );
xor ( n29228 , n29226 , n29227 );
and ( n29229 , n22892 , n771 );
xor ( n29230 , n29228 , n29229 );
xor ( n29231 , n29225 , n29230 );
xor ( n29232 , n29216 , n29231 );
xor ( n29233 , n29207 , n29232 );
and ( n29234 , n28156 , n28160 );
and ( n29235 , n28160 , n28166 );
and ( n29236 , n28156 , n28166 );
or ( n29237 , n29234 , n29235 , n29236 );
and ( n29238 , n28146 , n28147 );
and ( n29239 , n28147 , n28149 );
and ( n29240 , n28146 , n28149 );
or ( n29241 , n29238 , n29239 , n29240 );
and ( n29242 , n18144 , n1254 );
and ( n29243 , n19324 , n1134 );
xor ( n29244 , n29242 , n29243 );
and ( n29245 , n20233 , n1034 );
xor ( n29246 , n29244 , n29245 );
xor ( n29247 , n29241 , n29246 );
and ( n29248 , n15758 , n1738 );
and ( n29249 , n16637 , n1551 );
xor ( n29250 , n29248 , n29249 );
and ( n29251 , n17512 , n1424 );
xor ( n29252 , n29250 , n29251 );
xor ( n29253 , n29247 , n29252 );
xor ( n29254 , n29237 , n29253 );
and ( n29255 , n28162 , n28163 );
and ( n29256 , n28163 , n28165 );
and ( n29257 , n28162 , n28165 );
or ( n29258 , n29255 , n29256 , n29257 );
and ( n29259 , n28193 , n28194 );
and ( n29260 , n28194 , n28196 );
and ( n29261 , n28193 , n28196 );
or ( n29262 , n29259 , n29260 , n29261 );
xor ( n29263 , n29258 , n29262 );
and ( n29264 , n13322 , n2298 );
and ( n29265 , n14118 , n2100 );
xor ( n29266 , n29264 , n29265 );
and ( n29267 , n14938 , n1882 );
xor ( n29268 , n29266 , n29267 );
xor ( n29269 , n29263 , n29268 );
xor ( n29270 , n29254 , n29269 );
xor ( n29271 , n29233 , n29270 );
xor ( n29272 , n29203 , n29271 );
and ( n29273 , n28183 , n28187 );
and ( n29274 , n28187 , n28204 );
and ( n29275 , n28183 , n28204 );
or ( n29276 , n29273 , n29274 , n29275 );
and ( n29277 , n28230 , n28245 );
and ( n29278 , n28245 , n28262 );
and ( n29279 , n28230 , n28262 );
or ( n29280 , n29277 , n29278 , n29279 );
xor ( n29281 , n29276 , n29280 );
and ( n29282 , n28192 , n28197 );
and ( n29283 , n28197 , n28203 );
and ( n29284 , n28192 , n28203 );
or ( n29285 , n29282 , n29283 , n29284 );
and ( n29286 , n28234 , n28238 );
and ( n29287 , n28238 , n28244 );
and ( n29288 , n28234 , n28244 );
or ( n29289 , n29286 , n29287 , n29288 );
xor ( n29290 , n29285 , n29289 );
and ( n29291 , n28199 , n28200 );
and ( n29292 , n28200 , n28202 );
and ( n29293 , n28199 , n28202 );
or ( n29294 , n29291 , n29292 , n29293 );
and ( n29295 , n11015 , n2981 );
and ( n29296 , n11769 , n2739 );
xor ( n29297 , n29295 , n29296 );
and ( n29298 , n12320 , n2544 );
xor ( n29299 , n29297 , n29298 );
xor ( n29300 , n29294 , n29299 );
and ( n29301 , n8718 , n3749 );
and ( n29302 , n9400 , n3495 );
xor ( n29303 , n29301 , n29302 );
and ( n29304 , n10291 , n3271 );
xor ( n29305 , n29303 , n29304 );
xor ( n29306 , n29300 , n29305 );
xor ( n29307 , n29290 , n29306 );
xor ( n29308 , n29281 , n29307 );
xor ( n29309 , n29272 , n29308 );
xor ( n29310 , n29199 , n29309 );
xor ( n29311 , n29190 , n29310 );
and ( n29312 , n28296 , n28343 );
and ( n29313 , n28343 , n28414 );
and ( n29314 , n28296 , n28414 );
or ( n29315 , n29312 , n29313 , n29314 );
and ( n29316 , n28226 , n28263 );
and ( n29317 , n28263 , n28289 );
and ( n29318 , n28226 , n28289 );
or ( n29319 , n29316 , n29317 , n29318 );
and ( n29320 , n28300 , n28304 );
and ( n29321 , n28304 , n28342 );
and ( n29322 , n28300 , n28342 );
or ( n29323 , n29320 , n29321 , n29322 );
xor ( n29324 , n29319 , n29323 );
and ( n29325 , n28268 , n28272 );
and ( n29326 , n28272 , n28288 );
and ( n29327 , n28268 , n28288 );
or ( n29328 , n29325 , n29326 , n29327 );
and ( n29329 , n28250 , n28255 );
and ( n29330 , n28255 , n28261 );
and ( n29331 , n28250 , n28261 );
or ( n29332 , n29329 , n29330 , n29331 );
and ( n29333 , n28240 , n28241 );
and ( n29334 , n28241 , n28243 );
and ( n29335 , n28240 , n28243 );
or ( n29336 , n29333 , n29334 , n29335 );
and ( n29337 , n28251 , n28252 );
and ( n29338 , n28252 , n28254 );
and ( n29339 , n28251 , n28254 );
or ( n29340 , n29337 , n29338 , n29339 );
xor ( n29341 , n29336 , n29340 );
and ( n29342 , n7385 , n4730 );
and ( n29343 , n7808 , n4403 );
xor ( n29344 , n29342 , n29343 );
and ( n29345 , n8079 , n4102 );
xor ( n29346 , n29344 , n29345 );
xor ( n29347 , n29341 , n29346 );
xor ( n29348 , n29332 , n29347 );
and ( n29349 , n28257 , n28258 );
and ( n29350 , n28258 , n28260 );
and ( n29351 , n28257 , n28260 );
or ( n29352 , n29349 , n29350 , n29351 );
and ( n29353 , n6187 , n5765 );
and ( n29354 , n6569 , n5408 );
xor ( n29355 , n29353 , n29354 );
and ( n29356 , n6816 , n5103 );
xor ( n29357 , n29355 , n29356 );
xor ( n29358 , n29352 , n29357 );
and ( n29359 , n4959 , n6971 );
and ( n29360 , n5459 , n6504 );
xor ( n29361 , n29359 , n29360 );
and ( n29362 , n5819 , n6132 );
xor ( n29363 , n29361 , n29362 );
xor ( n29364 , n29358 , n29363 );
xor ( n29365 , n29348 , n29364 );
xor ( n29366 , n29328 , n29365 );
and ( n29367 , n28277 , n28281 );
and ( n29368 , n28281 , n28287 );
and ( n29369 , n28277 , n28287 );
or ( n29370 , n29367 , n29368 , n29369 );
and ( n29371 , n28313 , n28318 );
and ( n29372 , n28318 , n28324 );
and ( n29373 , n28313 , n28324 );
or ( n29374 , n29371 , n29372 , n29373 );
xor ( n29375 , n29370 , n29374 );
and ( n29376 , n28283 , n28284 );
and ( n29377 , n28284 , n28286 );
and ( n29378 , n28283 , n28286 );
or ( n29379 , n29376 , n29377 , n29378 );
and ( n29380 , n28314 , n28315 );
and ( n29381 , n28315 , n28317 );
and ( n29382 , n28314 , n28317 );
or ( n29383 , n29380 , n29381 , n29382 );
xor ( n29384 , n29379 , n29383 );
and ( n29385 , n4132 , n8243 );
and ( n29386 , n4438 , n7662 );
xor ( n29387 , n29385 , n29386 );
and ( n29388 , n4766 , n7310 );
xor ( n29389 , n29387 , n29388 );
xor ( n29390 , n29384 , n29389 );
xor ( n29391 , n29375 , n29390 );
xor ( n29392 , n29366 , n29391 );
xor ( n29393 , n29324 , n29392 );
xor ( n29394 , n29315 , n29393 );
and ( n29395 , n28348 , n28374 );
and ( n29396 , n28374 , n28413 );
and ( n29397 , n28348 , n28413 );
or ( n29398 , n29395 , n29396 , n29397 );
and ( n29399 , n28309 , n28325 );
and ( n29400 , n28325 , n28341 );
and ( n29401 , n28309 , n28341 );
or ( n29402 , n29399 , n29400 , n29401 );
and ( n29403 , n28352 , n28356 );
and ( n29404 , n28356 , n28373 );
and ( n29405 , n28352 , n28373 );
or ( n29406 , n29403 , n29404 , n29405 );
xor ( n29407 , n29402 , n29406 );
and ( n29408 , n28330 , n28334 );
and ( n29409 , n28334 , n28340 );
and ( n29410 , n28330 , n28340 );
or ( n29411 , n29408 , n29409 , n29410 );
and ( n29412 , n28320 , n28321 );
and ( n29413 , n28321 , n28323 );
and ( n29414 , n28320 , n28323 );
or ( n29415 , n29412 , n29413 , n29414 );
and ( n29416 , n3182 , n10239 );
and ( n29417 , n3545 , n9348 );
xor ( n29418 , n29416 , n29417 );
and ( n29419 , n3801 , n8669 );
xor ( n29420 , n29418 , n29419 );
xor ( n29421 , n29415 , n29420 );
and ( n29422 , n2462 , n12531 );
and ( n29423 , n2779 , n11718 );
xor ( n29424 , n29422 , n29423 );
and ( n29425 , n3024 , n10977 );
xor ( n29426 , n29424 , n29425 );
xor ( n29427 , n29421 , n29426 );
xor ( n29428 , n29411 , n29427 );
and ( n29429 , n28336 , n28337 );
and ( n29430 , n28337 , n28339 );
and ( n29431 , n28336 , n28339 );
or ( n29432 , n29429 , n29430 , n29431 );
and ( n29433 , n28362 , n28363 );
and ( n29434 , n28363 , n28365 );
and ( n29435 , n28362 , n28365 );
or ( n29436 , n29433 , n29434 , n29435 );
xor ( n29437 , n29432 , n29436 );
and ( n29438 , n1933 , n14838 );
and ( n29439 , n2120 , n14044 );
xor ( n29440 , n29438 , n29439 );
and ( n29441 , n2324 , n13256 );
xor ( n29442 , n29440 , n29441 );
xor ( n29443 , n29437 , n29442 );
xor ( n29444 , n29428 , n29443 );
xor ( n29445 , n29407 , n29444 );
xor ( n29446 , n29398 , n29445 );
and ( n29447 , n28379 , n28394 );
and ( n29448 , n28394 , n28412 );
and ( n29449 , n28379 , n28412 );
or ( n29450 , n29447 , n29448 , n29449 );
and ( n29451 , n28361 , n28366 );
and ( n29452 , n28366 , n28372 );
and ( n29453 , n28361 , n28372 );
or ( n29454 , n29451 , n29452 , n29453 );
and ( n29455 , n28383 , n28387 );
and ( n29456 , n28387 , n28393 );
and ( n29457 , n28383 , n28393 );
or ( n29458 , n29455 , n29456 , n29457 );
xor ( n29459 , n29454 , n29458 );
and ( n29460 , n28368 , n28369 );
and ( n29461 , n28369 , n28371 );
and ( n29462 , n28368 , n28371 );
or ( n29463 , n29460 , n29461 , n29462 );
and ( n29464 , n1383 , n17422 );
and ( n29465 , n1580 , n16550 );
xor ( n29466 , n29464 , n29465 );
and ( n29467 , n1694 , n15691 );
xor ( n29468 , n29466 , n29467 );
xor ( n29469 , n29463 , n29468 );
and ( n29470 , n1047 , n20156 );
and ( n29471 , n1164 , n19222 );
xor ( n29472 , n29470 , n29471 );
and ( n29473 , n1287 , n18407 );
xor ( n29474 , n29472 , n29473 );
xor ( n29475 , n29469 , n29474 );
xor ( n29476 , n29459 , n29475 );
xor ( n29477 , n29450 , n29476 );
and ( n29478 , n28399 , n28404 );
and ( n29479 , n28404 , n28411 );
and ( n29480 , n28399 , n28411 );
or ( n29481 , n29478 , n29479 , n29480 );
and ( n29482 , n28389 , n28390 );
and ( n29483 , n28390 , n28392 );
and ( n29484 , n28389 , n28392 );
or ( n29485 , n29482 , n29483 , n29484 );
and ( n29486 , n28400 , n28401 );
and ( n29487 , n28401 , n28403 );
and ( n29488 , n28400 , n28403 );
or ( n29489 , n29486 , n29487 , n29488 );
xor ( n29490 , n29485 , n29489 );
and ( n29491 , n783 , n23075 );
and ( n29492 , n856 , n22065 );
xor ( n29493 , n29491 , n29492 );
and ( n29494 , n925 , n20976 );
xor ( n29495 , n29493 , n29494 );
xor ( n29496 , n29490 , n29495 );
xor ( n29497 , n29481 , n29496 );
and ( n29498 , n28407 , n28408 );
and ( n29499 , n28408 , n28410 );
and ( n29500 , n28407 , n28410 );
or ( n29501 , n29498 , n29499 , n29500 );
and ( n29502 , n632 , n26216 );
and ( n29503 , n671 , n25163 );
xor ( n29504 , n29502 , n29503 );
and ( n29505 , n715 , n24137 );
xor ( n29506 , n29504 , n29505 );
xor ( n29507 , n29501 , n29506 );
buf ( n29508 , n411 );
and ( n29509 , n599 , n29508 );
and ( n29510 , n608 , n28406 );
xor ( n29511 , n29509 , n29510 );
and ( n29512 , n611 , n27296 );
xor ( n29513 , n29511 , n29512 );
xor ( n29514 , n29507 , n29513 );
xor ( n29515 , n29497 , n29514 );
xor ( n29516 , n29477 , n29515 );
xor ( n29517 , n29446 , n29516 );
xor ( n29518 , n29394 , n29517 );
xor ( n29519 , n29311 , n29518 );
xor ( n29520 , n29186 , n29519 );
and ( n29521 , n28092 , n28096 );
and ( n29522 , n28096 , n28207 );
and ( n29523 , n28092 , n28207 );
or ( n29524 , n29521 , n29522 , n29523 );
and ( n29525 , n28428 , n28462 );
xor ( n29526 , n29524 , n29525 );
and ( n29527 , n28432 , n28433 );
and ( n29528 , n28433 , n28461 );
and ( n29529 , n28432 , n28461 );
or ( n29530 , n29527 , n29528 , n29529 );
and ( n29531 , n28105 , n28130 );
and ( n29532 , n28130 , n28168 );
and ( n29533 , n28105 , n28168 );
or ( n29534 , n29531 , n29532 , n29533 );
and ( n29535 , n28438 , n28439 );
and ( n29536 , n28439 , n28460 );
and ( n29537 , n28438 , n28460 );
or ( n29538 , n29535 , n29536 , n29537 );
xor ( n29539 , n29534 , n29538 );
and ( n29540 , n28109 , n28113 );
and ( n29541 , n28113 , n28129 );
and ( n29542 , n28109 , n28129 );
or ( n29543 , n29540 , n29541 , n29542 );
and ( n29544 , n28444 , n28459 );
xor ( n29545 , n29543 , n29544 );
and ( n29546 , n28455 , n28457 );
and ( n29547 , n28448 , n28453 );
and ( n29548 , n28453 , n28458 );
and ( n29549 , n28448 , n28458 );
or ( n29550 , n29547 , n29548 , n29549 );
xor ( n29551 , n29546 , n29550 );
and ( n29552 , n28449 , n28450 );
and ( n29553 , n28450 , n28452 );
and ( n29554 , n28449 , n28452 );
or ( n29555 , n29552 , n29553 , n29554 );
and ( n29556 , n27361 , n606 );
and ( n29557 , n28456 , n615 );
xor ( n29558 , n29556 , n29557 );
buf ( n29559 , n411 );
and ( n29560 , n29559 , n612 );
xor ( n29561 , n29558 , n29560 );
xor ( n29562 , n29555 , n29561 );
and ( n29563 , n24214 , n719 );
and ( n29564 , n25243 , n663 );
xor ( n29565 , n29563 , n29564 );
and ( n29566 , n26296 , n635 );
xor ( n29567 , n29565 , n29566 );
xor ( n29568 , n29562 , n29567 );
xor ( n29569 , n29551 , n29568 );
xor ( n29570 , n29545 , n29569 );
xor ( n29571 , n29539 , n29570 );
xor ( n29572 , n29530 , n29571 );
xor ( n29573 , n29526 , n29572 );
xor ( n29574 , n29520 , n29573 );
xor ( n29575 , n29182 , n29574 );
and ( n29576 , n28075 , n28079 );
and ( n29577 , n28079 , n28465 );
and ( n29578 , n28075 , n28465 );
or ( n29579 , n29576 , n29577 , n29578 );
xor ( n29580 , n29575 , n29579 );
and ( n29581 , n28466 , n28470 );
and ( n29582 , n28471 , n28474 );
or ( n29583 , n29581 , n29582 );
xor ( n29584 , n29580 , n29583 );
buf ( n29585 , n29584 );
buf ( n29586 , n29585 );
not ( n29587 , n29586 );
nor ( n29588 , n29587 , n8739 );
xor ( n29589 , n29173 , n29588 );
and ( n29590 , n28071 , n28479 );
and ( n29591 , n28480 , n28483 );
or ( n29592 , n29590 , n29591 );
xor ( n29593 , n29589 , n29592 );
buf ( n29594 , n29593 );
buf ( n29595 , n29594 );
not ( n29596 , n29595 );
buf ( n29597 , n558 );
not ( n29598 , n29597 );
nor ( n29599 , n29596 , n29598 );
xor ( n29600 , n28831 , n29599 );
xor ( n29601 , n28495 , n28828 );
nor ( n29602 , n28487 , n29598 );
and ( n29603 , n29601 , n29602 );
xor ( n29604 , n29601 , n29602 );
xor ( n29605 , n28499 , n28826 );
nor ( n29606 , n27397 , n29598 );
and ( n29607 , n29605 , n29606 );
xor ( n29608 , n29605 , n29606 );
xor ( n29609 , n28503 , n28824 );
nor ( n29610 , n26326 , n29598 );
and ( n29611 , n29609 , n29610 );
xor ( n29612 , n29609 , n29610 );
xor ( n29613 , n28507 , n28822 );
nor ( n29614 , n25272 , n29598 );
and ( n29615 , n29613 , n29614 );
xor ( n29616 , n29613 , n29614 );
xor ( n29617 , n28511 , n28820 );
nor ( n29618 , n24242 , n29598 );
and ( n29619 , n29617 , n29618 );
xor ( n29620 , n29617 , n29618 );
xor ( n29621 , n28515 , n28818 );
nor ( n29622 , n23225 , n29598 );
and ( n29623 , n29621 , n29622 );
xor ( n29624 , n29621 , n29622 );
xor ( n29625 , n28519 , n28816 );
nor ( n29626 , n22231 , n29598 );
and ( n29627 , n29625 , n29626 );
xor ( n29628 , n29625 , n29626 );
xor ( n29629 , n28523 , n28814 );
nor ( n29630 , n21258 , n29598 );
and ( n29631 , n29629 , n29630 );
xor ( n29632 , n29629 , n29630 );
xor ( n29633 , n28527 , n28812 );
nor ( n29634 , n20303 , n29598 );
and ( n29635 , n29633 , n29634 );
xor ( n29636 , n29633 , n29634 );
xor ( n29637 , n28531 , n28810 );
nor ( n29638 , n19365 , n29598 );
and ( n29639 , n29637 , n29638 );
xor ( n29640 , n29637 , n29638 );
xor ( n29641 , n28535 , n28808 );
nor ( n29642 , n18448 , n29598 );
and ( n29643 , n29641 , n29642 );
xor ( n29644 , n29641 , n29642 );
xor ( n29645 , n28539 , n28806 );
nor ( n29646 , n17548 , n29598 );
and ( n29647 , n29645 , n29646 );
xor ( n29648 , n29645 , n29646 );
xor ( n29649 , n28543 , n28804 );
nor ( n29650 , n16669 , n29598 );
and ( n29651 , n29649 , n29650 );
xor ( n29652 , n29649 , n29650 );
xor ( n29653 , n28547 , n28802 );
nor ( n29654 , n15809 , n29598 );
and ( n29655 , n29653 , n29654 );
xor ( n29656 , n29653 , n29654 );
xor ( n29657 , n28551 , n28800 );
nor ( n29658 , n14968 , n29598 );
and ( n29659 , n29657 , n29658 );
xor ( n29660 , n29657 , n29658 );
xor ( n29661 , n28555 , n28798 );
nor ( n29662 , n14147 , n29598 );
and ( n29663 , n29661 , n29662 );
xor ( n29664 , n29661 , n29662 );
xor ( n29665 , n28559 , n28796 );
nor ( n29666 , n13349 , n29598 );
and ( n29667 , n29665 , n29666 );
xor ( n29668 , n29665 , n29666 );
xor ( n29669 , n28563 , n28794 );
nor ( n29670 , n12564 , n29598 );
and ( n29671 , n29669 , n29670 );
xor ( n29672 , n29669 , n29670 );
xor ( n29673 , n28567 , n28792 );
nor ( n29674 , n11799 , n29598 );
and ( n29675 , n29673 , n29674 );
xor ( n29676 , n29673 , n29674 );
xor ( n29677 , n28571 , n28790 );
nor ( n29678 , n11050 , n29598 );
and ( n29679 , n29677 , n29678 );
xor ( n29680 , n29677 , n29678 );
xor ( n29681 , n28575 , n28788 );
nor ( n29682 , n10321 , n29598 );
and ( n29683 , n29681 , n29682 );
xor ( n29684 , n29681 , n29682 );
xor ( n29685 , n28579 , n28786 );
nor ( n29686 , n9429 , n29598 );
and ( n29687 , n29685 , n29686 );
xor ( n29688 , n29685 , n29686 );
xor ( n29689 , n28583 , n28784 );
nor ( n29690 , n8949 , n29598 );
and ( n29691 , n29689 , n29690 );
xor ( n29692 , n29689 , n29690 );
xor ( n29693 , n28587 , n28782 );
nor ( n29694 , n9437 , n29598 );
and ( n29695 , n29693 , n29694 );
xor ( n29696 , n29693 , n29694 );
xor ( n29697 , n28591 , n28780 );
nor ( n29698 , n9446 , n29598 );
and ( n29699 , n29697 , n29698 );
xor ( n29700 , n29697 , n29698 );
xor ( n29701 , n28595 , n28778 );
nor ( n29702 , n9455 , n29598 );
and ( n29703 , n29701 , n29702 );
xor ( n29704 , n29701 , n29702 );
xor ( n29705 , n28599 , n28776 );
nor ( n29706 , n9464 , n29598 );
and ( n29707 , n29705 , n29706 );
xor ( n29708 , n29705 , n29706 );
xor ( n29709 , n28603 , n28774 );
nor ( n29710 , n9473 , n29598 );
and ( n29711 , n29709 , n29710 );
xor ( n29712 , n29709 , n29710 );
xor ( n29713 , n28607 , n28772 );
nor ( n29714 , n9482 , n29598 );
and ( n29715 , n29713 , n29714 );
xor ( n29716 , n29713 , n29714 );
xor ( n29717 , n28611 , n28770 );
nor ( n29718 , n9491 , n29598 );
and ( n29719 , n29717 , n29718 );
xor ( n29720 , n29717 , n29718 );
xor ( n29721 , n28615 , n28768 );
nor ( n29722 , n9500 , n29598 );
and ( n29723 , n29721 , n29722 );
xor ( n29724 , n29721 , n29722 );
xor ( n29725 , n28619 , n28766 );
nor ( n29726 , n9509 , n29598 );
and ( n29727 , n29725 , n29726 );
xor ( n29728 , n29725 , n29726 );
xor ( n29729 , n28623 , n28764 );
nor ( n29730 , n9518 , n29598 );
and ( n29731 , n29729 , n29730 );
xor ( n29732 , n29729 , n29730 );
xor ( n29733 , n28627 , n28762 );
nor ( n29734 , n9527 , n29598 );
and ( n29735 , n29733 , n29734 );
xor ( n29736 , n29733 , n29734 );
xor ( n29737 , n28631 , n28760 );
nor ( n29738 , n9536 , n29598 );
and ( n29739 , n29737 , n29738 );
xor ( n29740 , n29737 , n29738 );
xor ( n29741 , n28635 , n28758 );
nor ( n29742 , n9545 , n29598 );
and ( n29743 , n29741 , n29742 );
xor ( n29744 , n29741 , n29742 );
xor ( n29745 , n28639 , n28756 );
nor ( n29746 , n9554 , n29598 );
and ( n29747 , n29745 , n29746 );
xor ( n29748 , n29745 , n29746 );
xor ( n29749 , n28643 , n28754 );
nor ( n29750 , n9563 , n29598 );
and ( n29751 , n29749 , n29750 );
xor ( n29752 , n29749 , n29750 );
xor ( n29753 , n28647 , n28752 );
nor ( n29754 , n9572 , n29598 );
and ( n29755 , n29753 , n29754 );
xor ( n29756 , n29753 , n29754 );
xor ( n29757 , n28651 , n28750 );
nor ( n29758 , n9581 , n29598 );
and ( n29759 , n29757 , n29758 );
xor ( n29760 , n29757 , n29758 );
xor ( n29761 , n28655 , n28748 );
nor ( n29762 , n9590 , n29598 );
and ( n29763 , n29761 , n29762 );
xor ( n29764 , n29761 , n29762 );
xor ( n29765 , n28659 , n28746 );
nor ( n29766 , n9599 , n29598 );
and ( n29767 , n29765 , n29766 );
xor ( n29768 , n29765 , n29766 );
xor ( n29769 , n28663 , n28744 );
nor ( n29770 , n9608 , n29598 );
and ( n29771 , n29769 , n29770 );
xor ( n29772 , n29769 , n29770 );
xor ( n29773 , n28667 , n28742 );
nor ( n29774 , n9617 , n29598 );
and ( n29775 , n29773 , n29774 );
xor ( n29776 , n29773 , n29774 );
xor ( n29777 , n28671 , n28740 );
nor ( n29778 , n9626 , n29598 );
and ( n29779 , n29777 , n29778 );
xor ( n29780 , n29777 , n29778 );
xor ( n29781 , n28675 , n28738 );
nor ( n29782 , n9635 , n29598 );
and ( n29783 , n29781 , n29782 );
xor ( n29784 , n29781 , n29782 );
xor ( n29785 , n28679 , n28736 );
nor ( n29786 , n9644 , n29598 );
and ( n29787 , n29785 , n29786 );
xor ( n29788 , n29785 , n29786 );
xor ( n29789 , n28683 , n28734 );
nor ( n29790 , n9653 , n29598 );
and ( n29791 , n29789 , n29790 );
xor ( n29792 , n29789 , n29790 );
xor ( n29793 , n28687 , n28732 );
nor ( n29794 , n9662 , n29598 );
and ( n29795 , n29793 , n29794 );
xor ( n29796 , n29793 , n29794 );
xor ( n29797 , n28691 , n28730 );
nor ( n29798 , n9671 , n29598 );
and ( n29799 , n29797 , n29798 );
xor ( n29800 , n29797 , n29798 );
xor ( n29801 , n28695 , n28728 );
nor ( n29802 , n9680 , n29598 );
and ( n29803 , n29801 , n29802 );
xor ( n29804 , n29801 , n29802 );
xor ( n29805 , n28699 , n28726 );
nor ( n29806 , n9689 , n29598 );
and ( n29807 , n29805 , n29806 );
xor ( n29808 , n29805 , n29806 );
xor ( n29809 , n28703 , n28724 );
nor ( n29810 , n9698 , n29598 );
and ( n29811 , n29809 , n29810 );
xor ( n29812 , n29809 , n29810 );
xor ( n29813 , n28707 , n28722 );
nor ( n29814 , n9707 , n29598 );
and ( n29815 , n29813 , n29814 );
xor ( n29816 , n29813 , n29814 );
xor ( n29817 , n28711 , n28720 );
nor ( n29818 , n9716 , n29598 );
and ( n29819 , n29817 , n29818 );
xor ( n29820 , n29817 , n29818 );
xor ( n29821 , n28715 , n28718 );
nor ( n29822 , n9725 , n29598 );
and ( n29823 , n29821 , n29822 );
xor ( n29824 , n29821 , n29822 );
xor ( n29825 , n28716 , n28717 );
nor ( n29826 , n9734 , n29598 );
and ( n29827 , n29825 , n29826 );
xor ( n29828 , n29825 , n29826 );
nor ( n29829 , n9752 , n28489 );
nor ( n29830 , n9743 , n29598 );
and ( n29831 , n29829 , n29830 );
and ( n29832 , n29828 , n29831 );
or ( n29833 , n29827 , n29832 );
and ( n29834 , n29824 , n29833 );
or ( n29835 , n29823 , n29834 );
and ( n29836 , n29820 , n29835 );
or ( n29837 , n29819 , n29836 );
and ( n29838 , n29816 , n29837 );
or ( n29839 , n29815 , n29838 );
and ( n29840 , n29812 , n29839 );
or ( n29841 , n29811 , n29840 );
and ( n29842 , n29808 , n29841 );
or ( n29843 , n29807 , n29842 );
and ( n29844 , n29804 , n29843 );
or ( n29845 , n29803 , n29844 );
and ( n29846 , n29800 , n29845 );
or ( n29847 , n29799 , n29846 );
and ( n29848 , n29796 , n29847 );
or ( n29849 , n29795 , n29848 );
and ( n29850 , n29792 , n29849 );
or ( n29851 , n29791 , n29850 );
and ( n29852 , n29788 , n29851 );
or ( n29853 , n29787 , n29852 );
and ( n29854 , n29784 , n29853 );
or ( n29855 , n29783 , n29854 );
and ( n29856 , n29780 , n29855 );
or ( n29857 , n29779 , n29856 );
and ( n29858 , n29776 , n29857 );
or ( n29859 , n29775 , n29858 );
and ( n29860 , n29772 , n29859 );
or ( n29861 , n29771 , n29860 );
and ( n29862 , n29768 , n29861 );
or ( n29863 , n29767 , n29862 );
and ( n29864 , n29764 , n29863 );
or ( n29865 , n29763 , n29864 );
and ( n29866 , n29760 , n29865 );
or ( n29867 , n29759 , n29866 );
and ( n29868 , n29756 , n29867 );
or ( n29869 , n29755 , n29868 );
and ( n29870 , n29752 , n29869 );
or ( n29871 , n29751 , n29870 );
and ( n29872 , n29748 , n29871 );
or ( n29873 , n29747 , n29872 );
and ( n29874 , n29744 , n29873 );
or ( n29875 , n29743 , n29874 );
and ( n29876 , n29740 , n29875 );
or ( n29877 , n29739 , n29876 );
and ( n29878 , n29736 , n29877 );
or ( n29879 , n29735 , n29878 );
and ( n29880 , n29732 , n29879 );
or ( n29881 , n29731 , n29880 );
and ( n29882 , n29728 , n29881 );
or ( n29883 , n29727 , n29882 );
and ( n29884 , n29724 , n29883 );
or ( n29885 , n29723 , n29884 );
and ( n29886 , n29720 , n29885 );
or ( n29887 , n29719 , n29886 );
and ( n29888 , n29716 , n29887 );
or ( n29889 , n29715 , n29888 );
and ( n29890 , n29712 , n29889 );
or ( n29891 , n29711 , n29890 );
and ( n29892 , n29708 , n29891 );
or ( n29893 , n29707 , n29892 );
and ( n29894 , n29704 , n29893 );
or ( n29895 , n29703 , n29894 );
and ( n29896 , n29700 , n29895 );
or ( n29897 , n29699 , n29896 );
and ( n29898 , n29696 , n29897 );
or ( n29899 , n29695 , n29898 );
and ( n29900 , n29692 , n29899 );
or ( n29901 , n29691 , n29900 );
and ( n29902 , n29688 , n29901 );
or ( n29903 , n29687 , n29902 );
and ( n29904 , n29684 , n29903 );
or ( n29905 , n29683 , n29904 );
and ( n29906 , n29680 , n29905 );
or ( n29907 , n29679 , n29906 );
and ( n29908 , n29676 , n29907 );
or ( n29909 , n29675 , n29908 );
and ( n29910 , n29672 , n29909 );
or ( n29911 , n29671 , n29910 );
and ( n29912 , n29668 , n29911 );
or ( n29913 , n29667 , n29912 );
and ( n29914 , n29664 , n29913 );
or ( n29915 , n29663 , n29914 );
and ( n29916 , n29660 , n29915 );
or ( n29917 , n29659 , n29916 );
and ( n29918 , n29656 , n29917 );
or ( n29919 , n29655 , n29918 );
and ( n29920 , n29652 , n29919 );
or ( n29921 , n29651 , n29920 );
and ( n29922 , n29648 , n29921 );
or ( n29923 , n29647 , n29922 );
and ( n29924 , n29644 , n29923 );
or ( n29925 , n29643 , n29924 );
and ( n29926 , n29640 , n29925 );
or ( n29927 , n29639 , n29926 );
and ( n29928 , n29636 , n29927 );
or ( n29929 , n29635 , n29928 );
and ( n29930 , n29632 , n29929 );
or ( n29931 , n29631 , n29930 );
and ( n29932 , n29628 , n29931 );
or ( n29933 , n29627 , n29932 );
and ( n29934 , n29624 , n29933 );
or ( n29935 , n29623 , n29934 );
and ( n29936 , n29620 , n29935 );
or ( n29937 , n29619 , n29936 );
and ( n29938 , n29616 , n29937 );
or ( n29939 , n29615 , n29938 );
and ( n29940 , n29612 , n29939 );
or ( n29941 , n29611 , n29940 );
and ( n29942 , n29608 , n29941 );
or ( n29943 , n29607 , n29942 );
and ( n29944 , n29604 , n29943 );
or ( n29945 , n29603 , n29944 );
xor ( n29946 , n29600 , n29945 );
buf ( n29947 , n474 );
not ( n29948 , n29947 );
nor ( n29949 , n601 , n29948 );
buf ( n29950 , n29949 );
nor ( n29951 , n622 , n27737 );
xor ( n29952 , n29950 , n29951 );
buf ( n29953 , n29952 );
nor ( n29954 , n646 , n26660 );
xor ( n29955 , n29953 , n29954 );
and ( n29956 , n28835 , n28836 );
buf ( n29957 , n29956 );
xor ( n29958 , n29955 , n29957 );
nor ( n29959 , n684 , n25600 );
xor ( n29960 , n29958 , n29959 );
and ( n29961 , n28838 , n28839 );
and ( n29962 , n28840 , n28842 );
or ( n29963 , n29961 , n29962 );
xor ( n29964 , n29960 , n29963 );
nor ( n29965 , n733 , n24564 );
xor ( n29966 , n29964 , n29965 );
and ( n29967 , n28843 , n28844 );
and ( n29968 , n28845 , n28848 );
or ( n29969 , n29967 , n29968 );
xor ( n29970 , n29966 , n29969 );
nor ( n29971 , n796 , n23541 );
xor ( n29972 , n29970 , n29971 );
and ( n29973 , n28849 , n28850 );
and ( n29974 , n28851 , n28854 );
or ( n29975 , n29973 , n29974 );
xor ( n29976 , n29972 , n29975 );
nor ( n29977 , n868 , n22541 );
xor ( n29978 , n29976 , n29977 );
and ( n29979 , n28855 , n28856 );
and ( n29980 , n28857 , n28860 );
or ( n29981 , n29979 , n29980 );
xor ( n29982 , n29978 , n29981 );
nor ( n29983 , n958 , n21562 );
xor ( n29984 , n29982 , n29983 );
and ( n29985 , n28861 , n28862 );
and ( n29986 , n28863 , n28866 );
or ( n29987 , n29985 , n29986 );
xor ( n29988 , n29984 , n29987 );
nor ( n29989 , n1062 , n20601 );
xor ( n29990 , n29988 , n29989 );
and ( n29991 , n28867 , n28868 );
and ( n29992 , n28869 , n28872 );
or ( n29993 , n29991 , n29992 );
xor ( n29994 , n29990 , n29993 );
nor ( n29995 , n1176 , n19657 );
xor ( n29996 , n29994 , n29995 );
and ( n29997 , n28873 , n28874 );
and ( n29998 , n28875 , n28878 );
or ( n29999 , n29997 , n29998 );
xor ( n30000 , n29996 , n29999 );
nor ( n30001 , n1303 , n18734 );
xor ( n30002 , n30000 , n30001 );
and ( n30003 , n28879 , n28880 );
and ( n30004 , n28881 , n28884 );
or ( n30005 , n30003 , n30004 );
xor ( n30006 , n30002 , n30005 );
nor ( n30007 , n1445 , n17828 );
xor ( n30008 , n30006 , n30007 );
and ( n30009 , n28885 , n28886 );
and ( n30010 , n28887 , n28890 );
or ( n30011 , n30009 , n30010 );
xor ( n30012 , n30008 , n30011 );
nor ( n30013 , n1598 , n16943 );
xor ( n30014 , n30012 , n30013 );
and ( n30015 , n28891 , n28892 );
and ( n30016 , n28893 , n28896 );
or ( n30017 , n30015 , n30016 );
xor ( n30018 , n30014 , n30017 );
nor ( n30019 , n1766 , n16077 );
xor ( n30020 , n30018 , n30019 );
and ( n30021 , n28897 , n28898 );
and ( n30022 , n28899 , n28902 );
or ( n30023 , n30021 , n30022 );
xor ( n30024 , n30020 , n30023 );
nor ( n30025 , n1945 , n15230 );
xor ( n30026 , n30024 , n30025 );
and ( n30027 , n28903 , n28904 );
and ( n30028 , n28905 , n28908 );
or ( n30029 , n30027 , n30028 );
xor ( n30030 , n30026 , n30029 );
nor ( n30031 , n2137 , n14403 );
xor ( n30032 , n30030 , n30031 );
and ( n30033 , n28909 , n28910 );
and ( n30034 , n28911 , n28914 );
or ( n30035 , n30033 , n30034 );
xor ( n30036 , n30032 , n30035 );
nor ( n30037 , n2343 , n13599 );
xor ( n30038 , n30036 , n30037 );
and ( n30039 , n28915 , n28916 );
and ( n30040 , n28917 , n28920 );
or ( n30041 , n30039 , n30040 );
xor ( n30042 , n30038 , n30041 );
nor ( n30043 , n2566 , n12808 );
xor ( n30044 , n30042 , n30043 );
and ( n30045 , n28921 , n28922 );
and ( n30046 , n28923 , n28926 );
or ( n30047 , n30045 , n30046 );
xor ( n30048 , n30044 , n30047 );
nor ( n30049 , n2797 , n12037 );
xor ( n30050 , n30048 , n30049 );
and ( n30051 , n28927 , n28928 );
and ( n30052 , n28929 , n28932 );
or ( n30053 , n30051 , n30052 );
xor ( n30054 , n30050 , n30053 );
nor ( n30055 , n3043 , n11282 );
xor ( n30056 , n30054 , n30055 );
and ( n30057 , n28933 , n28934 );
and ( n30058 , n28935 , n28938 );
or ( n30059 , n30057 , n30058 );
xor ( n30060 , n30056 , n30059 );
nor ( n30061 , n3300 , n10547 );
xor ( n30062 , n30060 , n30061 );
and ( n30063 , n28939 , n28940 );
and ( n30064 , n28941 , n28944 );
or ( n30065 , n30063 , n30064 );
xor ( n30066 , n30062 , n30065 );
nor ( n30067 , n3570 , n9829 );
xor ( n30068 , n30066 , n30067 );
and ( n30069 , n28945 , n28946 );
and ( n30070 , n28947 , n28950 );
or ( n30071 , n30069 , n30070 );
xor ( n30072 , n30068 , n30071 );
nor ( n30073 , n3853 , n8955 );
xor ( n30074 , n30072 , n30073 );
and ( n30075 , n28951 , n28952 );
and ( n30076 , n28953 , n28956 );
or ( n30077 , n30075 , n30076 );
xor ( n30078 , n30074 , n30077 );
nor ( n30079 , n4151 , n603 );
xor ( n30080 , n30078 , n30079 );
and ( n30081 , n28957 , n28958 );
and ( n30082 , n28959 , n28962 );
or ( n30083 , n30081 , n30082 );
xor ( n30084 , n30080 , n30083 );
nor ( n30085 , n4458 , n652 );
xor ( n30086 , n30084 , n30085 );
and ( n30087 , n28963 , n28964 );
and ( n30088 , n28965 , n28968 );
or ( n30089 , n30087 , n30088 );
xor ( n30090 , n30086 , n30089 );
nor ( n30091 , n4786 , n624 );
xor ( n30092 , n30090 , n30091 );
and ( n30093 , n28969 , n28970 );
and ( n30094 , n28971 , n28974 );
or ( n30095 , n30093 , n30094 );
xor ( n30096 , n30092 , n30095 );
nor ( n30097 , n5126 , n648 );
xor ( n30098 , n30096 , n30097 );
and ( n30099 , n28975 , n28976 );
and ( n30100 , n28977 , n28980 );
or ( n30101 , n30099 , n30100 );
xor ( n30102 , n30098 , n30101 );
nor ( n30103 , n5477 , n686 );
xor ( n30104 , n30102 , n30103 );
and ( n30105 , n28981 , n28982 );
and ( n30106 , n28983 , n28986 );
or ( n30107 , n30105 , n30106 );
xor ( n30108 , n30104 , n30107 );
nor ( n30109 , n5838 , n735 );
xor ( n30110 , n30108 , n30109 );
and ( n30111 , n28987 , n28988 );
and ( n30112 , n28989 , n28992 );
or ( n30113 , n30111 , n30112 );
xor ( n30114 , n30110 , n30113 );
nor ( n30115 , n6212 , n798 );
xor ( n30116 , n30114 , n30115 );
and ( n30117 , n28993 , n28994 );
and ( n30118 , n28995 , n28998 );
or ( n30119 , n30117 , n30118 );
xor ( n30120 , n30116 , n30119 );
nor ( n30121 , n6596 , n870 );
xor ( n30122 , n30120 , n30121 );
and ( n30123 , n28999 , n29000 );
and ( n30124 , n29001 , n29004 );
or ( n30125 , n30123 , n30124 );
xor ( n30126 , n30122 , n30125 );
nor ( n30127 , n6997 , n960 );
xor ( n30128 , n30126 , n30127 );
and ( n30129 , n29005 , n29006 );
and ( n30130 , n29007 , n29010 );
or ( n30131 , n30129 , n30130 );
xor ( n30132 , n30128 , n30131 );
nor ( n30133 , n7413 , n1064 );
xor ( n30134 , n30132 , n30133 );
and ( n30135 , n29011 , n29012 );
and ( n30136 , n29013 , n29016 );
or ( n30137 , n30135 , n30136 );
xor ( n30138 , n30134 , n30137 );
nor ( n30139 , n7841 , n1178 );
xor ( n30140 , n30138 , n30139 );
and ( n30141 , n29017 , n29018 );
and ( n30142 , n29019 , n29022 );
or ( n30143 , n30141 , n30142 );
xor ( n30144 , n30140 , n30143 );
nor ( n30145 , n8281 , n1305 );
xor ( n30146 , n30144 , n30145 );
and ( n30147 , n29023 , n29024 );
and ( n30148 , n29025 , n29028 );
or ( n30149 , n30147 , n30148 );
xor ( n30150 , n30146 , n30149 );
nor ( n30151 , n8737 , n1447 );
xor ( n30152 , n30150 , n30151 );
and ( n30153 , n29029 , n29030 );
and ( n30154 , n29031 , n29034 );
or ( n30155 , n30153 , n30154 );
xor ( n30156 , n30152 , n30155 );
nor ( n30157 , n9420 , n1600 );
xor ( n30158 , n30156 , n30157 );
and ( n30159 , n29035 , n29036 );
and ( n30160 , n29037 , n29040 );
or ( n30161 , n30159 , n30160 );
xor ( n30162 , n30158 , n30161 );
nor ( n30163 , n10312 , n1768 );
xor ( n30164 , n30162 , n30163 );
and ( n30165 , n29041 , n29042 );
and ( n30166 , n29043 , n29046 );
or ( n30167 , n30165 , n30166 );
xor ( n30168 , n30164 , n30167 );
nor ( n30169 , n11041 , n1947 );
xor ( n30170 , n30168 , n30169 );
and ( n30171 , n29047 , n29048 );
and ( n30172 , n29049 , n29052 );
or ( n30173 , n30171 , n30172 );
xor ( n30174 , n30170 , n30173 );
nor ( n30175 , n11790 , n2139 );
xor ( n30176 , n30174 , n30175 );
and ( n30177 , n29053 , n29054 );
and ( n30178 , n29055 , n29058 );
or ( n30179 , n30177 , n30178 );
xor ( n30180 , n30176 , n30179 );
nor ( n30181 , n12555 , n2345 );
xor ( n30182 , n30180 , n30181 );
and ( n30183 , n29059 , n29060 );
and ( n30184 , n29061 , n29064 );
or ( n30185 , n30183 , n30184 );
xor ( n30186 , n30182 , n30185 );
nor ( n30187 , n13340 , n2568 );
xor ( n30188 , n30186 , n30187 );
and ( n30189 , n29065 , n29066 );
and ( n30190 , n29067 , n29070 );
or ( n30191 , n30189 , n30190 );
xor ( n30192 , n30188 , n30191 );
nor ( n30193 , n14138 , n2799 );
xor ( n30194 , n30192 , n30193 );
and ( n30195 , n29071 , n29072 );
and ( n30196 , n29073 , n29076 );
or ( n30197 , n30195 , n30196 );
xor ( n30198 , n30194 , n30197 );
nor ( n30199 , n14959 , n3045 );
xor ( n30200 , n30198 , n30199 );
and ( n30201 , n29077 , n29078 );
and ( n30202 , n29079 , n29082 );
or ( n30203 , n30201 , n30202 );
xor ( n30204 , n30200 , n30203 );
nor ( n30205 , n15800 , n3302 );
xor ( n30206 , n30204 , n30205 );
and ( n30207 , n29083 , n29084 );
and ( n30208 , n29085 , n29088 );
or ( n30209 , n30207 , n30208 );
xor ( n30210 , n30206 , n30209 );
nor ( n30211 , n16660 , n3572 );
xor ( n30212 , n30210 , n30211 );
and ( n30213 , n29089 , n29090 );
and ( n30214 , n29091 , n29094 );
or ( n30215 , n30213 , n30214 );
xor ( n30216 , n30212 , n30215 );
nor ( n30217 , n17539 , n3855 );
xor ( n30218 , n30216 , n30217 );
and ( n30219 , n29095 , n29096 );
and ( n30220 , n29097 , n29100 );
or ( n30221 , n30219 , n30220 );
xor ( n30222 , n30218 , n30221 );
nor ( n30223 , n18439 , n4153 );
xor ( n30224 , n30222 , n30223 );
and ( n30225 , n29101 , n29102 );
and ( n30226 , n29103 , n29106 );
or ( n30227 , n30225 , n30226 );
xor ( n30228 , n30224 , n30227 );
nor ( n30229 , n19356 , n4460 );
xor ( n30230 , n30228 , n30229 );
and ( n30231 , n29107 , n29108 );
and ( n30232 , n29109 , n29112 );
or ( n30233 , n30231 , n30232 );
xor ( n30234 , n30230 , n30233 );
nor ( n30235 , n20294 , n4788 );
xor ( n30236 , n30234 , n30235 );
and ( n30237 , n29113 , n29114 );
and ( n30238 , n29115 , n29118 );
or ( n30239 , n30237 , n30238 );
xor ( n30240 , n30236 , n30239 );
nor ( n30241 , n21249 , n5128 );
xor ( n30242 , n30240 , n30241 );
and ( n30243 , n29119 , n29120 );
and ( n30244 , n29121 , n29124 );
or ( n30245 , n30243 , n30244 );
xor ( n30246 , n30242 , n30245 );
nor ( n30247 , n22222 , n5479 );
xor ( n30248 , n30246 , n30247 );
and ( n30249 , n29125 , n29126 );
and ( n30250 , n29127 , n29130 );
or ( n30251 , n30249 , n30250 );
xor ( n30252 , n30248 , n30251 );
nor ( n30253 , n23216 , n5840 );
xor ( n30254 , n30252 , n30253 );
and ( n30255 , n29131 , n29132 );
and ( n30256 , n29133 , n29136 );
or ( n30257 , n30255 , n30256 );
xor ( n30258 , n30254 , n30257 );
nor ( n30259 , n24233 , n6214 );
xor ( n30260 , n30258 , n30259 );
and ( n30261 , n29137 , n29138 );
and ( n30262 , n29139 , n29142 );
or ( n30263 , n30261 , n30262 );
xor ( n30264 , n30260 , n30263 );
nor ( n30265 , n25263 , n6598 );
xor ( n30266 , n30264 , n30265 );
and ( n30267 , n29143 , n29144 );
and ( n30268 , n29145 , n29148 );
or ( n30269 , n30267 , n30268 );
xor ( n30270 , n30266 , n30269 );
nor ( n30271 , n26317 , n6999 );
xor ( n30272 , n30270 , n30271 );
and ( n30273 , n29149 , n29150 );
and ( n30274 , n29151 , n29154 );
or ( n30275 , n30273 , n30274 );
xor ( n30276 , n30272 , n30275 );
nor ( n30277 , n27388 , n7415 );
xor ( n30278 , n30276 , n30277 );
and ( n30279 , n29155 , n29156 );
and ( n30280 , n29157 , n29160 );
or ( n30281 , n30279 , n30280 );
xor ( n30282 , n30278 , n30281 );
nor ( n30283 , n28478 , n7843 );
xor ( n30284 , n30282 , n30283 );
and ( n30285 , n29161 , n29162 );
and ( n30286 , n29163 , n29166 );
or ( n30287 , n30285 , n30286 );
xor ( n30288 , n30284 , n30287 );
nor ( n30289 , n29587 , n8283 );
xor ( n30290 , n30288 , n30289 );
and ( n30291 , n29167 , n29168 );
and ( n30292 , n29169 , n29172 );
or ( n30293 , n30291 , n30292 );
xor ( n30294 , n30290 , n30293 );
and ( n30295 , n29524 , n29525 );
and ( n30296 , n29525 , n29572 );
and ( n30297 , n29524 , n29572 );
or ( n30298 , n30295 , n30296 , n30297 );
and ( n30299 , n29186 , n29519 );
and ( n30300 , n29519 , n29573 );
and ( n30301 , n29186 , n29573 );
or ( n30302 , n30299 , n30300 , n30301 );
xor ( n30303 , n30298 , n30302 );
and ( n30304 , n29190 , n29310 );
and ( n30305 , n29310 , n29518 );
and ( n30306 , n29190 , n29518 );
or ( n30307 , n30304 , n30305 , n30306 );
and ( n30308 , n29315 , n29393 );
and ( n30309 , n29393 , n29517 );
and ( n30310 , n29315 , n29517 );
or ( n30311 , n30308 , n30309 , n30310 );
and ( n30312 , n29203 , n29271 );
and ( n30313 , n29271 , n29308 );
and ( n30314 , n29203 , n29308 );
or ( n30315 , n30312 , n30313 , n30314 );
and ( n30316 , n29319 , n29323 );
and ( n30317 , n29323 , n29392 );
and ( n30318 , n29319 , n29392 );
or ( n30319 , n30316 , n30317 , n30318 );
xor ( n30320 , n30315 , n30319 );
and ( n30321 , n29276 , n29280 );
and ( n30322 , n29280 , n29307 );
and ( n30323 , n29276 , n29307 );
or ( n30324 , n30321 , n30322 , n30323 );
and ( n30325 , n29237 , n29253 );
and ( n30326 , n29253 , n29269 );
and ( n30327 , n29237 , n29269 );
or ( n30328 , n30325 , n30326 , n30327 );
and ( n30329 , n29220 , n29224 );
and ( n30330 , n29224 , n29230 );
and ( n30331 , n29220 , n29230 );
or ( n30332 , n30329 , n30330 , n30331 );
and ( n30333 , n29241 , n29246 );
and ( n30334 , n29246 , n29252 );
and ( n30335 , n29241 , n29252 );
or ( n30336 , n30333 , n30334 , n30335 );
xor ( n30337 , n30332 , n30336 );
and ( n30338 , n29226 , n29227 );
and ( n30339 , n29227 , n29229 );
and ( n30340 , n29226 , n29229 );
or ( n30341 , n30338 , n30339 , n30340 );
and ( n30342 , n29242 , n29243 );
and ( n30343 , n29243 , n29245 );
and ( n30344 , n29242 , n29245 );
or ( n30345 , n30342 , n30343 , n30344 );
xor ( n30346 , n30341 , n30345 );
and ( n30347 , n21216 , n1034 );
and ( n30348 , n22186 , n940 );
xor ( n30349 , n30347 , n30348 );
and ( n30350 , n22892 , n840 );
xor ( n30351 , n30349 , n30350 );
xor ( n30352 , n30346 , n30351 );
xor ( n30353 , n30337 , n30352 );
xor ( n30354 , n30328 , n30353 );
and ( n30355 , n29258 , n29262 );
and ( n30356 , n29262 , n29268 );
and ( n30357 , n29258 , n29268 );
or ( n30358 , n30355 , n30356 , n30357 );
and ( n30359 , n29248 , n29249 );
and ( n30360 , n29249 , n29251 );
and ( n30361 , n29248 , n29251 );
or ( n30362 , n30359 , n30360 , n30361 );
and ( n30363 , n18144 , n1424 );
and ( n30364 , n19324 , n1254 );
xor ( n30365 , n30363 , n30364 );
and ( n30366 , n20233 , n1134 );
xor ( n30367 , n30365 , n30366 );
xor ( n30368 , n30362 , n30367 );
and ( n30369 , n15758 , n1882 );
and ( n30370 , n16637 , n1738 );
xor ( n30371 , n30369 , n30370 );
and ( n30372 , n17512 , n1551 );
xor ( n30373 , n30371 , n30372 );
xor ( n30374 , n30368 , n30373 );
xor ( n30375 , n30358 , n30374 );
and ( n30376 , n29264 , n29265 );
and ( n30377 , n29265 , n29267 );
and ( n30378 , n29264 , n29267 );
or ( n30379 , n30376 , n30377 , n30378 );
and ( n30380 , n29295 , n29296 );
and ( n30381 , n29296 , n29298 );
and ( n30382 , n29295 , n29298 );
or ( n30383 , n30380 , n30381 , n30382 );
xor ( n30384 , n30379 , n30383 );
and ( n30385 , n13322 , n2544 );
and ( n30386 , n14118 , n2298 );
xor ( n30387 , n30385 , n30386 );
and ( n30388 , n14938 , n2100 );
xor ( n30389 , n30387 , n30388 );
xor ( n30390 , n30384 , n30389 );
xor ( n30391 , n30375 , n30390 );
xor ( n30392 , n30354 , n30391 );
xor ( n30393 , n30324 , n30392 );
and ( n30394 , n29285 , n29289 );
and ( n30395 , n29289 , n29306 );
and ( n30396 , n29285 , n29306 );
or ( n30397 , n30394 , n30395 , n30396 );
and ( n30398 , n29332 , n29347 );
and ( n30399 , n29347 , n29364 );
and ( n30400 , n29332 , n29364 );
or ( n30401 , n30398 , n30399 , n30400 );
xor ( n30402 , n30397 , n30401 );
and ( n30403 , n29294 , n29299 );
and ( n30404 , n29299 , n29305 );
and ( n30405 , n29294 , n29305 );
or ( n30406 , n30403 , n30404 , n30405 );
and ( n30407 , n29336 , n29340 );
and ( n30408 , n29340 , n29346 );
and ( n30409 , n29336 , n29346 );
or ( n30410 , n30407 , n30408 , n30409 );
xor ( n30411 , n30406 , n30410 );
and ( n30412 , n29301 , n29302 );
and ( n30413 , n29302 , n29304 );
and ( n30414 , n29301 , n29304 );
or ( n30415 , n30412 , n30413 , n30414 );
and ( n30416 , n11015 , n3271 );
and ( n30417 , n11769 , n2981 );
xor ( n30418 , n30416 , n30417 );
and ( n30419 , n12320 , n2739 );
xor ( n30420 , n30418 , n30419 );
xor ( n30421 , n30415 , n30420 );
and ( n30422 , n8718 , n4102 );
and ( n30423 , n9400 , n3749 );
xor ( n30424 , n30422 , n30423 );
and ( n30425 , n10291 , n3495 );
xor ( n30426 , n30424 , n30425 );
xor ( n30427 , n30421 , n30426 );
xor ( n30428 , n30411 , n30427 );
xor ( n30429 , n30402 , n30428 );
xor ( n30430 , n30393 , n30429 );
xor ( n30431 , n30320 , n30430 );
xor ( n30432 , n30311 , n30431 );
and ( n30433 , n29398 , n29445 );
and ( n30434 , n29445 , n29516 );
and ( n30435 , n29398 , n29516 );
or ( n30436 , n30433 , n30434 , n30435 );
and ( n30437 , n29328 , n29365 );
and ( n30438 , n29365 , n29391 );
and ( n30439 , n29328 , n29391 );
or ( n30440 , n30437 , n30438 , n30439 );
and ( n30441 , n29402 , n29406 );
and ( n30442 , n29406 , n29444 );
and ( n30443 , n29402 , n29444 );
or ( n30444 , n30441 , n30442 , n30443 );
xor ( n30445 , n30440 , n30444 );
and ( n30446 , n29370 , n29374 );
and ( n30447 , n29374 , n29390 );
and ( n30448 , n29370 , n29390 );
or ( n30449 , n30446 , n30447 , n30448 );
and ( n30450 , n29352 , n29357 );
and ( n30451 , n29357 , n29363 );
and ( n30452 , n29352 , n29363 );
or ( n30453 , n30450 , n30451 , n30452 );
and ( n30454 , n29342 , n29343 );
and ( n30455 , n29343 , n29345 );
and ( n30456 , n29342 , n29345 );
or ( n30457 , n30454 , n30455 , n30456 );
and ( n30458 , n29353 , n29354 );
and ( n30459 , n29354 , n29356 );
and ( n30460 , n29353 , n29356 );
or ( n30461 , n30458 , n30459 , n30460 );
xor ( n30462 , n30457 , n30461 );
and ( n30463 , n7385 , n5103 );
and ( n30464 , n7808 , n4730 );
xor ( n30465 , n30463 , n30464 );
and ( n30466 , n8079 , n4403 );
xor ( n30467 , n30465 , n30466 );
xor ( n30468 , n30462 , n30467 );
xor ( n30469 , n30453 , n30468 );
and ( n30470 , n29359 , n29360 );
and ( n30471 , n29360 , n29362 );
and ( n30472 , n29359 , n29362 );
or ( n30473 , n30470 , n30471 , n30472 );
buf ( n30474 , n6187 );
and ( n30475 , n6569 , n5765 );
xor ( n30476 , n30474 , n30475 );
and ( n30477 , n6816 , n5408 );
xor ( n30478 , n30476 , n30477 );
xor ( n30479 , n30473 , n30478 );
and ( n30480 , n4959 , n7310 );
and ( n30481 , n5459 , n6971 );
xor ( n30482 , n30480 , n30481 );
and ( n30483 , n5819 , n6504 );
xor ( n30484 , n30482 , n30483 );
xor ( n30485 , n30479 , n30484 );
xor ( n30486 , n30469 , n30485 );
xor ( n30487 , n30449 , n30486 );
and ( n30488 , n29379 , n29383 );
and ( n30489 , n29383 , n29389 );
and ( n30490 , n29379 , n29389 );
or ( n30491 , n30488 , n30489 , n30490 );
and ( n30492 , n29415 , n29420 );
and ( n30493 , n29420 , n29426 );
and ( n30494 , n29415 , n29426 );
or ( n30495 , n30492 , n30493 , n30494 );
xor ( n30496 , n30491 , n30495 );
and ( n30497 , n29385 , n29386 );
and ( n30498 , n29386 , n29388 );
and ( n30499 , n29385 , n29388 );
or ( n30500 , n30497 , n30498 , n30499 );
and ( n30501 , n29416 , n29417 );
and ( n30502 , n29417 , n29419 );
and ( n30503 , n29416 , n29419 );
or ( n30504 , n30501 , n30502 , n30503 );
xor ( n30505 , n30500 , n30504 );
and ( n30506 , n4132 , n8669 );
and ( n30507 , n4438 , n8243 );
xor ( n30508 , n30506 , n30507 );
and ( n30509 , n4766 , n7662 );
xor ( n30510 , n30508 , n30509 );
xor ( n30511 , n30505 , n30510 );
xor ( n30512 , n30496 , n30511 );
xor ( n30513 , n30487 , n30512 );
xor ( n30514 , n30445 , n30513 );
xor ( n30515 , n30436 , n30514 );
and ( n30516 , n29450 , n29476 );
and ( n30517 , n29476 , n29515 );
and ( n30518 , n29450 , n29515 );
or ( n30519 , n30516 , n30517 , n30518 );
and ( n30520 , n29411 , n29427 );
and ( n30521 , n29427 , n29443 );
and ( n30522 , n29411 , n29443 );
or ( n30523 , n30520 , n30521 , n30522 );
and ( n30524 , n29454 , n29458 );
and ( n30525 , n29458 , n29475 );
and ( n30526 , n29454 , n29475 );
or ( n30527 , n30524 , n30525 , n30526 );
xor ( n30528 , n30523 , n30527 );
and ( n30529 , n29432 , n29436 );
and ( n30530 , n29436 , n29442 );
and ( n30531 , n29432 , n29442 );
or ( n30532 , n30529 , n30530 , n30531 );
and ( n30533 , n29422 , n29423 );
and ( n30534 , n29423 , n29425 );
and ( n30535 , n29422 , n29425 );
or ( n30536 , n30533 , n30534 , n30535 );
and ( n30537 , n3182 , n10977 );
and ( n30538 , n3545 , n10239 );
xor ( n30539 , n30537 , n30538 );
and ( n30540 , n3801 , n9348 );
xor ( n30541 , n30539 , n30540 );
xor ( n30542 , n30536 , n30541 );
and ( n30543 , n2462 , n13256 );
and ( n30544 , n2779 , n12531 );
xor ( n30545 , n30543 , n30544 );
and ( n30546 , n3024 , n11718 );
xor ( n30547 , n30545 , n30546 );
xor ( n30548 , n30542 , n30547 );
xor ( n30549 , n30532 , n30548 );
and ( n30550 , n29438 , n29439 );
and ( n30551 , n29439 , n29441 );
and ( n30552 , n29438 , n29441 );
or ( n30553 , n30550 , n30551 , n30552 );
and ( n30554 , n29464 , n29465 );
and ( n30555 , n29465 , n29467 );
and ( n30556 , n29464 , n29467 );
or ( n30557 , n30554 , n30555 , n30556 );
xor ( n30558 , n30553 , n30557 );
and ( n30559 , n1933 , n15691 );
and ( n30560 , n2120 , n14838 );
xor ( n30561 , n30559 , n30560 );
and ( n30562 , n2324 , n14044 );
xor ( n30563 , n30561 , n30562 );
xor ( n30564 , n30558 , n30563 );
xor ( n30565 , n30549 , n30564 );
xor ( n30566 , n30528 , n30565 );
xor ( n30567 , n30519 , n30566 );
and ( n30568 , n29481 , n29496 );
and ( n30569 , n29496 , n29514 );
and ( n30570 , n29481 , n29514 );
or ( n30571 , n30568 , n30569 , n30570 );
and ( n30572 , n29463 , n29468 );
and ( n30573 , n29468 , n29474 );
and ( n30574 , n29463 , n29474 );
or ( n30575 , n30572 , n30573 , n30574 );
and ( n30576 , n29485 , n29489 );
and ( n30577 , n29489 , n29495 );
and ( n30578 , n29485 , n29495 );
or ( n30579 , n30576 , n30577 , n30578 );
xor ( n30580 , n30575 , n30579 );
and ( n30581 , n29470 , n29471 );
and ( n30582 , n29471 , n29473 );
and ( n30583 , n29470 , n29473 );
or ( n30584 , n30581 , n30582 , n30583 );
and ( n30585 , n1383 , n18407 );
and ( n30586 , n1580 , n17422 );
xor ( n30587 , n30585 , n30586 );
and ( n30588 , n1694 , n16550 );
xor ( n30589 , n30587 , n30588 );
xor ( n30590 , n30584 , n30589 );
and ( n30591 , n1047 , n20976 );
and ( n30592 , n1164 , n20156 );
xor ( n30593 , n30591 , n30592 );
and ( n30594 , n1287 , n19222 );
xor ( n30595 , n30593 , n30594 );
xor ( n30596 , n30590 , n30595 );
xor ( n30597 , n30580 , n30596 );
xor ( n30598 , n30571 , n30597 );
and ( n30599 , n29501 , n29506 );
and ( n30600 , n29506 , n29513 );
and ( n30601 , n29501 , n29513 );
or ( n30602 , n30599 , n30600 , n30601 );
and ( n30603 , n29491 , n29492 );
and ( n30604 , n29492 , n29494 );
and ( n30605 , n29491 , n29494 );
or ( n30606 , n30603 , n30604 , n30605 );
and ( n30607 , n29502 , n29503 );
and ( n30608 , n29503 , n29505 );
and ( n30609 , n29502 , n29505 );
or ( n30610 , n30607 , n30608 , n30609 );
xor ( n30611 , n30606 , n30610 );
and ( n30612 , n783 , n24137 );
and ( n30613 , n856 , n23075 );
xor ( n30614 , n30612 , n30613 );
and ( n30615 , n925 , n22065 );
xor ( n30616 , n30614 , n30615 );
xor ( n30617 , n30611 , n30616 );
xor ( n30618 , n30602 , n30617 );
and ( n30619 , n29509 , n29510 );
and ( n30620 , n29510 , n29512 );
and ( n30621 , n29509 , n29512 );
or ( n30622 , n30619 , n30620 , n30621 );
and ( n30623 , n632 , n27296 );
and ( n30624 , n671 , n26216 );
xor ( n30625 , n30623 , n30624 );
and ( n30626 , n715 , n25163 );
xor ( n30627 , n30625 , n30626 );
xor ( n30628 , n30622 , n30627 );
buf ( n30629 , n410 );
and ( n30630 , n599 , n30629 );
and ( n30631 , n608 , n29508 );
xor ( n30632 , n30630 , n30631 );
and ( n30633 , n611 , n28406 );
xor ( n30634 , n30632 , n30633 );
xor ( n30635 , n30628 , n30634 );
xor ( n30636 , n30618 , n30635 );
xor ( n30637 , n30598 , n30636 );
xor ( n30638 , n30567 , n30637 );
xor ( n30639 , n30515 , n30638 );
xor ( n30640 , n30432 , n30639 );
xor ( n30641 , n30307 , n30640 );
and ( n30642 , n29194 , n29198 );
and ( n30643 , n29198 , n29309 );
and ( n30644 , n29194 , n29309 );
or ( n30645 , n30642 , n30643 , n30644 );
and ( n30646 , n29530 , n29571 );
xor ( n30647 , n30645 , n30646 );
and ( n30648 , n29534 , n29538 );
and ( n30649 , n29538 , n29570 );
and ( n30650 , n29534 , n29570 );
or ( n30651 , n30648 , n30649 , n30650 );
and ( n30652 , n29543 , n29544 );
and ( n30653 , n29544 , n29569 );
and ( n30654 , n29543 , n29569 );
or ( n30655 , n30652 , n30653 , n30654 );
and ( n30656 , n29207 , n29232 );
and ( n30657 , n29232 , n29270 );
and ( n30658 , n29207 , n29270 );
or ( n30659 , n30656 , n30657 , n30658 );
xor ( n30660 , n30655 , n30659 );
and ( n30661 , n29546 , n29550 );
and ( n30662 , n29550 , n29568 );
and ( n30663 , n29546 , n29568 );
or ( n30664 , n30661 , n30662 , n30663 );
and ( n30665 , n29211 , n29215 );
and ( n30666 , n29215 , n29231 );
and ( n30667 , n29211 , n29231 );
or ( n30668 , n30665 , n30666 , n30667 );
xor ( n30669 , n30664 , n30668 );
and ( n30670 , n29555 , n29561 );
and ( n30671 , n29561 , n29567 );
and ( n30672 , n29555 , n29567 );
or ( n30673 , n30670 , n30671 , n30672 );
and ( n30674 , n29563 , n29564 );
and ( n30675 , n29564 , n29566 );
and ( n30676 , n29563 , n29566 );
or ( n30677 , n30674 , n30675 , n30676 );
and ( n30678 , n27361 , n635 );
and ( n30679 , n28456 , n606 );
xor ( n30680 , n30678 , n30679 );
and ( n30681 , n29559 , n615 );
xor ( n30682 , n30680 , n30681 );
xor ( n30683 , n30677 , n30682 );
and ( n30684 , n24214 , n771 );
and ( n30685 , n25243 , n719 );
xor ( n30686 , n30684 , n30685 );
and ( n30687 , n26296 , n663 );
xor ( n30688 , n30686 , n30687 );
xor ( n30689 , n30683 , n30688 );
xor ( n30690 , n30673 , n30689 );
and ( n30691 , n29556 , n29557 );
and ( n30692 , n29557 , n29560 );
and ( n30693 , n29556 , n29560 );
or ( n30694 , n30691 , n30692 , n30693 );
buf ( n30695 , n410 );
and ( n30696 , n30695 , n612 );
xor ( n30697 , n30694 , n30696 );
xor ( n30698 , n30690 , n30697 );
xor ( n30699 , n30669 , n30698 );
xor ( n30700 , n30660 , n30699 );
xor ( n30701 , n30651 , n30700 );
xor ( n30702 , n30647 , n30701 );
xor ( n30703 , n30641 , n30702 );
xor ( n30704 , n30303 , n30703 );
and ( n30705 , n29177 , n29181 );
and ( n30706 , n29181 , n29574 );
and ( n30707 , n29177 , n29574 );
or ( n30708 , n30705 , n30706 , n30707 );
xor ( n30709 , n30704 , n30708 );
and ( n30710 , n29575 , n29579 );
and ( n30711 , n29580 , n29583 );
or ( n30712 , n30710 , n30711 );
xor ( n30713 , n30709 , n30712 );
buf ( n30714 , n30713 );
buf ( n30715 , n30714 );
not ( n30716 , n30715 );
nor ( n30717 , n30716 , n8739 );
xor ( n30718 , n30294 , n30717 );
and ( n30719 , n29173 , n29588 );
and ( n30720 , n29589 , n29592 );
or ( n30721 , n30719 , n30720 );
xor ( n30722 , n30718 , n30721 );
buf ( n30723 , n30722 );
buf ( n30724 , n30723 );
not ( n30725 , n30724 );
buf ( n30726 , n559 );
not ( n30727 , n30726 );
nor ( n30728 , n30725 , n30727 );
xor ( n30729 , n29946 , n30728 );
xor ( n30730 , n29604 , n29943 );
nor ( n30731 , n29596 , n30727 );
and ( n30732 , n30730 , n30731 );
xor ( n30733 , n30730 , n30731 );
xor ( n30734 , n29608 , n29941 );
nor ( n30735 , n28487 , n30727 );
and ( n30736 , n30734 , n30735 );
xor ( n30737 , n30734 , n30735 );
xor ( n30738 , n29612 , n29939 );
nor ( n30739 , n27397 , n30727 );
and ( n30740 , n30738 , n30739 );
xor ( n30741 , n30738 , n30739 );
xor ( n30742 , n29616 , n29937 );
nor ( n30743 , n26326 , n30727 );
and ( n30744 , n30742 , n30743 );
xor ( n30745 , n30742 , n30743 );
xor ( n30746 , n29620 , n29935 );
nor ( n30747 , n25272 , n30727 );
and ( n30748 , n30746 , n30747 );
xor ( n30749 , n30746 , n30747 );
xor ( n30750 , n29624 , n29933 );
nor ( n30751 , n24242 , n30727 );
and ( n30752 , n30750 , n30751 );
xor ( n30753 , n30750 , n30751 );
xor ( n30754 , n29628 , n29931 );
nor ( n30755 , n23225 , n30727 );
and ( n30756 , n30754 , n30755 );
xor ( n30757 , n30754 , n30755 );
xor ( n30758 , n29632 , n29929 );
nor ( n30759 , n22231 , n30727 );
and ( n30760 , n30758 , n30759 );
xor ( n30761 , n30758 , n30759 );
xor ( n30762 , n29636 , n29927 );
nor ( n30763 , n21258 , n30727 );
and ( n30764 , n30762 , n30763 );
xor ( n30765 , n30762 , n30763 );
xor ( n30766 , n29640 , n29925 );
nor ( n30767 , n20303 , n30727 );
and ( n30768 , n30766 , n30767 );
xor ( n30769 , n30766 , n30767 );
xor ( n30770 , n29644 , n29923 );
nor ( n30771 , n19365 , n30727 );
and ( n30772 , n30770 , n30771 );
xor ( n30773 , n30770 , n30771 );
xor ( n30774 , n29648 , n29921 );
nor ( n30775 , n18448 , n30727 );
and ( n30776 , n30774 , n30775 );
xor ( n30777 , n30774 , n30775 );
xor ( n30778 , n29652 , n29919 );
nor ( n30779 , n17548 , n30727 );
and ( n30780 , n30778 , n30779 );
xor ( n30781 , n30778 , n30779 );
xor ( n30782 , n29656 , n29917 );
nor ( n30783 , n16669 , n30727 );
and ( n30784 , n30782 , n30783 );
xor ( n30785 , n30782 , n30783 );
xor ( n30786 , n29660 , n29915 );
nor ( n30787 , n15809 , n30727 );
and ( n30788 , n30786 , n30787 );
xor ( n30789 , n30786 , n30787 );
xor ( n30790 , n29664 , n29913 );
nor ( n30791 , n14968 , n30727 );
and ( n30792 , n30790 , n30791 );
xor ( n30793 , n30790 , n30791 );
xor ( n30794 , n29668 , n29911 );
nor ( n30795 , n14147 , n30727 );
and ( n30796 , n30794 , n30795 );
xor ( n30797 , n30794 , n30795 );
xor ( n30798 , n29672 , n29909 );
nor ( n30799 , n13349 , n30727 );
and ( n30800 , n30798 , n30799 );
xor ( n30801 , n30798 , n30799 );
xor ( n30802 , n29676 , n29907 );
nor ( n30803 , n12564 , n30727 );
and ( n30804 , n30802 , n30803 );
xor ( n30805 , n30802 , n30803 );
xor ( n30806 , n29680 , n29905 );
nor ( n30807 , n11799 , n30727 );
and ( n30808 , n30806 , n30807 );
xor ( n30809 , n30806 , n30807 );
xor ( n30810 , n29684 , n29903 );
nor ( n30811 , n11050 , n30727 );
and ( n30812 , n30810 , n30811 );
xor ( n30813 , n30810 , n30811 );
xor ( n30814 , n29688 , n29901 );
nor ( n30815 , n10321 , n30727 );
and ( n30816 , n30814 , n30815 );
xor ( n30817 , n30814 , n30815 );
xor ( n30818 , n29692 , n29899 );
nor ( n30819 , n9429 , n30727 );
and ( n30820 , n30818 , n30819 );
xor ( n30821 , n30818 , n30819 );
xor ( n30822 , n29696 , n29897 );
nor ( n30823 , n8949 , n30727 );
and ( n30824 , n30822 , n30823 );
xor ( n30825 , n30822 , n30823 );
xor ( n30826 , n29700 , n29895 );
nor ( n30827 , n9437 , n30727 );
and ( n30828 , n30826 , n30827 );
xor ( n30829 , n30826 , n30827 );
xor ( n30830 , n29704 , n29893 );
nor ( n30831 , n9446 , n30727 );
and ( n30832 , n30830 , n30831 );
xor ( n30833 , n30830 , n30831 );
xor ( n30834 , n29708 , n29891 );
nor ( n30835 , n9455 , n30727 );
and ( n30836 , n30834 , n30835 );
xor ( n30837 , n30834 , n30835 );
xor ( n30838 , n29712 , n29889 );
nor ( n30839 , n9464 , n30727 );
and ( n30840 , n30838 , n30839 );
xor ( n30841 , n30838 , n30839 );
xor ( n30842 , n29716 , n29887 );
nor ( n30843 , n9473 , n30727 );
and ( n30844 , n30842 , n30843 );
xor ( n30845 , n30842 , n30843 );
xor ( n30846 , n29720 , n29885 );
nor ( n30847 , n9482 , n30727 );
and ( n30848 , n30846 , n30847 );
xor ( n30849 , n30846 , n30847 );
xor ( n30850 , n29724 , n29883 );
nor ( n30851 , n9491 , n30727 );
and ( n30852 , n30850 , n30851 );
xor ( n30853 , n30850 , n30851 );
xor ( n30854 , n29728 , n29881 );
nor ( n30855 , n9500 , n30727 );
and ( n30856 , n30854 , n30855 );
xor ( n30857 , n30854 , n30855 );
xor ( n30858 , n29732 , n29879 );
nor ( n30859 , n9509 , n30727 );
and ( n30860 , n30858 , n30859 );
xor ( n30861 , n30858 , n30859 );
xor ( n30862 , n29736 , n29877 );
nor ( n30863 , n9518 , n30727 );
and ( n30864 , n30862 , n30863 );
xor ( n30865 , n30862 , n30863 );
xor ( n30866 , n29740 , n29875 );
nor ( n30867 , n9527 , n30727 );
and ( n30868 , n30866 , n30867 );
xor ( n30869 , n30866 , n30867 );
xor ( n30870 , n29744 , n29873 );
nor ( n30871 , n9536 , n30727 );
and ( n30872 , n30870 , n30871 );
xor ( n30873 , n30870 , n30871 );
xor ( n30874 , n29748 , n29871 );
nor ( n30875 , n9545 , n30727 );
and ( n30876 , n30874 , n30875 );
xor ( n30877 , n30874 , n30875 );
xor ( n30878 , n29752 , n29869 );
nor ( n30879 , n9554 , n30727 );
and ( n30880 , n30878 , n30879 );
xor ( n30881 , n30878 , n30879 );
xor ( n30882 , n29756 , n29867 );
nor ( n30883 , n9563 , n30727 );
and ( n30884 , n30882 , n30883 );
xor ( n30885 , n30882 , n30883 );
xor ( n30886 , n29760 , n29865 );
nor ( n30887 , n9572 , n30727 );
and ( n30888 , n30886 , n30887 );
xor ( n30889 , n30886 , n30887 );
xor ( n30890 , n29764 , n29863 );
nor ( n30891 , n9581 , n30727 );
and ( n30892 , n30890 , n30891 );
xor ( n30893 , n30890 , n30891 );
xor ( n30894 , n29768 , n29861 );
nor ( n30895 , n9590 , n30727 );
and ( n30896 , n30894 , n30895 );
xor ( n30897 , n30894 , n30895 );
xor ( n30898 , n29772 , n29859 );
nor ( n30899 , n9599 , n30727 );
and ( n30900 , n30898 , n30899 );
xor ( n30901 , n30898 , n30899 );
xor ( n30902 , n29776 , n29857 );
nor ( n30903 , n9608 , n30727 );
and ( n30904 , n30902 , n30903 );
xor ( n30905 , n30902 , n30903 );
xor ( n30906 , n29780 , n29855 );
nor ( n30907 , n9617 , n30727 );
and ( n30908 , n30906 , n30907 );
xor ( n30909 , n30906 , n30907 );
xor ( n30910 , n29784 , n29853 );
nor ( n30911 , n9626 , n30727 );
and ( n30912 , n30910 , n30911 );
xor ( n30913 , n30910 , n30911 );
xor ( n30914 , n29788 , n29851 );
nor ( n30915 , n9635 , n30727 );
and ( n30916 , n30914 , n30915 );
xor ( n30917 , n30914 , n30915 );
xor ( n30918 , n29792 , n29849 );
nor ( n30919 , n9644 , n30727 );
and ( n30920 , n30918 , n30919 );
xor ( n30921 , n30918 , n30919 );
xor ( n30922 , n29796 , n29847 );
nor ( n30923 , n9653 , n30727 );
and ( n30924 , n30922 , n30923 );
xor ( n30925 , n30922 , n30923 );
xor ( n30926 , n29800 , n29845 );
nor ( n30927 , n9662 , n30727 );
and ( n30928 , n30926 , n30927 );
xor ( n30929 , n30926 , n30927 );
xor ( n30930 , n29804 , n29843 );
nor ( n30931 , n9671 , n30727 );
and ( n30932 , n30930 , n30931 );
xor ( n30933 , n30930 , n30931 );
xor ( n30934 , n29808 , n29841 );
nor ( n30935 , n9680 , n30727 );
and ( n30936 , n30934 , n30935 );
xor ( n30937 , n30934 , n30935 );
xor ( n30938 , n29812 , n29839 );
nor ( n30939 , n9689 , n30727 );
and ( n30940 , n30938 , n30939 );
xor ( n30941 , n30938 , n30939 );
xor ( n30942 , n29816 , n29837 );
nor ( n30943 , n9698 , n30727 );
and ( n30944 , n30942 , n30943 );
xor ( n30945 , n30942 , n30943 );
xor ( n30946 , n29820 , n29835 );
nor ( n30947 , n9707 , n30727 );
and ( n30948 , n30946 , n30947 );
xor ( n30949 , n30946 , n30947 );
xor ( n30950 , n29824 , n29833 );
nor ( n30951 , n9716 , n30727 );
and ( n30952 , n30950 , n30951 );
xor ( n30953 , n30950 , n30951 );
xor ( n30954 , n29828 , n29831 );
nor ( n30955 , n9725 , n30727 );
and ( n30956 , n30954 , n30955 );
xor ( n30957 , n30954 , n30955 );
xor ( n30958 , n29829 , n29830 );
nor ( n30959 , n9734 , n30727 );
and ( n30960 , n30958 , n30959 );
xor ( n30961 , n30958 , n30959 );
nor ( n30962 , n9752 , n29598 );
nor ( n30963 , n9743 , n30727 );
and ( n30964 , n30962 , n30963 );
and ( n30965 , n30961 , n30964 );
or ( n30966 , n30960 , n30965 );
and ( n30967 , n30957 , n30966 );
or ( n30968 , n30956 , n30967 );
and ( n30969 , n30953 , n30968 );
or ( n30970 , n30952 , n30969 );
and ( n30971 , n30949 , n30970 );
or ( n30972 , n30948 , n30971 );
and ( n30973 , n30945 , n30972 );
or ( n30974 , n30944 , n30973 );
and ( n30975 , n30941 , n30974 );
or ( n30976 , n30940 , n30975 );
and ( n30977 , n30937 , n30976 );
or ( n30978 , n30936 , n30977 );
and ( n30979 , n30933 , n30978 );
or ( n30980 , n30932 , n30979 );
and ( n30981 , n30929 , n30980 );
or ( n30982 , n30928 , n30981 );
and ( n30983 , n30925 , n30982 );
or ( n30984 , n30924 , n30983 );
and ( n30985 , n30921 , n30984 );
or ( n30986 , n30920 , n30985 );
and ( n30987 , n30917 , n30986 );
or ( n30988 , n30916 , n30987 );
and ( n30989 , n30913 , n30988 );
or ( n30990 , n30912 , n30989 );
and ( n30991 , n30909 , n30990 );
or ( n30992 , n30908 , n30991 );
and ( n30993 , n30905 , n30992 );
or ( n30994 , n30904 , n30993 );
and ( n30995 , n30901 , n30994 );
or ( n30996 , n30900 , n30995 );
and ( n30997 , n30897 , n30996 );
or ( n30998 , n30896 , n30997 );
and ( n30999 , n30893 , n30998 );
or ( n31000 , n30892 , n30999 );
and ( n31001 , n30889 , n31000 );
or ( n31002 , n30888 , n31001 );
and ( n31003 , n30885 , n31002 );
or ( n31004 , n30884 , n31003 );
and ( n31005 , n30881 , n31004 );
or ( n31006 , n30880 , n31005 );
and ( n31007 , n30877 , n31006 );
or ( n31008 , n30876 , n31007 );
and ( n31009 , n30873 , n31008 );
or ( n31010 , n30872 , n31009 );
and ( n31011 , n30869 , n31010 );
or ( n31012 , n30868 , n31011 );
and ( n31013 , n30865 , n31012 );
or ( n31014 , n30864 , n31013 );
and ( n31015 , n30861 , n31014 );
or ( n31016 , n30860 , n31015 );
and ( n31017 , n30857 , n31016 );
or ( n31018 , n30856 , n31017 );
and ( n31019 , n30853 , n31018 );
or ( n31020 , n30852 , n31019 );
and ( n31021 , n30849 , n31020 );
or ( n31022 , n30848 , n31021 );
and ( n31023 , n30845 , n31022 );
or ( n31024 , n30844 , n31023 );
and ( n31025 , n30841 , n31024 );
or ( n31026 , n30840 , n31025 );
and ( n31027 , n30837 , n31026 );
or ( n31028 , n30836 , n31027 );
and ( n31029 , n30833 , n31028 );
or ( n31030 , n30832 , n31029 );
and ( n31031 , n30829 , n31030 );
or ( n31032 , n30828 , n31031 );
and ( n31033 , n30825 , n31032 );
or ( n31034 , n30824 , n31033 );
and ( n31035 , n30821 , n31034 );
or ( n31036 , n30820 , n31035 );
and ( n31037 , n30817 , n31036 );
or ( n31038 , n30816 , n31037 );
and ( n31039 , n30813 , n31038 );
or ( n31040 , n30812 , n31039 );
and ( n31041 , n30809 , n31040 );
or ( n31042 , n30808 , n31041 );
and ( n31043 , n30805 , n31042 );
or ( n31044 , n30804 , n31043 );
and ( n31045 , n30801 , n31044 );
or ( n31046 , n30800 , n31045 );
and ( n31047 , n30797 , n31046 );
or ( n31048 , n30796 , n31047 );
and ( n31049 , n30793 , n31048 );
or ( n31050 , n30792 , n31049 );
and ( n31051 , n30789 , n31050 );
or ( n31052 , n30788 , n31051 );
and ( n31053 , n30785 , n31052 );
or ( n31054 , n30784 , n31053 );
and ( n31055 , n30781 , n31054 );
or ( n31056 , n30780 , n31055 );
and ( n31057 , n30777 , n31056 );
or ( n31058 , n30776 , n31057 );
and ( n31059 , n30773 , n31058 );
or ( n31060 , n30772 , n31059 );
and ( n31061 , n30769 , n31060 );
or ( n31062 , n30768 , n31061 );
and ( n31063 , n30765 , n31062 );
or ( n31064 , n30764 , n31063 );
and ( n31065 , n30761 , n31064 );
or ( n31066 , n30760 , n31065 );
and ( n31067 , n30757 , n31066 );
or ( n31068 , n30756 , n31067 );
and ( n31069 , n30753 , n31068 );
or ( n31070 , n30752 , n31069 );
and ( n31071 , n30749 , n31070 );
or ( n31072 , n30748 , n31071 );
and ( n31073 , n30745 , n31072 );
or ( n31074 , n30744 , n31073 );
and ( n31075 , n30741 , n31074 );
or ( n31076 , n30740 , n31075 );
and ( n31077 , n30737 , n31076 );
or ( n31078 , n30736 , n31077 );
and ( n31079 , n30733 , n31078 );
or ( n31080 , n30732 , n31079 );
xor ( n31081 , n30729 , n31080 );
buf ( n31082 , n473 );
not ( n31083 , n31082 );
nor ( n31084 , n601 , n31083 );
buf ( n31085 , n31084 );
nor ( n31086 , n622 , n28833 );
xor ( n31087 , n31085 , n31086 );
buf ( n31088 , n31087 );
nor ( n31089 , n646 , n27737 );
xor ( n31090 , n31088 , n31089 );
and ( n31091 , n29950 , n29951 );
buf ( n31092 , n31091 );
xor ( n31093 , n31090 , n31092 );
nor ( n31094 , n684 , n26660 );
xor ( n31095 , n31093 , n31094 );
and ( n31096 , n29953 , n29954 );
and ( n31097 , n29955 , n29957 );
or ( n31098 , n31096 , n31097 );
xor ( n31099 , n31095 , n31098 );
nor ( n31100 , n733 , n25600 );
xor ( n31101 , n31099 , n31100 );
and ( n31102 , n29958 , n29959 );
and ( n31103 , n29960 , n29963 );
or ( n31104 , n31102 , n31103 );
xor ( n31105 , n31101 , n31104 );
nor ( n31106 , n796 , n24564 );
xor ( n31107 , n31105 , n31106 );
and ( n31108 , n29964 , n29965 );
and ( n31109 , n29966 , n29969 );
or ( n31110 , n31108 , n31109 );
xor ( n31111 , n31107 , n31110 );
nor ( n31112 , n868 , n23541 );
xor ( n31113 , n31111 , n31112 );
and ( n31114 , n29970 , n29971 );
and ( n31115 , n29972 , n29975 );
or ( n31116 , n31114 , n31115 );
xor ( n31117 , n31113 , n31116 );
nor ( n31118 , n958 , n22541 );
xor ( n31119 , n31117 , n31118 );
and ( n31120 , n29976 , n29977 );
and ( n31121 , n29978 , n29981 );
or ( n31122 , n31120 , n31121 );
xor ( n31123 , n31119 , n31122 );
nor ( n31124 , n1062 , n21562 );
xor ( n31125 , n31123 , n31124 );
and ( n31126 , n29982 , n29983 );
and ( n31127 , n29984 , n29987 );
or ( n31128 , n31126 , n31127 );
xor ( n31129 , n31125 , n31128 );
nor ( n31130 , n1176 , n20601 );
xor ( n31131 , n31129 , n31130 );
and ( n31132 , n29988 , n29989 );
and ( n31133 , n29990 , n29993 );
or ( n31134 , n31132 , n31133 );
xor ( n31135 , n31131 , n31134 );
nor ( n31136 , n1303 , n19657 );
xor ( n31137 , n31135 , n31136 );
and ( n31138 , n29994 , n29995 );
and ( n31139 , n29996 , n29999 );
or ( n31140 , n31138 , n31139 );
xor ( n31141 , n31137 , n31140 );
nor ( n31142 , n1445 , n18734 );
xor ( n31143 , n31141 , n31142 );
and ( n31144 , n30000 , n30001 );
and ( n31145 , n30002 , n30005 );
or ( n31146 , n31144 , n31145 );
xor ( n31147 , n31143 , n31146 );
nor ( n31148 , n1598 , n17828 );
xor ( n31149 , n31147 , n31148 );
and ( n31150 , n30006 , n30007 );
and ( n31151 , n30008 , n30011 );
or ( n31152 , n31150 , n31151 );
xor ( n31153 , n31149 , n31152 );
nor ( n31154 , n1766 , n16943 );
xor ( n31155 , n31153 , n31154 );
and ( n31156 , n30012 , n30013 );
and ( n31157 , n30014 , n30017 );
or ( n31158 , n31156 , n31157 );
xor ( n31159 , n31155 , n31158 );
nor ( n31160 , n1945 , n16077 );
xor ( n31161 , n31159 , n31160 );
and ( n31162 , n30018 , n30019 );
and ( n31163 , n30020 , n30023 );
or ( n31164 , n31162 , n31163 );
xor ( n31165 , n31161 , n31164 );
nor ( n31166 , n2137 , n15230 );
xor ( n31167 , n31165 , n31166 );
and ( n31168 , n30024 , n30025 );
and ( n31169 , n30026 , n30029 );
or ( n31170 , n31168 , n31169 );
xor ( n31171 , n31167 , n31170 );
nor ( n31172 , n2343 , n14403 );
xor ( n31173 , n31171 , n31172 );
and ( n31174 , n30030 , n30031 );
and ( n31175 , n30032 , n30035 );
or ( n31176 , n31174 , n31175 );
xor ( n31177 , n31173 , n31176 );
nor ( n31178 , n2566 , n13599 );
xor ( n31179 , n31177 , n31178 );
and ( n31180 , n30036 , n30037 );
and ( n31181 , n30038 , n30041 );
or ( n31182 , n31180 , n31181 );
xor ( n31183 , n31179 , n31182 );
nor ( n31184 , n2797 , n12808 );
xor ( n31185 , n31183 , n31184 );
and ( n31186 , n30042 , n30043 );
and ( n31187 , n30044 , n30047 );
or ( n31188 , n31186 , n31187 );
xor ( n31189 , n31185 , n31188 );
nor ( n31190 , n3043 , n12037 );
xor ( n31191 , n31189 , n31190 );
and ( n31192 , n30048 , n30049 );
and ( n31193 , n30050 , n30053 );
or ( n31194 , n31192 , n31193 );
xor ( n31195 , n31191 , n31194 );
nor ( n31196 , n3300 , n11282 );
xor ( n31197 , n31195 , n31196 );
and ( n31198 , n30054 , n30055 );
and ( n31199 , n30056 , n30059 );
or ( n31200 , n31198 , n31199 );
xor ( n31201 , n31197 , n31200 );
nor ( n31202 , n3570 , n10547 );
xor ( n31203 , n31201 , n31202 );
and ( n31204 , n30060 , n30061 );
and ( n31205 , n30062 , n30065 );
or ( n31206 , n31204 , n31205 );
xor ( n31207 , n31203 , n31206 );
nor ( n31208 , n3853 , n9829 );
xor ( n31209 , n31207 , n31208 );
and ( n31210 , n30066 , n30067 );
and ( n31211 , n30068 , n30071 );
or ( n31212 , n31210 , n31211 );
xor ( n31213 , n31209 , n31212 );
nor ( n31214 , n4151 , n8955 );
xor ( n31215 , n31213 , n31214 );
and ( n31216 , n30072 , n30073 );
and ( n31217 , n30074 , n30077 );
or ( n31218 , n31216 , n31217 );
xor ( n31219 , n31215 , n31218 );
nor ( n31220 , n4458 , n603 );
xor ( n31221 , n31219 , n31220 );
and ( n31222 , n30078 , n30079 );
and ( n31223 , n30080 , n30083 );
or ( n31224 , n31222 , n31223 );
xor ( n31225 , n31221 , n31224 );
nor ( n31226 , n4786 , n652 );
xor ( n31227 , n31225 , n31226 );
and ( n31228 , n30084 , n30085 );
and ( n31229 , n30086 , n30089 );
or ( n31230 , n31228 , n31229 );
xor ( n31231 , n31227 , n31230 );
nor ( n31232 , n5126 , n624 );
xor ( n31233 , n31231 , n31232 );
and ( n31234 , n30090 , n30091 );
and ( n31235 , n30092 , n30095 );
or ( n31236 , n31234 , n31235 );
xor ( n31237 , n31233 , n31236 );
nor ( n31238 , n5477 , n648 );
xor ( n31239 , n31237 , n31238 );
and ( n31240 , n30096 , n30097 );
and ( n31241 , n30098 , n30101 );
or ( n31242 , n31240 , n31241 );
xor ( n31243 , n31239 , n31242 );
nor ( n31244 , n5838 , n686 );
xor ( n31245 , n31243 , n31244 );
and ( n31246 , n30102 , n30103 );
and ( n31247 , n30104 , n30107 );
or ( n31248 , n31246 , n31247 );
xor ( n31249 , n31245 , n31248 );
nor ( n31250 , n6212 , n735 );
xor ( n31251 , n31249 , n31250 );
and ( n31252 , n30108 , n30109 );
and ( n31253 , n30110 , n30113 );
or ( n31254 , n31252 , n31253 );
xor ( n31255 , n31251 , n31254 );
nor ( n31256 , n6596 , n798 );
xor ( n31257 , n31255 , n31256 );
and ( n31258 , n30114 , n30115 );
and ( n31259 , n30116 , n30119 );
or ( n31260 , n31258 , n31259 );
xor ( n31261 , n31257 , n31260 );
nor ( n31262 , n6997 , n870 );
xor ( n31263 , n31261 , n31262 );
and ( n31264 , n30120 , n30121 );
and ( n31265 , n30122 , n30125 );
or ( n31266 , n31264 , n31265 );
xor ( n31267 , n31263 , n31266 );
nor ( n31268 , n7413 , n960 );
xor ( n31269 , n31267 , n31268 );
and ( n31270 , n30126 , n30127 );
and ( n31271 , n30128 , n30131 );
or ( n31272 , n31270 , n31271 );
xor ( n31273 , n31269 , n31272 );
nor ( n31274 , n7841 , n1064 );
xor ( n31275 , n31273 , n31274 );
and ( n31276 , n30132 , n30133 );
and ( n31277 , n30134 , n30137 );
or ( n31278 , n31276 , n31277 );
xor ( n31279 , n31275 , n31278 );
nor ( n31280 , n8281 , n1178 );
xor ( n31281 , n31279 , n31280 );
and ( n31282 , n30138 , n30139 );
and ( n31283 , n30140 , n30143 );
or ( n31284 , n31282 , n31283 );
xor ( n31285 , n31281 , n31284 );
nor ( n31286 , n8737 , n1305 );
xor ( n31287 , n31285 , n31286 );
and ( n31288 , n30144 , n30145 );
and ( n31289 , n30146 , n30149 );
or ( n31290 , n31288 , n31289 );
xor ( n31291 , n31287 , n31290 );
nor ( n31292 , n9420 , n1447 );
xor ( n31293 , n31291 , n31292 );
and ( n31294 , n30150 , n30151 );
and ( n31295 , n30152 , n30155 );
or ( n31296 , n31294 , n31295 );
xor ( n31297 , n31293 , n31296 );
nor ( n31298 , n10312 , n1600 );
xor ( n31299 , n31297 , n31298 );
and ( n31300 , n30156 , n30157 );
and ( n31301 , n30158 , n30161 );
or ( n31302 , n31300 , n31301 );
xor ( n31303 , n31299 , n31302 );
nor ( n31304 , n11041 , n1768 );
xor ( n31305 , n31303 , n31304 );
and ( n31306 , n30162 , n30163 );
and ( n31307 , n30164 , n30167 );
or ( n31308 , n31306 , n31307 );
xor ( n31309 , n31305 , n31308 );
nor ( n31310 , n11790 , n1947 );
xor ( n31311 , n31309 , n31310 );
and ( n31312 , n30168 , n30169 );
and ( n31313 , n30170 , n30173 );
or ( n31314 , n31312 , n31313 );
xor ( n31315 , n31311 , n31314 );
nor ( n31316 , n12555 , n2139 );
xor ( n31317 , n31315 , n31316 );
and ( n31318 , n30174 , n30175 );
and ( n31319 , n30176 , n30179 );
or ( n31320 , n31318 , n31319 );
xor ( n31321 , n31317 , n31320 );
nor ( n31322 , n13340 , n2345 );
xor ( n31323 , n31321 , n31322 );
and ( n31324 , n30180 , n30181 );
and ( n31325 , n30182 , n30185 );
or ( n31326 , n31324 , n31325 );
xor ( n31327 , n31323 , n31326 );
nor ( n31328 , n14138 , n2568 );
xor ( n31329 , n31327 , n31328 );
and ( n31330 , n30186 , n30187 );
and ( n31331 , n30188 , n30191 );
or ( n31332 , n31330 , n31331 );
xor ( n31333 , n31329 , n31332 );
nor ( n31334 , n14959 , n2799 );
xor ( n31335 , n31333 , n31334 );
and ( n31336 , n30192 , n30193 );
and ( n31337 , n30194 , n30197 );
or ( n31338 , n31336 , n31337 );
xor ( n31339 , n31335 , n31338 );
nor ( n31340 , n15800 , n3045 );
xor ( n31341 , n31339 , n31340 );
and ( n31342 , n30198 , n30199 );
and ( n31343 , n30200 , n30203 );
or ( n31344 , n31342 , n31343 );
xor ( n31345 , n31341 , n31344 );
nor ( n31346 , n16660 , n3302 );
xor ( n31347 , n31345 , n31346 );
and ( n31348 , n30204 , n30205 );
and ( n31349 , n30206 , n30209 );
or ( n31350 , n31348 , n31349 );
xor ( n31351 , n31347 , n31350 );
nor ( n31352 , n17539 , n3572 );
xor ( n31353 , n31351 , n31352 );
and ( n31354 , n30210 , n30211 );
and ( n31355 , n30212 , n30215 );
or ( n31356 , n31354 , n31355 );
xor ( n31357 , n31353 , n31356 );
nor ( n31358 , n18439 , n3855 );
xor ( n31359 , n31357 , n31358 );
and ( n31360 , n30216 , n30217 );
and ( n31361 , n30218 , n30221 );
or ( n31362 , n31360 , n31361 );
xor ( n31363 , n31359 , n31362 );
nor ( n31364 , n19356 , n4153 );
xor ( n31365 , n31363 , n31364 );
and ( n31366 , n30222 , n30223 );
and ( n31367 , n30224 , n30227 );
or ( n31368 , n31366 , n31367 );
xor ( n31369 , n31365 , n31368 );
nor ( n31370 , n20294 , n4460 );
xor ( n31371 , n31369 , n31370 );
and ( n31372 , n30228 , n30229 );
and ( n31373 , n30230 , n30233 );
or ( n31374 , n31372 , n31373 );
xor ( n31375 , n31371 , n31374 );
nor ( n31376 , n21249 , n4788 );
xor ( n31377 , n31375 , n31376 );
and ( n31378 , n30234 , n30235 );
and ( n31379 , n30236 , n30239 );
or ( n31380 , n31378 , n31379 );
xor ( n31381 , n31377 , n31380 );
nor ( n31382 , n22222 , n5128 );
xor ( n31383 , n31381 , n31382 );
and ( n31384 , n30240 , n30241 );
and ( n31385 , n30242 , n30245 );
or ( n31386 , n31384 , n31385 );
xor ( n31387 , n31383 , n31386 );
nor ( n31388 , n23216 , n5479 );
xor ( n31389 , n31387 , n31388 );
and ( n31390 , n30246 , n30247 );
and ( n31391 , n30248 , n30251 );
or ( n31392 , n31390 , n31391 );
xor ( n31393 , n31389 , n31392 );
nor ( n31394 , n24233 , n5840 );
xor ( n31395 , n31393 , n31394 );
and ( n31396 , n30252 , n30253 );
and ( n31397 , n30254 , n30257 );
or ( n31398 , n31396 , n31397 );
xor ( n31399 , n31395 , n31398 );
nor ( n31400 , n25263 , n6214 );
xor ( n31401 , n31399 , n31400 );
and ( n31402 , n30258 , n30259 );
and ( n31403 , n30260 , n30263 );
or ( n31404 , n31402 , n31403 );
xor ( n31405 , n31401 , n31404 );
nor ( n31406 , n26317 , n6598 );
xor ( n31407 , n31405 , n31406 );
and ( n31408 , n30264 , n30265 );
and ( n31409 , n30266 , n30269 );
or ( n31410 , n31408 , n31409 );
xor ( n31411 , n31407 , n31410 );
nor ( n31412 , n27388 , n6999 );
xor ( n31413 , n31411 , n31412 );
and ( n31414 , n30270 , n30271 );
and ( n31415 , n30272 , n30275 );
or ( n31416 , n31414 , n31415 );
xor ( n31417 , n31413 , n31416 );
nor ( n31418 , n28478 , n7415 );
xor ( n31419 , n31417 , n31418 );
and ( n31420 , n30276 , n30277 );
and ( n31421 , n30278 , n30281 );
or ( n31422 , n31420 , n31421 );
xor ( n31423 , n31419 , n31422 );
nor ( n31424 , n29587 , n7843 );
xor ( n31425 , n31423 , n31424 );
and ( n31426 , n30282 , n30283 );
and ( n31427 , n30284 , n30287 );
or ( n31428 , n31426 , n31427 );
xor ( n31429 , n31425 , n31428 );
nor ( n31430 , n30716 , n8283 );
xor ( n31431 , n31429 , n31430 );
and ( n31432 , n30288 , n30289 );
and ( n31433 , n30290 , n30293 );
or ( n31434 , n31432 , n31433 );
xor ( n31435 , n31431 , n31434 );
and ( n31436 , n30645 , n30646 );
and ( n31437 , n30646 , n30701 );
and ( n31438 , n30645 , n30701 );
or ( n31439 , n31436 , n31437 , n31438 );
and ( n31440 , n30307 , n30640 );
and ( n31441 , n30640 , n30702 );
and ( n31442 , n30307 , n30702 );
or ( n31443 , n31440 , n31441 , n31442 );
xor ( n31444 , n31439 , n31443 );
and ( n31445 , n30311 , n30431 );
and ( n31446 , n30431 , n30639 );
and ( n31447 , n30311 , n30639 );
or ( n31448 , n31445 , n31446 , n31447 );
and ( n31449 , n30436 , n30514 );
and ( n31450 , n30514 , n30638 );
and ( n31451 , n30436 , n30638 );
or ( n31452 , n31449 , n31450 , n31451 );
and ( n31453 , n30324 , n30392 );
and ( n31454 , n30392 , n30429 );
and ( n31455 , n30324 , n30429 );
or ( n31456 , n31453 , n31454 , n31455 );
and ( n31457 , n30440 , n30444 );
and ( n31458 , n30444 , n30513 );
and ( n31459 , n30440 , n30513 );
or ( n31460 , n31457 , n31458 , n31459 );
xor ( n31461 , n31456 , n31460 );
and ( n31462 , n30397 , n30401 );
and ( n31463 , n30401 , n30428 );
and ( n31464 , n30397 , n30428 );
or ( n31465 , n31462 , n31463 , n31464 );
and ( n31466 , n30406 , n30410 );
and ( n31467 , n30410 , n30427 );
and ( n31468 , n30406 , n30427 );
or ( n31469 , n31466 , n31467 , n31468 );
and ( n31470 , n30453 , n30468 );
and ( n31471 , n30468 , n30485 );
and ( n31472 , n30453 , n30485 );
or ( n31473 , n31470 , n31471 , n31472 );
xor ( n31474 , n31469 , n31473 );
and ( n31475 , n30415 , n30420 );
and ( n31476 , n30420 , n30426 );
and ( n31477 , n30415 , n30426 );
or ( n31478 , n31475 , n31476 , n31477 );
and ( n31479 , n30457 , n30461 );
and ( n31480 , n30461 , n30467 );
and ( n31481 , n30457 , n30467 );
or ( n31482 , n31479 , n31480 , n31481 );
xor ( n31483 , n31478 , n31482 );
and ( n31484 , n30422 , n30423 );
and ( n31485 , n30423 , n30425 );
and ( n31486 , n30422 , n30425 );
or ( n31487 , n31484 , n31485 , n31486 );
and ( n31488 , n11015 , n3495 );
and ( n31489 , n11769 , n3271 );
xor ( n31490 , n31488 , n31489 );
and ( n31491 , n12320 , n2981 );
xor ( n31492 , n31490 , n31491 );
xor ( n31493 , n31487 , n31492 );
and ( n31494 , n8718 , n4403 );
and ( n31495 , n9400 , n4102 );
xor ( n31496 , n31494 , n31495 );
and ( n31497 , n10291 , n3749 );
xor ( n31498 , n31496 , n31497 );
xor ( n31499 , n31493 , n31498 );
xor ( n31500 , n31483 , n31499 );
xor ( n31501 , n31474 , n31500 );
xor ( n31502 , n31465 , n31501 );
and ( n31503 , n30358 , n30374 );
and ( n31504 , n30374 , n30390 );
and ( n31505 , n30358 , n30390 );
or ( n31506 , n31503 , n31504 , n31505 );
and ( n31507 , n30379 , n30383 );
and ( n31508 , n30383 , n30389 );
and ( n31509 , n30379 , n30389 );
or ( n31510 , n31507 , n31508 , n31509 );
and ( n31511 , n30369 , n30370 );
and ( n31512 , n30370 , n30372 );
and ( n31513 , n30369 , n30372 );
or ( n31514 , n31511 , n31512 , n31513 );
and ( n31515 , n18144 , n1551 );
and ( n31516 , n19324 , n1424 );
xor ( n31517 , n31515 , n31516 );
and ( n31518 , n20233 , n1254 );
xor ( n31519 , n31517 , n31518 );
xor ( n31520 , n31514 , n31519 );
and ( n31521 , n15758 , n2100 );
and ( n31522 , n16637 , n1882 );
xor ( n31523 , n31521 , n31522 );
and ( n31524 , n17512 , n1738 );
xor ( n31525 , n31523 , n31524 );
xor ( n31526 , n31520 , n31525 );
xor ( n31527 , n31510 , n31526 );
and ( n31528 , n30385 , n30386 );
and ( n31529 , n30386 , n30388 );
and ( n31530 , n30385 , n30388 );
or ( n31531 , n31528 , n31529 , n31530 );
and ( n31532 , n30416 , n30417 );
and ( n31533 , n30417 , n30419 );
and ( n31534 , n30416 , n30419 );
or ( n31535 , n31532 , n31533 , n31534 );
xor ( n31536 , n31531 , n31535 );
and ( n31537 , n13322 , n2739 );
and ( n31538 , n14118 , n2544 );
xor ( n31539 , n31537 , n31538 );
and ( n31540 , n14938 , n2298 );
xor ( n31541 , n31539 , n31540 );
xor ( n31542 , n31536 , n31541 );
xor ( n31543 , n31527 , n31542 );
xor ( n31544 , n31506 , n31543 );
and ( n31545 , n30341 , n30345 );
and ( n31546 , n30345 , n30351 );
and ( n31547 , n30341 , n30351 );
or ( n31548 , n31545 , n31546 , n31547 );
and ( n31549 , n30362 , n30367 );
and ( n31550 , n30367 , n30373 );
and ( n31551 , n30362 , n30373 );
or ( n31552 , n31549 , n31550 , n31551 );
xor ( n31553 , n31548 , n31552 );
and ( n31554 , n30347 , n30348 );
and ( n31555 , n30348 , n30350 );
and ( n31556 , n30347 , n30350 );
or ( n31557 , n31554 , n31555 , n31556 );
and ( n31558 , n30363 , n30364 );
and ( n31559 , n30364 , n30366 );
and ( n31560 , n30363 , n30366 );
or ( n31561 , n31558 , n31559 , n31560 );
xor ( n31562 , n31557 , n31561 );
and ( n31563 , n21216 , n1134 );
and ( n31564 , n22186 , n1034 );
xor ( n31565 , n31563 , n31564 );
and ( n31566 , n22892 , n940 );
xor ( n31567 , n31565 , n31566 );
xor ( n31568 , n31562 , n31567 );
xor ( n31569 , n31553 , n31568 );
xor ( n31570 , n31544 , n31569 );
xor ( n31571 , n31502 , n31570 );
xor ( n31572 , n31461 , n31571 );
xor ( n31573 , n31452 , n31572 );
and ( n31574 , n30519 , n30566 );
and ( n31575 , n30566 , n30637 );
and ( n31576 , n30519 , n30637 );
or ( n31577 , n31574 , n31575 , n31576 );
and ( n31578 , n30449 , n30486 );
and ( n31579 , n30486 , n30512 );
and ( n31580 , n30449 , n30512 );
or ( n31581 , n31578 , n31579 , n31580 );
and ( n31582 , n30523 , n30527 );
and ( n31583 , n30527 , n30565 );
and ( n31584 , n30523 , n30565 );
or ( n31585 , n31582 , n31583 , n31584 );
xor ( n31586 , n31581 , n31585 );
and ( n31587 , n30491 , n30495 );
and ( n31588 , n30495 , n30511 );
and ( n31589 , n30491 , n30511 );
or ( n31590 , n31587 , n31588 , n31589 );
and ( n31591 , n30473 , n30478 );
and ( n31592 , n30478 , n30484 );
and ( n31593 , n30473 , n30484 );
or ( n31594 , n31591 , n31592 , n31593 );
and ( n31595 , n30463 , n30464 );
and ( n31596 , n30464 , n30466 );
and ( n31597 , n30463 , n30466 );
or ( n31598 , n31595 , n31596 , n31597 );
and ( n31599 , n30474 , n30475 );
and ( n31600 , n30475 , n30477 );
and ( n31601 , n30474 , n30477 );
or ( n31602 , n31599 , n31600 , n31601 );
xor ( n31603 , n31598 , n31602 );
and ( n31604 , n7385 , n5408 );
and ( n31605 , n7808 , n5103 );
xor ( n31606 , n31604 , n31605 );
and ( n31607 , n8079 , n4730 );
xor ( n31608 , n31606 , n31607 );
xor ( n31609 , n31603 , n31608 );
xor ( n31610 , n31594 , n31609 );
and ( n31611 , n30480 , n30481 );
and ( n31612 , n30481 , n30483 );
and ( n31613 , n30480 , n30483 );
or ( n31614 , n31611 , n31612 , n31613 );
and ( n31615 , n6816 , n5765 );
buf ( n31616 , n31615 );
xor ( n31617 , n31614 , n31616 );
and ( n31618 , n4959 , n7662 );
and ( n31619 , n5459 , n7310 );
xor ( n31620 , n31618 , n31619 );
and ( n31621 , n5819 , n6971 );
xor ( n31622 , n31620 , n31621 );
xor ( n31623 , n31617 , n31622 );
xor ( n31624 , n31610 , n31623 );
xor ( n31625 , n31590 , n31624 );
and ( n31626 , n30500 , n30504 );
and ( n31627 , n30504 , n30510 );
and ( n31628 , n30500 , n30510 );
or ( n31629 , n31626 , n31627 , n31628 );
and ( n31630 , n30536 , n30541 );
and ( n31631 , n30541 , n30547 );
and ( n31632 , n30536 , n30547 );
or ( n31633 , n31630 , n31631 , n31632 );
xor ( n31634 , n31629 , n31633 );
and ( n31635 , n30506 , n30507 );
and ( n31636 , n30507 , n30509 );
and ( n31637 , n30506 , n30509 );
or ( n31638 , n31635 , n31636 , n31637 );
and ( n31639 , n30537 , n30538 );
and ( n31640 , n30538 , n30540 );
and ( n31641 , n30537 , n30540 );
or ( n31642 , n31639 , n31640 , n31641 );
xor ( n31643 , n31638 , n31642 );
and ( n31644 , n4132 , n9348 );
and ( n31645 , n4438 , n8669 );
xor ( n31646 , n31644 , n31645 );
and ( n31647 , n4766 , n8243 );
xor ( n31648 , n31646 , n31647 );
xor ( n31649 , n31643 , n31648 );
xor ( n31650 , n31634 , n31649 );
xor ( n31651 , n31625 , n31650 );
xor ( n31652 , n31586 , n31651 );
xor ( n31653 , n31577 , n31652 );
and ( n31654 , n30571 , n30597 );
and ( n31655 , n30597 , n30636 );
and ( n31656 , n30571 , n30636 );
or ( n31657 , n31654 , n31655 , n31656 );
and ( n31658 , n30532 , n30548 );
and ( n31659 , n30548 , n30564 );
and ( n31660 , n30532 , n30564 );
or ( n31661 , n31658 , n31659 , n31660 );
and ( n31662 , n30575 , n30579 );
and ( n31663 , n30579 , n30596 );
and ( n31664 , n30575 , n30596 );
or ( n31665 , n31662 , n31663 , n31664 );
xor ( n31666 , n31661 , n31665 );
and ( n31667 , n30553 , n30557 );
and ( n31668 , n30557 , n30563 );
and ( n31669 , n30553 , n30563 );
or ( n31670 , n31667 , n31668 , n31669 );
and ( n31671 , n30543 , n30544 );
and ( n31672 , n30544 , n30546 );
and ( n31673 , n30543 , n30546 );
or ( n31674 , n31671 , n31672 , n31673 );
and ( n31675 , n3182 , n11718 );
and ( n31676 , n3545 , n10977 );
xor ( n31677 , n31675 , n31676 );
and ( n31678 , n3801 , n10239 );
xor ( n31679 , n31677 , n31678 );
xor ( n31680 , n31674 , n31679 );
and ( n31681 , n2462 , n14044 );
and ( n31682 , n2779 , n13256 );
xor ( n31683 , n31681 , n31682 );
and ( n31684 , n3024 , n12531 );
xor ( n31685 , n31683 , n31684 );
xor ( n31686 , n31680 , n31685 );
xor ( n31687 , n31670 , n31686 );
and ( n31688 , n30559 , n30560 );
and ( n31689 , n30560 , n30562 );
and ( n31690 , n30559 , n30562 );
or ( n31691 , n31688 , n31689 , n31690 );
and ( n31692 , n30585 , n30586 );
and ( n31693 , n30586 , n30588 );
and ( n31694 , n30585 , n30588 );
or ( n31695 , n31692 , n31693 , n31694 );
xor ( n31696 , n31691 , n31695 );
and ( n31697 , n1933 , n16550 );
and ( n31698 , n2120 , n15691 );
xor ( n31699 , n31697 , n31698 );
and ( n31700 , n2324 , n14838 );
xor ( n31701 , n31699 , n31700 );
xor ( n31702 , n31696 , n31701 );
xor ( n31703 , n31687 , n31702 );
xor ( n31704 , n31666 , n31703 );
xor ( n31705 , n31657 , n31704 );
and ( n31706 , n30602 , n30617 );
and ( n31707 , n30617 , n30635 );
and ( n31708 , n30602 , n30635 );
or ( n31709 , n31706 , n31707 , n31708 );
and ( n31710 , n30584 , n30589 );
and ( n31711 , n30589 , n30595 );
and ( n31712 , n30584 , n30595 );
or ( n31713 , n31710 , n31711 , n31712 );
and ( n31714 , n30606 , n30610 );
and ( n31715 , n30610 , n30616 );
and ( n31716 , n30606 , n30616 );
or ( n31717 , n31714 , n31715 , n31716 );
xor ( n31718 , n31713 , n31717 );
and ( n31719 , n30591 , n30592 );
and ( n31720 , n30592 , n30594 );
and ( n31721 , n30591 , n30594 );
or ( n31722 , n31719 , n31720 , n31721 );
and ( n31723 , n1383 , n19222 );
and ( n31724 , n1580 , n18407 );
xor ( n31725 , n31723 , n31724 );
and ( n31726 , n1694 , n17422 );
xor ( n31727 , n31725 , n31726 );
xor ( n31728 , n31722 , n31727 );
and ( n31729 , n1047 , n22065 );
and ( n31730 , n1164 , n20976 );
xor ( n31731 , n31729 , n31730 );
and ( n31732 , n1287 , n20156 );
xor ( n31733 , n31731 , n31732 );
xor ( n31734 , n31728 , n31733 );
xor ( n31735 , n31718 , n31734 );
xor ( n31736 , n31709 , n31735 );
and ( n31737 , n30622 , n30627 );
and ( n31738 , n30627 , n30634 );
and ( n31739 , n30622 , n30634 );
or ( n31740 , n31737 , n31738 , n31739 );
and ( n31741 , n30612 , n30613 );
and ( n31742 , n30613 , n30615 );
and ( n31743 , n30612 , n30615 );
or ( n31744 , n31741 , n31742 , n31743 );
and ( n31745 , n30623 , n30624 );
and ( n31746 , n30624 , n30626 );
and ( n31747 , n30623 , n30626 );
or ( n31748 , n31745 , n31746 , n31747 );
xor ( n31749 , n31744 , n31748 );
and ( n31750 , n783 , n25163 );
and ( n31751 , n856 , n24137 );
xor ( n31752 , n31750 , n31751 );
and ( n31753 , n925 , n23075 );
xor ( n31754 , n31752 , n31753 );
xor ( n31755 , n31749 , n31754 );
xor ( n31756 , n31740 , n31755 );
and ( n31757 , n30630 , n30631 );
and ( n31758 , n30631 , n30633 );
and ( n31759 , n30630 , n30633 );
or ( n31760 , n31757 , n31758 , n31759 );
buf ( n31761 , n409 );
and ( n31762 , n599 , n31761 );
and ( n31763 , n608 , n30629 );
xor ( n31764 , n31762 , n31763 );
and ( n31765 , n611 , n29508 );
xor ( n31766 , n31764 , n31765 );
xor ( n31767 , n31760 , n31766 );
and ( n31768 , n632 , n28406 );
and ( n31769 , n671 , n27296 );
xor ( n31770 , n31768 , n31769 );
and ( n31771 , n715 , n26216 );
xor ( n31772 , n31770 , n31771 );
xor ( n31773 , n31767 , n31772 );
xor ( n31774 , n31756 , n31773 );
xor ( n31775 , n31736 , n31774 );
xor ( n31776 , n31705 , n31775 );
xor ( n31777 , n31653 , n31776 );
xor ( n31778 , n31573 , n31777 );
xor ( n31779 , n31448 , n31778 );
and ( n31780 , n30315 , n30319 );
and ( n31781 , n30319 , n30430 );
and ( n31782 , n30315 , n30430 );
or ( n31783 , n31780 , n31781 , n31782 );
and ( n31784 , n30651 , n30700 );
xor ( n31785 , n31783 , n31784 );
and ( n31786 , n30694 , n30696 );
and ( n31787 , n30655 , n30659 );
and ( n31788 , n30659 , n30699 );
and ( n31789 , n30655 , n30699 );
or ( n31790 , n31787 , n31788 , n31789 );
xor ( n31791 , n31786 , n31790 );
and ( n31792 , n30328 , n30353 );
and ( n31793 , n30353 , n30391 );
and ( n31794 , n30328 , n30391 );
or ( n31795 , n31792 , n31793 , n31794 );
and ( n31796 , n30664 , n30668 );
and ( n31797 , n30668 , n30698 );
and ( n31798 , n30664 , n30698 );
or ( n31799 , n31796 , n31797 , n31798 );
xor ( n31800 , n31795 , n31799 );
and ( n31801 , n30332 , n30336 );
and ( n31802 , n30336 , n30352 );
and ( n31803 , n30332 , n30352 );
or ( n31804 , n31801 , n31802 , n31803 );
and ( n31805 , n30673 , n30689 );
and ( n31806 , n30689 , n30697 );
and ( n31807 , n30673 , n30697 );
or ( n31808 , n31805 , n31806 , n31807 );
xor ( n31809 , n31804 , n31808 );
and ( n31810 , n30677 , n30682 );
and ( n31811 , n30682 , n30688 );
and ( n31812 , n30677 , n30688 );
or ( n31813 , n31810 , n31811 , n31812 );
and ( n31814 , n30684 , n30685 );
and ( n31815 , n30685 , n30687 );
and ( n31816 , n30684 , n30687 );
or ( n31817 , n31814 , n31815 , n31816 );
and ( n31818 , n27361 , n663 );
and ( n31819 , n28456 , n635 );
xor ( n31820 , n31818 , n31819 );
and ( n31821 , n29559 , n606 );
xor ( n31822 , n31820 , n31821 );
xor ( n31823 , n31817 , n31822 );
and ( n31824 , n24214 , n840 );
and ( n31825 , n25243 , n771 );
xor ( n31826 , n31824 , n31825 );
and ( n31827 , n26296 , n719 );
xor ( n31828 , n31826 , n31827 );
xor ( n31829 , n31823 , n31828 );
xor ( n31830 , n31813 , n31829 );
and ( n31831 , n30678 , n30679 );
and ( n31832 , n30679 , n30681 );
and ( n31833 , n30678 , n30681 );
or ( n31834 , n31831 , n31832 , n31833 );
and ( n31835 , n30695 , n615 );
buf ( n31836 , n409 );
and ( n31837 , n31836 , n612 );
xor ( n31838 , n31835 , n31837 );
xor ( n31839 , n31834 , n31838 );
xor ( n31840 , n31830 , n31839 );
xor ( n31841 , n31809 , n31840 );
xor ( n31842 , n31800 , n31841 );
xor ( n31843 , n31791 , n31842 );
xor ( n31844 , n31785 , n31843 );
xor ( n31845 , n31779 , n31844 );
xor ( n31846 , n31444 , n31845 );
and ( n31847 , n30298 , n30302 );
and ( n31848 , n30302 , n30703 );
and ( n31849 , n30298 , n30703 );
or ( n31850 , n31847 , n31848 , n31849 );
xor ( n31851 , n31846 , n31850 );
and ( n31852 , n30704 , n30708 );
and ( n31853 , n30709 , n30712 );
or ( n31854 , n31852 , n31853 );
xor ( n31855 , n31851 , n31854 );
buf ( n31856 , n31855 );
buf ( n31857 , n31856 );
not ( n31858 , n31857 );
nor ( n31859 , n31858 , n8739 );
xor ( n31860 , n31435 , n31859 );
and ( n31861 , n30294 , n30717 );
and ( n31862 , n30718 , n30721 );
or ( n31863 , n31861 , n31862 );
xor ( n31864 , n31860 , n31863 );
buf ( n31865 , n31864 );
buf ( n31866 , n31865 );
not ( n31867 , n31866 );
buf ( n31868 , n560 );
not ( n31869 , n31868 );
nor ( n31870 , n31867 , n31869 );
xor ( n31871 , n31081 , n31870 );
xor ( n31872 , n30733 , n31078 );
nor ( n31873 , n30725 , n31869 );
and ( n31874 , n31872 , n31873 );
xor ( n31875 , n31872 , n31873 );
xor ( n31876 , n30737 , n31076 );
nor ( n31877 , n29596 , n31869 );
and ( n31878 , n31876 , n31877 );
xor ( n31879 , n31876 , n31877 );
xor ( n31880 , n30741 , n31074 );
nor ( n31881 , n28487 , n31869 );
and ( n31882 , n31880 , n31881 );
xor ( n31883 , n31880 , n31881 );
xor ( n31884 , n30745 , n31072 );
nor ( n31885 , n27397 , n31869 );
and ( n31886 , n31884 , n31885 );
xor ( n31887 , n31884 , n31885 );
xor ( n31888 , n30749 , n31070 );
nor ( n31889 , n26326 , n31869 );
and ( n31890 , n31888 , n31889 );
xor ( n31891 , n31888 , n31889 );
xor ( n31892 , n30753 , n31068 );
nor ( n31893 , n25272 , n31869 );
and ( n31894 , n31892 , n31893 );
xor ( n31895 , n31892 , n31893 );
xor ( n31896 , n30757 , n31066 );
nor ( n31897 , n24242 , n31869 );
and ( n31898 , n31896 , n31897 );
xor ( n31899 , n31896 , n31897 );
xor ( n31900 , n30761 , n31064 );
nor ( n31901 , n23225 , n31869 );
and ( n31902 , n31900 , n31901 );
xor ( n31903 , n31900 , n31901 );
xor ( n31904 , n30765 , n31062 );
nor ( n31905 , n22231 , n31869 );
and ( n31906 , n31904 , n31905 );
xor ( n31907 , n31904 , n31905 );
xor ( n31908 , n30769 , n31060 );
nor ( n31909 , n21258 , n31869 );
and ( n31910 , n31908 , n31909 );
xor ( n31911 , n31908 , n31909 );
xor ( n31912 , n30773 , n31058 );
nor ( n31913 , n20303 , n31869 );
and ( n31914 , n31912 , n31913 );
xor ( n31915 , n31912 , n31913 );
xor ( n31916 , n30777 , n31056 );
nor ( n31917 , n19365 , n31869 );
and ( n31918 , n31916 , n31917 );
xor ( n31919 , n31916 , n31917 );
xor ( n31920 , n30781 , n31054 );
nor ( n31921 , n18448 , n31869 );
and ( n31922 , n31920 , n31921 );
xor ( n31923 , n31920 , n31921 );
xor ( n31924 , n30785 , n31052 );
nor ( n31925 , n17548 , n31869 );
and ( n31926 , n31924 , n31925 );
xor ( n31927 , n31924 , n31925 );
xor ( n31928 , n30789 , n31050 );
nor ( n31929 , n16669 , n31869 );
and ( n31930 , n31928 , n31929 );
xor ( n31931 , n31928 , n31929 );
xor ( n31932 , n30793 , n31048 );
nor ( n31933 , n15809 , n31869 );
and ( n31934 , n31932 , n31933 );
xor ( n31935 , n31932 , n31933 );
xor ( n31936 , n30797 , n31046 );
nor ( n31937 , n14968 , n31869 );
and ( n31938 , n31936 , n31937 );
xor ( n31939 , n31936 , n31937 );
xor ( n31940 , n30801 , n31044 );
nor ( n31941 , n14147 , n31869 );
and ( n31942 , n31940 , n31941 );
xor ( n31943 , n31940 , n31941 );
xor ( n31944 , n30805 , n31042 );
nor ( n31945 , n13349 , n31869 );
and ( n31946 , n31944 , n31945 );
xor ( n31947 , n31944 , n31945 );
xor ( n31948 , n30809 , n31040 );
nor ( n31949 , n12564 , n31869 );
and ( n31950 , n31948 , n31949 );
xor ( n31951 , n31948 , n31949 );
xor ( n31952 , n30813 , n31038 );
nor ( n31953 , n11799 , n31869 );
and ( n31954 , n31952 , n31953 );
xor ( n31955 , n31952 , n31953 );
xor ( n31956 , n30817 , n31036 );
nor ( n31957 , n11050 , n31869 );
and ( n31958 , n31956 , n31957 );
xor ( n31959 , n31956 , n31957 );
xor ( n31960 , n30821 , n31034 );
nor ( n31961 , n10321 , n31869 );
and ( n31962 , n31960 , n31961 );
xor ( n31963 , n31960 , n31961 );
xor ( n31964 , n30825 , n31032 );
nor ( n31965 , n9429 , n31869 );
and ( n31966 , n31964 , n31965 );
xor ( n31967 , n31964 , n31965 );
xor ( n31968 , n30829 , n31030 );
nor ( n31969 , n8949 , n31869 );
and ( n31970 , n31968 , n31969 );
xor ( n31971 , n31968 , n31969 );
xor ( n31972 , n30833 , n31028 );
nor ( n31973 , n9437 , n31869 );
and ( n31974 , n31972 , n31973 );
xor ( n31975 , n31972 , n31973 );
xor ( n31976 , n30837 , n31026 );
nor ( n31977 , n9446 , n31869 );
and ( n31978 , n31976 , n31977 );
xor ( n31979 , n31976 , n31977 );
xor ( n31980 , n30841 , n31024 );
nor ( n31981 , n9455 , n31869 );
and ( n31982 , n31980 , n31981 );
xor ( n31983 , n31980 , n31981 );
xor ( n31984 , n30845 , n31022 );
nor ( n31985 , n9464 , n31869 );
and ( n31986 , n31984 , n31985 );
xor ( n31987 , n31984 , n31985 );
xor ( n31988 , n30849 , n31020 );
nor ( n31989 , n9473 , n31869 );
and ( n31990 , n31988 , n31989 );
xor ( n31991 , n31988 , n31989 );
xor ( n31992 , n30853 , n31018 );
nor ( n31993 , n9482 , n31869 );
and ( n31994 , n31992 , n31993 );
xor ( n31995 , n31992 , n31993 );
xor ( n31996 , n30857 , n31016 );
nor ( n31997 , n9491 , n31869 );
and ( n31998 , n31996 , n31997 );
xor ( n31999 , n31996 , n31997 );
xor ( n32000 , n30861 , n31014 );
nor ( n32001 , n9500 , n31869 );
and ( n32002 , n32000 , n32001 );
xor ( n32003 , n32000 , n32001 );
xor ( n32004 , n30865 , n31012 );
nor ( n32005 , n9509 , n31869 );
and ( n32006 , n32004 , n32005 );
xor ( n32007 , n32004 , n32005 );
xor ( n32008 , n30869 , n31010 );
nor ( n32009 , n9518 , n31869 );
and ( n32010 , n32008 , n32009 );
xor ( n32011 , n32008 , n32009 );
xor ( n32012 , n30873 , n31008 );
nor ( n32013 , n9527 , n31869 );
and ( n32014 , n32012 , n32013 );
xor ( n32015 , n32012 , n32013 );
xor ( n32016 , n30877 , n31006 );
nor ( n32017 , n9536 , n31869 );
and ( n32018 , n32016 , n32017 );
xor ( n32019 , n32016 , n32017 );
xor ( n32020 , n30881 , n31004 );
nor ( n32021 , n9545 , n31869 );
and ( n32022 , n32020 , n32021 );
xor ( n32023 , n32020 , n32021 );
xor ( n32024 , n30885 , n31002 );
nor ( n32025 , n9554 , n31869 );
and ( n32026 , n32024 , n32025 );
xor ( n32027 , n32024 , n32025 );
xor ( n32028 , n30889 , n31000 );
nor ( n32029 , n9563 , n31869 );
and ( n32030 , n32028 , n32029 );
xor ( n32031 , n32028 , n32029 );
xor ( n32032 , n30893 , n30998 );
nor ( n32033 , n9572 , n31869 );
and ( n32034 , n32032 , n32033 );
xor ( n32035 , n32032 , n32033 );
xor ( n32036 , n30897 , n30996 );
nor ( n32037 , n9581 , n31869 );
and ( n32038 , n32036 , n32037 );
xor ( n32039 , n32036 , n32037 );
xor ( n32040 , n30901 , n30994 );
nor ( n32041 , n9590 , n31869 );
and ( n32042 , n32040 , n32041 );
xor ( n32043 , n32040 , n32041 );
xor ( n32044 , n30905 , n30992 );
nor ( n32045 , n9599 , n31869 );
and ( n32046 , n32044 , n32045 );
xor ( n32047 , n32044 , n32045 );
xor ( n32048 , n30909 , n30990 );
nor ( n32049 , n9608 , n31869 );
and ( n32050 , n32048 , n32049 );
xor ( n32051 , n32048 , n32049 );
xor ( n32052 , n30913 , n30988 );
nor ( n32053 , n9617 , n31869 );
and ( n32054 , n32052 , n32053 );
xor ( n32055 , n32052 , n32053 );
xor ( n32056 , n30917 , n30986 );
nor ( n32057 , n9626 , n31869 );
and ( n32058 , n32056 , n32057 );
xor ( n32059 , n32056 , n32057 );
xor ( n32060 , n30921 , n30984 );
nor ( n32061 , n9635 , n31869 );
and ( n32062 , n32060 , n32061 );
xor ( n32063 , n32060 , n32061 );
xor ( n32064 , n30925 , n30982 );
nor ( n32065 , n9644 , n31869 );
and ( n32066 , n32064 , n32065 );
xor ( n32067 , n32064 , n32065 );
xor ( n32068 , n30929 , n30980 );
nor ( n32069 , n9653 , n31869 );
and ( n32070 , n32068 , n32069 );
xor ( n32071 , n32068 , n32069 );
xor ( n32072 , n30933 , n30978 );
nor ( n32073 , n9662 , n31869 );
and ( n32074 , n32072 , n32073 );
xor ( n32075 , n32072 , n32073 );
xor ( n32076 , n30937 , n30976 );
nor ( n32077 , n9671 , n31869 );
and ( n32078 , n32076 , n32077 );
xor ( n32079 , n32076 , n32077 );
xor ( n32080 , n30941 , n30974 );
nor ( n32081 , n9680 , n31869 );
and ( n32082 , n32080 , n32081 );
xor ( n32083 , n32080 , n32081 );
xor ( n32084 , n30945 , n30972 );
nor ( n32085 , n9689 , n31869 );
and ( n32086 , n32084 , n32085 );
xor ( n32087 , n32084 , n32085 );
xor ( n32088 , n30949 , n30970 );
nor ( n32089 , n9698 , n31869 );
and ( n32090 , n32088 , n32089 );
xor ( n32091 , n32088 , n32089 );
xor ( n32092 , n30953 , n30968 );
nor ( n32093 , n9707 , n31869 );
and ( n32094 , n32092 , n32093 );
xor ( n32095 , n32092 , n32093 );
xor ( n32096 , n30957 , n30966 );
nor ( n32097 , n9716 , n31869 );
and ( n32098 , n32096 , n32097 );
xor ( n32099 , n32096 , n32097 );
xor ( n32100 , n30961 , n30964 );
nor ( n32101 , n9725 , n31869 );
and ( n32102 , n32100 , n32101 );
xor ( n32103 , n32100 , n32101 );
xor ( n32104 , n30962 , n30963 );
nor ( n32105 , n9734 , n31869 );
and ( n32106 , n32104 , n32105 );
xor ( n32107 , n32104 , n32105 );
nor ( n32108 , n9752 , n30727 );
nor ( n32109 , n9743 , n31869 );
and ( n32110 , n32108 , n32109 );
and ( n32111 , n32107 , n32110 );
or ( n32112 , n32106 , n32111 );
and ( n32113 , n32103 , n32112 );
or ( n32114 , n32102 , n32113 );
and ( n32115 , n32099 , n32114 );
or ( n32116 , n32098 , n32115 );
and ( n32117 , n32095 , n32116 );
or ( n32118 , n32094 , n32117 );
and ( n32119 , n32091 , n32118 );
or ( n32120 , n32090 , n32119 );
and ( n32121 , n32087 , n32120 );
or ( n32122 , n32086 , n32121 );
and ( n32123 , n32083 , n32122 );
or ( n32124 , n32082 , n32123 );
and ( n32125 , n32079 , n32124 );
or ( n32126 , n32078 , n32125 );
and ( n32127 , n32075 , n32126 );
or ( n32128 , n32074 , n32127 );
and ( n32129 , n32071 , n32128 );
or ( n32130 , n32070 , n32129 );
and ( n32131 , n32067 , n32130 );
or ( n32132 , n32066 , n32131 );
and ( n32133 , n32063 , n32132 );
or ( n32134 , n32062 , n32133 );
and ( n32135 , n32059 , n32134 );
or ( n32136 , n32058 , n32135 );
and ( n32137 , n32055 , n32136 );
or ( n32138 , n32054 , n32137 );
and ( n32139 , n32051 , n32138 );
or ( n32140 , n32050 , n32139 );
and ( n32141 , n32047 , n32140 );
or ( n32142 , n32046 , n32141 );
and ( n32143 , n32043 , n32142 );
or ( n32144 , n32042 , n32143 );
and ( n32145 , n32039 , n32144 );
or ( n32146 , n32038 , n32145 );
and ( n32147 , n32035 , n32146 );
or ( n32148 , n32034 , n32147 );
and ( n32149 , n32031 , n32148 );
or ( n32150 , n32030 , n32149 );
and ( n32151 , n32027 , n32150 );
or ( n32152 , n32026 , n32151 );
and ( n32153 , n32023 , n32152 );
or ( n32154 , n32022 , n32153 );
and ( n32155 , n32019 , n32154 );
or ( n32156 , n32018 , n32155 );
and ( n32157 , n32015 , n32156 );
or ( n32158 , n32014 , n32157 );
and ( n32159 , n32011 , n32158 );
or ( n32160 , n32010 , n32159 );
and ( n32161 , n32007 , n32160 );
or ( n32162 , n32006 , n32161 );
and ( n32163 , n32003 , n32162 );
or ( n32164 , n32002 , n32163 );
and ( n32165 , n31999 , n32164 );
or ( n32166 , n31998 , n32165 );
and ( n32167 , n31995 , n32166 );
or ( n32168 , n31994 , n32167 );
and ( n32169 , n31991 , n32168 );
or ( n32170 , n31990 , n32169 );
and ( n32171 , n31987 , n32170 );
or ( n32172 , n31986 , n32171 );
and ( n32173 , n31983 , n32172 );
or ( n32174 , n31982 , n32173 );
and ( n32175 , n31979 , n32174 );
or ( n32176 , n31978 , n32175 );
and ( n32177 , n31975 , n32176 );
or ( n32178 , n31974 , n32177 );
and ( n32179 , n31971 , n32178 );
or ( n32180 , n31970 , n32179 );
and ( n32181 , n31967 , n32180 );
or ( n32182 , n31966 , n32181 );
and ( n32183 , n31963 , n32182 );
or ( n32184 , n31962 , n32183 );
and ( n32185 , n31959 , n32184 );
or ( n32186 , n31958 , n32185 );
and ( n32187 , n31955 , n32186 );
or ( n32188 , n31954 , n32187 );
and ( n32189 , n31951 , n32188 );
or ( n32190 , n31950 , n32189 );
and ( n32191 , n31947 , n32190 );
or ( n32192 , n31946 , n32191 );
and ( n32193 , n31943 , n32192 );
or ( n32194 , n31942 , n32193 );
and ( n32195 , n31939 , n32194 );
or ( n32196 , n31938 , n32195 );
and ( n32197 , n31935 , n32196 );
or ( n32198 , n31934 , n32197 );
and ( n32199 , n31931 , n32198 );
or ( n32200 , n31930 , n32199 );
and ( n32201 , n31927 , n32200 );
or ( n32202 , n31926 , n32201 );
and ( n32203 , n31923 , n32202 );
or ( n32204 , n31922 , n32203 );
and ( n32205 , n31919 , n32204 );
or ( n32206 , n31918 , n32205 );
and ( n32207 , n31915 , n32206 );
or ( n32208 , n31914 , n32207 );
and ( n32209 , n31911 , n32208 );
or ( n32210 , n31910 , n32209 );
and ( n32211 , n31907 , n32210 );
or ( n32212 , n31906 , n32211 );
and ( n32213 , n31903 , n32212 );
or ( n32214 , n31902 , n32213 );
and ( n32215 , n31899 , n32214 );
or ( n32216 , n31898 , n32215 );
and ( n32217 , n31895 , n32216 );
or ( n32218 , n31894 , n32217 );
and ( n32219 , n31891 , n32218 );
or ( n32220 , n31890 , n32219 );
and ( n32221 , n31887 , n32220 );
or ( n32222 , n31886 , n32221 );
and ( n32223 , n31883 , n32222 );
or ( n32224 , n31882 , n32223 );
and ( n32225 , n31879 , n32224 );
or ( n32226 , n31878 , n32225 );
and ( n32227 , n31875 , n32226 );
or ( n32228 , n31874 , n32227 );
xor ( n32229 , n31871 , n32228 );
buf ( n32230 , n472 );
not ( n32231 , n32230 );
nor ( n32232 , n601 , n32231 );
buf ( n32233 , n32232 );
nor ( n32234 , n622 , n29948 );
xor ( n32235 , n32233 , n32234 );
buf ( n32236 , n32235 );
nor ( n32237 , n646 , n28833 );
xor ( n32238 , n32236 , n32237 );
and ( n32239 , n31085 , n31086 );
buf ( n32240 , n32239 );
xor ( n32241 , n32238 , n32240 );
nor ( n32242 , n684 , n27737 );
xor ( n32243 , n32241 , n32242 );
and ( n32244 , n31088 , n31089 );
and ( n32245 , n31090 , n31092 );
or ( n32246 , n32244 , n32245 );
xor ( n32247 , n32243 , n32246 );
nor ( n32248 , n733 , n26660 );
xor ( n32249 , n32247 , n32248 );
and ( n32250 , n31093 , n31094 );
and ( n32251 , n31095 , n31098 );
or ( n32252 , n32250 , n32251 );
xor ( n32253 , n32249 , n32252 );
nor ( n32254 , n796 , n25600 );
xor ( n32255 , n32253 , n32254 );
and ( n32256 , n31099 , n31100 );
and ( n32257 , n31101 , n31104 );
or ( n32258 , n32256 , n32257 );
xor ( n32259 , n32255 , n32258 );
nor ( n32260 , n868 , n24564 );
xor ( n32261 , n32259 , n32260 );
and ( n32262 , n31105 , n31106 );
and ( n32263 , n31107 , n31110 );
or ( n32264 , n32262 , n32263 );
xor ( n32265 , n32261 , n32264 );
nor ( n32266 , n958 , n23541 );
xor ( n32267 , n32265 , n32266 );
and ( n32268 , n31111 , n31112 );
and ( n32269 , n31113 , n31116 );
or ( n32270 , n32268 , n32269 );
xor ( n32271 , n32267 , n32270 );
nor ( n32272 , n1062 , n22541 );
xor ( n32273 , n32271 , n32272 );
and ( n32274 , n31117 , n31118 );
and ( n32275 , n31119 , n31122 );
or ( n32276 , n32274 , n32275 );
xor ( n32277 , n32273 , n32276 );
nor ( n32278 , n1176 , n21562 );
xor ( n32279 , n32277 , n32278 );
and ( n32280 , n31123 , n31124 );
and ( n32281 , n31125 , n31128 );
or ( n32282 , n32280 , n32281 );
xor ( n32283 , n32279 , n32282 );
nor ( n32284 , n1303 , n20601 );
xor ( n32285 , n32283 , n32284 );
and ( n32286 , n31129 , n31130 );
and ( n32287 , n31131 , n31134 );
or ( n32288 , n32286 , n32287 );
xor ( n32289 , n32285 , n32288 );
nor ( n32290 , n1445 , n19657 );
xor ( n32291 , n32289 , n32290 );
and ( n32292 , n31135 , n31136 );
and ( n32293 , n31137 , n31140 );
or ( n32294 , n32292 , n32293 );
xor ( n32295 , n32291 , n32294 );
nor ( n32296 , n1598 , n18734 );
xor ( n32297 , n32295 , n32296 );
and ( n32298 , n31141 , n31142 );
and ( n32299 , n31143 , n31146 );
or ( n32300 , n32298 , n32299 );
xor ( n32301 , n32297 , n32300 );
nor ( n32302 , n1766 , n17828 );
xor ( n32303 , n32301 , n32302 );
and ( n32304 , n31147 , n31148 );
and ( n32305 , n31149 , n31152 );
or ( n32306 , n32304 , n32305 );
xor ( n32307 , n32303 , n32306 );
nor ( n32308 , n1945 , n16943 );
xor ( n32309 , n32307 , n32308 );
and ( n32310 , n31153 , n31154 );
and ( n32311 , n31155 , n31158 );
or ( n32312 , n32310 , n32311 );
xor ( n32313 , n32309 , n32312 );
nor ( n32314 , n2137 , n16077 );
xor ( n32315 , n32313 , n32314 );
and ( n32316 , n31159 , n31160 );
and ( n32317 , n31161 , n31164 );
or ( n32318 , n32316 , n32317 );
xor ( n32319 , n32315 , n32318 );
nor ( n32320 , n2343 , n15230 );
xor ( n32321 , n32319 , n32320 );
and ( n32322 , n31165 , n31166 );
and ( n32323 , n31167 , n31170 );
or ( n32324 , n32322 , n32323 );
xor ( n32325 , n32321 , n32324 );
nor ( n32326 , n2566 , n14403 );
xor ( n32327 , n32325 , n32326 );
and ( n32328 , n31171 , n31172 );
and ( n32329 , n31173 , n31176 );
or ( n32330 , n32328 , n32329 );
xor ( n32331 , n32327 , n32330 );
nor ( n32332 , n2797 , n13599 );
xor ( n32333 , n32331 , n32332 );
and ( n32334 , n31177 , n31178 );
and ( n32335 , n31179 , n31182 );
or ( n32336 , n32334 , n32335 );
xor ( n32337 , n32333 , n32336 );
nor ( n32338 , n3043 , n12808 );
xor ( n32339 , n32337 , n32338 );
and ( n32340 , n31183 , n31184 );
and ( n32341 , n31185 , n31188 );
or ( n32342 , n32340 , n32341 );
xor ( n32343 , n32339 , n32342 );
nor ( n32344 , n3300 , n12037 );
xor ( n32345 , n32343 , n32344 );
and ( n32346 , n31189 , n31190 );
and ( n32347 , n31191 , n31194 );
or ( n32348 , n32346 , n32347 );
xor ( n32349 , n32345 , n32348 );
nor ( n32350 , n3570 , n11282 );
xor ( n32351 , n32349 , n32350 );
and ( n32352 , n31195 , n31196 );
and ( n32353 , n31197 , n31200 );
or ( n32354 , n32352 , n32353 );
xor ( n32355 , n32351 , n32354 );
nor ( n32356 , n3853 , n10547 );
xor ( n32357 , n32355 , n32356 );
and ( n32358 , n31201 , n31202 );
and ( n32359 , n31203 , n31206 );
or ( n32360 , n32358 , n32359 );
xor ( n32361 , n32357 , n32360 );
nor ( n32362 , n4151 , n9829 );
xor ( n32363 , n32361 , n32362 );
and ( n32364 , n31207 , n31208 );
and ( n32365 , n31209 , n31212 );
or ( n32366 , n32364 , n32365 );
xor ( n32367 , n32363 , n32366 );
nor ( n32368 , n4458 , n8955 );
xor ( n32369 , n32367 , n32368 );
and ( n32370 , n31213 , n31214 );
and ( n32371 , n31215 , n31218 );
or ( n32372 , n32370 , n32371 );
xor ( n32373 , n32369 , n32372 );
nor ( n32374 , n4786 , n603 );
xor ( n32375 , n32373 , n32374 );
and ( n32376 , n31219 , n31220 );
and ( n32377 , n31221 , n31224 );
or ( n32378 , n32376 , n32377 );
xor ( n32379 , n32375 , n32378 );
nor ( n32380 , n5126 , n652 );
xor ( n32381 , n32379 , n32380 );
and ( n32382 , n31225 , n31226 );
and ( n32383 , n31227 , n31230 );
or ( n32384 , n32382 , n32383 );
xor ( n32385 , n32381 , n32384 );
nor ( n32386 , n5477 , n624 );
xor ( n32387 , n32385 , n32386 );
and ( n32388 , n31231 , n31232 );
and ( n32389 , n31233 , n31236 );
or ( n32390 , n32388 , n32389 );
xor ( n32391 , n32387 , n32390 );
nor ( n32392 , n5838 , n648 );
xor ( n32393 , n32391 , n32392 );
and ( n32394 , n31237 , n31238 );
and ( n32395 , n31239 , n31242 );
or ( n32396 , n32394 , n32395 );
xor ( n32397 , n32393 , n32396 );
nor ( n32398 , n6212 , n686 );
xor ( n32399 , n32397 , n32398 );
and ( n32400 , n31243 , n31244 );
and ( n32401 , n31245 , n31248 );
or ( n32402 , n32400 , n32401 );
xor ( n32403 , n32399 , n32402 );
nor ( n32404 , n6596 , n735 );
xor ( n32405 , n32403 , n32404 );
and ( n32406 , n31249 , n31250 );
and ( n32407 , n31251 , n31254 );
or ( n32408 , n32406 , n32407 );
xor ( n32409 , n32405 , n32408 );
nor ( n32410 , n6997 , n798 );
xor ( n32411 , n32409 , n32410 );
and ( n32412 , n31255 , n31256 );
and ( n32413 , n31257 , n31260 );
or ( n32414 , n32412 , n32413 );
xor ( n32415 , n32411 , n32414 );
nor ( n32416 , n7413 , n870 );
xor ( n32417 , n32415 , n32416 );
and ( n32418 , n31261 , n31262 );
and ( n32419 , n31263 , n31266 );
or ( n32420 , n32418 , n32419 );
xor ( n32421 , n32417 , n32420 );
nor ( n32422 , n7841 , n960 );
xor ( n32423 , n32421 , n32422 );
and ( n32424 , n31267 , n31268 );
and ( n32425 , n31269 , n31272 );
or ( n32426 , n32424 , n32425 );
xor ( n32427 , n32423 , n32426 );
nor ( n32428 , n8281 , n1064 );
xor ( n32429 , n32427 , n32428 );
and ( n32430 , n31273 , n31274 );
and ( n32431 , n31275 , n31278 );
or ( n32432 , n32430 , n32431 );
xor ( n32433 , n32429 , n32432 );
nor ( n32434 , n8737 , n1178 );
xor ( n32435 , n32433 , n32434 );
and ( n32436 , n31279 , n31280 );
and ( n32437 , n31281 , n31284 );
or ( n32438 , n32436 , n32437 );
xor ( n32439 , n32435 , n32438 );
nor ( n32440 , n9420 , n1305 );
xor ( n32441 , n32439 , n32440 );
and ( n32442 , n31285 , n31286 );
and ( n32443 , n31287 , n31290 );
or ( n32444 , n32442 , n32443 );
xor ( n32445 , n32441 , n32444 );
nor ( n32446 , n10312 , n1447 );
xor ( n32447 , n32445 , n32446 );
and ( n32448 , n31291 , n31292 );
and ( n32449 , n31293 , n31296 );
or ( n32450 , n32448 , n32449 );
xor ( n32451 , n32447 , n32450 );
nor ( n32452 , n11041 , n1600 );
xor ( n32453 , n32451 , n32452 );
and ( n32454 , n31297 , n31298 );
and ( n32455 , n31299 , n31302 );
or ( n32456 , n32454 , n32455 );
xor ( n32457 , n32453 , n32456 );
nor ( n32458 , n11790 , n1768 );
xor ( n32459 , n32457 , n32458 );
and ( n32460 , n31303 , n31304 );
and ( n32461 , n31305 , n31308 );
or ( n32462 , n32460 , n32461 );
xor ( n32463 , n32459 , n32462 );
nor ( n32464 , n12555 , n1947 );
xor ( n32465 , n32463 , n32464 );
and ( n32466 , n31309 , n31310 );
and ( n32467 , n31311 , n31314 );
or ( n32468 , n32466 , n32467 );
xor ( n32469 , n32465 , n32468 );
nor ( n32470 , n13340 , n2139 );
xor ( n32471 , n32469 , n32470 );
and ( n32472 , n31315 , n31316 );
and ( n32473 , n31317 , n31320 );
or ( n32474 , n32472 , n32473 );
xor ( n32475 , n32471 , n32474 );
nor ( n32476 , n14138 , n2345 );
xor ( n32477 , n32475 , n32476 );
and ( n32478 , n31321 , n31322 );
and ( n32479 , n31323 , n31326 );
or ( n32480 , n32478 , n32479 );
xor ( n32481 , n32477 , n32480 );
nor ( n32482 , n14959 , n2568 );
xor ( n32483 , n32481 , n32482 );
and ( n32484 , n31327 , n31328 );
and ( n32485 , n31329 , n31332 );
or ( n32486 , n32484 , n32485 );
xor ( n32487 , n32483 , n32486 );
nor ( n32488 , n15800 , n2799 );
xor ( n32489 , n32487 , n32488 );
and ( n32490 , n31333 , n31334 );
and ( n32491 , n31335 , n31338 );
or ( n32492 , n32490 , n32491 );
xor ( n32493 , n32489 , n32492 );
nor ( n32494 , n16660 , n3045 );
xor ( n32495 , n32493 , n32494 );
and ( n32496 , n31339 , n31340 );
and ( n32497 , n31341 , n31344 );
or ( n32498 , n32496 , n32497 );
xor ( n32499 , n32495 , n32498 );
nor ( n32500 , n17539 , n3302 );
xor ( n32501 , n32499 , n32500 );
and ( n32502 , n31345 , n31346 );
and ( n32503 , n31347 , n31350 );
or ( n32504 , n32502 , n32503 );
xor ( n32505 , n32501 , n32504 );
nor ( n32506 , n18439 , n3572 );
xor ( n32507 , n32505 , n32506 );
and ( n32508 , n31351 , n31352 );
and ( n32509 , n31353 , n31356 );
or ( n32510 , n32508 , n32509 );
xor ( n32511 , n32507 , n32510 );
nor ( n32512 , n19356 , n3855 );
xor ( n32513 , n32511 , n32512 );
and ( n32514 , n31357 , n31358 );
and ( n32515 , n31359 , n31362 );
or ( n32516 , n32514 , n32515 );
xor ( n32517 , n32513 , n32516 );
nor ( n32518 , n20294 , n4153 );
xor ( n32519 , n32517 , n32518 );
and ( n32520 , n31363 , n31364 );
and ( n32521 , n31365 , n31368 );
or ( n32522 , n32520 , n32521 );
xor ( n32523 , n32519 , n32522 );
nor ( n32524 , n21249 , n4460 );
xor ( n32525 , n32523 , n32524 );
and ( n32526 , n31369 , n31370 );
and ( n32527 , n31371 , n31374 );
or ( n32528 , n32526 , n32527 );
xor ( n32529 , n32525 , n32528 );
nor ( n32530 , n22222 , n4788 );
xor ( n32531 , n32529 , n32530 );
and ( n32532 , n31375 , n31376 );
and ( n32533 , n31377 , n31380 );
or ( n32534 , n32532 , n32533 );
xor ( n32535 , n32531 , n32534 );
nor ( n32536 , n23216 , n5128 );
xor ( n32537 , n32535 , n32536 );
and ( n32538 , n31381 , n31382 );
and ( n32539 , n31383 , n31386 );
or ( n32540 , n32538 , n32539 );
xor ( n32541 , n32537 , n32540 );
nor ( n32542 , n24233 , n5479 );
xor ( n32543 , n32541 , n32542 );
and ( n32544 , n31387 , n31388 );
and ( n32545 , n31389 , n31392 );
or ( n32546 , n32544 , n32545 );
xor ( n32547 , n32543 , n32546 );
nor ( n32548 , n25263 , n5840 );
xor ( n32549 , n32547 , n32548 );
and ( n32550 , n31393 , n31394 );
and ( n32551 , n31395 , n31398 );
or ( n32552 , n32550 , n32551 );
xor ( n32553 , n32549 , n32552 );
nor ( n32554 , n26317 , n6214 );
xor ( n32555 , n32553 , n32554 );
and ( n32556 , n31399 , n31400 );
and ( n32557 , n31401 , n31404 );
or ( n32558 , n32556 , n32557 );
xor ( n32559 , n32555 , n32558 );
nor ( n32560 , n27388 , n6598 );
xor ( n32561 , n32559 , n32560 );
and ( n32562 , n31405 , n31406 );
and ( n32563 , n31407 , n31410 );
or ( n32564 , n32562 , n32563 );
xor ( n32565 , n32561 , n32564 );
nor ( n32566 , n28478 , n6999 );
xor ( n32567 , n32565 , n32566 );
and ( n32568 , n31411 , n31412 );
and ( n32569 , n31413 , n31416 );
or ( n32570 , n32568 , n32569 );
xor ( n32571 , n32567 , n32570 );
nor ( n32572 , n29587 , n7415 );
xor ( n32573 , n32571 , n32572 );
and ( n32574 , n31417 , n31418 );
and ( n32575 , n31419 , n31422 );
or ( n32576 , n32574 , n32575 );
xor ( n32577 , n32573 , n32576 );
nor ( n32578 , n30716 , n7843 );
xor ( n32579 , n32577 , n32578 );
and ( n32580 , n31423 , n31424 );
and ( n32581 , n31425 , n31428 );
or ( n32582 , n32580 , n32581 );
xor ( n32583 , n32579 , n32582 );
nor ( n32584 , n31858 , n8283 );
xor ( n32585 , n32583 , n32584 );
and ( n32586 , n31429 , n31430 );
and ( n32587 , n31431 , n31434 );
or ( n32588 , n32586 , n32587 );
xor ( n32589 , n32585 , n32588 );
and ( n32590 , n31783 , n31784 );
and ( n32591 , n31784 , n31843 );
and ( n32592 , n31783 , n31843 );
or ( n32593 , n32590 , n32591 , n32592 );
and ( n32594 , n31448 , n31778 );
and ( n32595 , n31778 , n31844 );
and ( n32596 , n31448 , n31844 );
or ( n32597 , n32594 , n32595 , n32596 );
xor ( n32598 , n32593 , n32597 );
and ( n32599 , n31452 , n31572 );
and ( n32600 , n31572 , n31777 );
and ( n32601 , n31452 , n31777 );
or ( n32602 , n32599 , n32600 , n32601 );
and ( n32603 , n31456 , n31460 );
and ( n32604 , n31460 , n31571 );
and ( n32605 , n31456 , n31571 );
or ( n32606 , n32603 , n32604 , n32605 );
and ( n32607 , n31786 , n31790 );
and ( n32608 , n31790 , n31842 );
and ( n32609 , n31786 , n31842 );
or ( n32610 , n32607 , n32608 , n32609 );
xor ( n32611 , n32606 , n32610 );
and ( n32612 , n31834 , n31838 );
and ( n32613 , n31795 , n31799 );
and ( n32614 , n31799 , n31841 );
and ( n32615 , n31795 , n31841 );
or ( n32616 , n32613 , n32614 , n32615 );
xor ( n32617 , n32612 , n32616 );
and ( n32618 , n31506 , n31543 );
and ( n32619 , n31543 , n31569 );
and ( n32620 , n31506 , n31569 );
or ( n32621 , n32618 , n32619 , n32620 );
and ( n32622 , n31804 , n31808 );
and ( n32623 , n31808 , n31840 );
and ( n32624 , n31804 , n31840 );
or ( n32625 , n32622 , n32623 , n32624 );
xor ( n32626 , n32621 , n32625 );
and ( n32627 , n31548 , n31552 );
and ( n32628 , n31552 , n31568 );
and ( n32629 , n31548 , n31568 );
or ( n32630 , n32627 , n32628 , n32629 );
and ( n32631 , n31813 , n31829 );
and ( n32632 , n31829 , n31839 );
and ( n32633 , n31813 , n31839 );
or ( n32634 , n32631 , n32632 , n32633 );
xor ( n32635 , n32630 , n32634 );
and ( n32636 , n31817 , n31822 );
and ( n32637 , n31822 , n31828 );
and ( n32638 , n31817 , n31828 );
or ( n32639 , n32636 , n32637 , n32638 );
and ( n32640 , n31818 , n31819 );
and ( n32641 , n31819 , n31821 );
and ( n32642 , n31818 , n31821 );
or ( n32643 , n32640 , n32641 , n32642 );
and ( n32644 , n31835 , n31837 );
xor ( n32645 , n32643 , n32644 );
and ( n32646 , n30695 , n606 );
and ( n32647 , n31836 , n615 );
xor ( n32648 , n32646 , n32647 );
buf ( n32649 , n408 );
and ( n32650 , n32649 , n612 );
xor ( n32651 , n32648 , n32650 );
xor ( n32652 , n32645 , n32651 );
xor ( n32653 , n32639 , n32652 );
and ( n32654 , n31824 , n31825 );
and ( n32655 , n31825 , n31827 );
and ( n32656 , n31824 , n31827 );
or ( n32657 , n32654 , n32655 , n32656 );
and ( n32658 , n27361 , n719 );
and ( n32659 , n28456 , n663 );
xor ( n32660 , n32658 , n32659 );
and ( n32661 , n29559 , n635 );
xor ( n32662 , n32660 , n32661 );
xor ( n32663 , n32657 , n32662 );
and ( n32664 , n24214 , n940 );
and ( n32665 , n25243 , n840 );
xor ( n32666 , n32664 , n32665 );
and ( n32667 , n26296 , n771 );
xor ( n32668 , n32666 , n32667 );
xor ( n32669 , n32663 , n32668 );
xor ( n32670 , n32653 , n32669 );
xor ( n32671 , n32635 , n32670 );
xor ( n32672 , n32626 , n32671 );
xor ( n32673 , n32617 , n32672 );
xor ( n32674 , n32611 , n32673 );
xor ( n32675 , n32602 , n32674 );
and ( n32676 , n31577 , n31652 );
and ( n32677 , n31652 , n31776 );
and ( n32678 , n31577 , n31776 );
or ( n32679 , n32676 , n32677 , n32678 );
and ( n32680 , n31581 , n31585 );
and ( n32681 , n31585 , n31651 );
and ( n32682 , n31581 , n31651 );
or ( n32683 , n32680 , n32681 , n32682 );
and ( n32684 , n31465 , n31501 );
and ( n32685 , n31501 , n31570 );
and ( n32686 , n31465 , n31570 );
or ( n32687 , n32684 , n32685 , n32686 );
xor ( n32688 , n32683 , n32687 );
and ( n32689 , n31469 , n31473 );
and ( n32690 , n31473 , n31500 );
and ( n32691 , n31469 , n31500 );
or ( n32692 , n32689 , n32690 , n32691 );
and ( n32693 , n31510 , n31526 );
and ( n32694 , n31526 , n31542 );
and ( n32695 , n31510 , n31542 );
or ( n32696 , n32693 , n32694 , n32695 );
and ( n32697 , n31557 , n31561 );
and ( n32698 , n31561 , n31567 );
and ( n32699 , n31557 , n31567 );
or ( n32700 , n32697 , n32698 , n32699 );
and ( n32701 , n31514 , n31519 );
and ( n32702 , n31519 , n31525 );
and ( n32703 , n31514 , n31525 );
or ( n32704 , n32701 , n32702 , n32703 );
xor ( n32705 , n32700 , n32704 );
and ( n32706 , n31563 , n31564 );
and ( n32707 , n31564 , n31566 );
and ( n32708 , n31563 , n31566 );
or ( n32709 , n32706 , n32707 , n32708 );
and ( n32710 , n31515 , n31516 );
and ( n32711 , n31516 , n31518 );
and ( n32712 , n31515 , n31518 );
or ( n32713 , n32710 , n32711 , n32712 );
xor ( n32714 , n32709 , n32713 );
and ( n32715 , n21216 , n1254 );
and ( n32716 , n22186 , n1134 );
xor ( n32717 , n32715 , n32716 );
and ( n32718 , n22892 , n1034 );
xor ( n32719 , n32717 , n32718 );
xor ( n32720 , n32714 , n32719 );
xor ( n32721 , n32705 , n32720 );
xor ( n32722 , n32696 , n32721 );
and ( n32723 , n31531 , n31535 );
and ( n32724 , n31535 , n31541 );
and ( n32725 , n31531 , n31541 );
or ( n32726 , n32723 , n32724 , n32725 );
and ( n32727 , n31521 , n31522 );
and ( n32728 , n31522 , n31524 );
and ( n32729 , n31521 , n31524 );
or ( n32730 , n32727 , n32728 , n32729 );
and ( n32731 , n18144 , n1738 );
and ( n32732 , n19324 , n1551 );
xor ( n32733 , n32731 , n32732 );
and ( n32734 , n20233 , n1424 );
xor ( n32735 , n32733 , n32734 );
xor ( n32736 , n32730 , n32735 );
and ( n32737 , n15758 , n2298 );
and ( n32738 , n16637 , n2100 );
xor ( n32739 , n32737 , n32738 );
and ( n32740 , n17512 , n1882 );
xor ( n32741 , n32739 , n32740 );
xor ( n32742 , n32736 , n32741 );
xor ( n32743 , n32726 , n32742 );
and ( n32744 , n31537 , n31538 );
and ( n32745 , n31538 , n31540 );
and ( n32746 , n31537 , n31540 );
or ( n32747 , n32744 , n32745 , n32746 );
and ( n32748 , n31488 , n31489 );
and ( n32749 , n31489 , n31491 );
and ( n32750 , n31488 , n31491 );
or ( n32751 , n32748 , n32749 , n32750 );
xor ( n32752 , n32747 , n32751 );
and ( n32753 , n13322 , n2981 );
and ( n32754 , n14118 , n2739 );
xor ( n32755 , n32753 , n32754 );
and ( n32756 , n14938 , n2544 );
xor ( n32757 , n32755 , n32756 );
xor ( n32758 , n32752 , n32757 );
xor ( n32759 , n32743 , n32758 );
xor ( n32760 , n32722 , n32759 );
xor ( n32761 , n32692 , n32760 );
and ( n32762 , n31478 , n31482 );
and ( n32763 , n31482 , n31499 );
and ( n32764 , n31478 , n31499 );
or ( n32765 , n32762 , n32763 , n32764 );
and ( n32766 , n31594 , n31609 );
and ( n32767 , n31609 , n31623 );
and ( n32768 , n31594 , n31623 );
or ( n32769 , n32766 , n32767 , n32768 );
xor ( n32770 , n32765 , n32769 );
and ( n32771 , n31487 , n31492 );
and ( n32772 , n31492 , n31498 );
and ( n32773 , n31487 , n31498 );
or ( n32774 , n32771 , n32772 , n32773 );
and ( n32775 , n31598 , n31602 );
and ( n32776 , n31602 , n31608 );
and ( n32777 , n31598 , n31608 );
or ( n32778 , n32775 , n32776 , n32777 );
xor ( n32779 , n32774 , n32778 );
and ( n32780 , n31494 , n31495 );
and ( n32781 , n31495 , n31497 );
and ( n32782 , n31494 , n31497 );
or ( n32783 , n32780 , n32781 , n32782 );
and ( n32784 , n11015 , n3749 );
and ( n32785 , n11769 , n3495 );
xor ( n32786 , n32784 , n32785 );
and ( n32787 , n12320 , n3271 );
xor ( n32788 , n32786 , n32787 );
xor ( n32789 , n32783 , n32788 );
and ( n32790 , n8718 , n4730 );
and ( n32791 , n9400 , n4403 );
xor ( n32792 , n32790 , n32791 );
and ( n32793 , n10291 , n4102 );
xor ( n32794 , n32792 , n32793 );
xor ( n32795 , n32789 , n32794 );
xor ( n32796 , n32779 , n32795 );
xor ( n32797 , n32770 , n32796 );
xor ( n32798 , n32761 , n32797 );
xor ( n32799 , n32688 , n32798 );
xor ( n32800 , n32679 , n32799 );
and ( n32801 , n31657 , n31704 );
and ( n32802 , n31704 , n31775 );
and ( n32803 , n31657 , n31775 );
or ( n32804 , n32801 , n32802 , n32803 );
and ( n32805 , n31590 , n31624 );
and ( n32806 , n31624 , n31650 );
and ( n32807 , n31590 , n31650 );
or ( n32808 , n32805 , n32806 , n32807 );
and ( n32809 , n31661 , n31665 );
and ( n32810 , n31665 , n31703 );
and ( n32811 , n31661 , n31703 );
or ( n32812 , n32809 , n32810 , n32811 );
xor ( n32813 , n32808 , n32812 );
and ( n32814 , n31629 , n31633 );
and ( n32815 , n31633 , n31649 );
and ( n32816 , n31629 , n31649 );
or ( n32817 , n32814 , n32815 , n32816 );
and ( n32818 , n31614 , n31616 );
and ( n32819 , n31616 , n31622 );
and ( n32820 , n31614 , n31622 );
or ( n32821 , n32818 , n32819 , n32820 );
and ( n32822 , n31604 , n31605 );
and ( n32823 , n31605 , n31607 );
and ( n32824 , n31604 , n31607 );
or ( n32825 , n32822 , n32823 , n32824 );
and ( n32826 , n6187 , n6504 );
and ( n32827 , n6569 , n6132 );
and ( n32828 , n32826 , n32827 );
and ( n32829 , n32827 , n31615 );
and ( n32830 , n32826 , n31615 );
or ( n32831 , n32828 , n32829 , n32830 );
xor ( n32832 , n32825 , n32831 );
and ( n32833 , n7385 , n5765 );
and ( n32834 , n7808 , n5408 );
xor ( n32835 , n32833 , n32834 );
and ( n32836 , n8079 , n5103 );
xor ( n32837 , n32835 , n32836 );
xor ( n32838 , n32832 , n32837 );
xor ( n32839 , n32821 , n32838 );
and ( n32840 , n31618 , n31619 );
and ( n32841 , n31619 , n31621 );
and ( n32842 , n31618 , n31621 );
or ( n32843 , n32840 , n32841 , n32842 );
and ( n32844 , n6187 , n6971 );
buf ( n32845 , n6569 );
xor ( n32846 , n32844 , n32845 );
and ( n32847 , n6816 , n6132 );
xor ( n32848 , n32846 , n32847 );
xor ( n32849 , n32843 , n32848 );
and ( n32850 , n4959 , n8243 );
and ( n32851 , n5459 , n7662 );
xor ( n32852 , n32850 , n32851 );
and ( n32853 , n5819 , n7310 );
xor ( n32854 , n32852 , n32853 );
xor ( n32855 , n32849 , n32854 );
xor ( n32856 , n32839 , n32855 );
xor ( n32857 , n32817 , n32856 );
and ( n32858 , n31638 , n31642 );
and ( n32859 , n31642 , n31648 );
and ( n32860 , n31638 , n31648 );
or ( n32861 , n32858 , n32859 , n32860 );
and ( n32862 , n31674 , n31679 );
and ( n32863 , n31679 , n31685 );
and ( n32864 , n31674 , n31685 );
or ( n32865 , n32862 , n32863 , n32864 );
xor ( n32866 , n32861 , n32865 );
and ( n32867 , n31675 , n31676 );
and ( n32868 , n31676 , n31678 );
and ( n32869 , n31675 , n31678 );
or ( n32870 , n32867 , n32868 , n32869 );
and ( n32871 , n31644 , n31645 );
and ( n32872 , n31645 , n31647 );
and ( n32873 , n31644 , n31647 );
or ( n32874 , n32871 , n32872 , n32873 );
xor ( n32875 , n32870 , n32874 );
and ( n32876 , n4132 , n10239 );
and ( n32877 , n4438 , n9348 );
xor ( n32878 , n32876 , n32877 );
and ( n32879 , n4766 , n8669 );
xor ( n32880 , n32878 , n32879 );
xor ( n32881 , n32875 , n32880 );
xor ( n32882 , n32866 , n32881 );
xor ( n32883 , n32857 , n32882 );
xor ( n32884 , n32813 , n32883 );
xor ( n32885 , n32804 , n32884 );
and ( n32886 , n31709 , n31735 );
and ( n32887 , n31735 , n31774 );
and ( n32888 , n31709 , n31774 );
or ( n32889 , n32886 , n32887 , n32888 );
and ( n32890 , n31670 , n31686 );
and ( n32891 , n31686 , n31702 );
and ( n32892 , n31670 , n31702 );
or ( n32893 , n32890 , n32891 , n32892 );
and ( n32894 , n31713 , n31717 );
and ( n32895 , n31717 , n31734 );
and ( n32896 , n31713 , n31734 );
or ( n32897 , n32894 , n32895 , n32896 );
xor ( n32898 , n32893 , n32897 );
and ( n32899 , n31691 , n31695 );
and ( n32900 , n31695 , n31701 );
and ( n32901 , n31691 , n31701 );
or ( n32902 , n32899 , n32900 , n32901 );
and ( n32903 , n31681 , n31682 );
and ( n32904 , n31682 , n31684 );
and ( n32905 , n31681 , n31684 );
or ( n32906 , n32903 , n32904 , n32905 );
and ( n32907 , n3182 , n12531 );
and ( n32908 , n3545 , n11718 );
xor ( n32909 , n32907 , n32908 );
and ( n32910 , n3801 , n10977 );
xor ( n32911 , n32909 , n32910 );
xor ( n32912 , n32906 , n32911 );
and ( n32913 , n2462 , n14838 );
and ( n32914 , n2779 , n14044 );
xor ( n32915 , n32913 , n32914 );
and ( n32916 , n3024 , n13256 );
xor ( n32917 , n32915 , n32916 );
xor ( n32918 , n32912 , n32917 );
xor ( n32919 , n32902 , n32918 );
and ( n32920 , n31697 , n31698 );
and ( n32921 , n31698 , n31700 );
and ( n32922 , n31697 , n31700 );
or ( n32923 , n32920 , n32921 , n32922 );
and ( n32924 , n31723 , n31724 );
and ( n32925 , n31724 , n31726 );
and ( n32926 , n31723 , n31726 );
or ( n32927 , n32924 , n32925 , n32926 );
xor ( n32928 , n32923 , n32927 );
and ( n32929 , n1933 , n17422 );
and ( n32930 , n2120 , n16550 );
xor ( n32931 , n32929 , n32930 );
and ( n32932 , n2324 , n15691 );
xor ( n32933 , n32931 , n32932 );
xor ( n32934 , n32928 , n32933 );
xor ( n32935 , n32919 , n32934 );
xor ( n32936 , n32898 , n32935 );
xor ( n32937 , n32889 , n32936 );
and ( n32938 , n31740 , n31755 );
and ( n32939 , n31755 , n31773 );
and ( n32940 , n31740 , n31773 );
or ( n32941 , n32938 , n32939 , n32940 );
and ( n32942 , n31722 , n31727 );
and ( n32943 , n31727 , n31733 );
and ( n32944 , n31722 , n31733 );
or ( n32945 , n32942 , n32943 , n32944 );
and ( n32946 , n31744 , n31748 );
and ( n32947 , n31748 , n31754 );
and ( n32948 , n31744 , n31754 );
or ( n32949 , n32946 , n32947 , n32948 );
xor ( n32950 , n32945 , n32949 );
and ( n32951 , n31729 , n31730 );
and ( n32952 , n31730 , n31732 );
and ( n32953 , n31729 , n31732 );
or ( n32954 , n32951 , n32952 , n32953 );
and ( n32955 , n1383 , n20156 );
and ( n32956 , n1580 , n19222 );
xor ( n32957 , n32955 , n32956 );
and ( n32958 , n1694 , n18407 );
xor ( n32959 , n32957 , n32958 );
xor ( n32960 , n32954 , n32959 );
and ( n32961 , n1047 , n23075 );
and ( n32962 , n1164 , n22065 );
xor ( n32963 , n32961 , n32962 );
and ( n32964 , n1287 , n20976 );
xor ( n32965 , n32963 , n32964 );
xor ( n32966 , n32960 , n32965 );
xor ( n32967 , n32950 , n32966 );
xor ( n32968 , n32941 , n32967 );
and ( n32969 , n31760 , n31766 );
and ( n32970 , n31766 , n31772 );
and ( n32971 , n31760 , n31772 );
or ( n32972 , n32969 , n32970 , n32971 );
and ( n32973 , n31768 , n31769 );
and ( n32974 , n31769 , n31771 );
and ( n32975 , n31768 , n31771 );
or ( n32976 , n32973 , n32974 , n32975 );
and ( n32977 , n31750 , n31751 );
and ( n32978 , n31751 , n31753 );
and ( n32979 , n31750 , n31753 );
or ( n32980 , n32977 , n32978 , n32979 );
xor ( n32981 , n32976 , n32980 );
and ( n32982 , n783 , n26216 );
and ( n32983 , n856 , n25163 );
xor ( n32984 , n32982 , n32983 );
and ( n32985 , n925 , n24137 );
xor ( n32986 , n32984 , n32985 );
xor ( n32987 , n32981 , n32986 );
xor ( n32988 , n32972 , n32987 );
and ( n32989 , n31762 , n31763 );
and ( n32990 , n31763 , n31765 );
and ( n32991 , n31762 , n31765 );
or ( n32992 , n32989 , n32990 , n32991 );
and ( n32993 , n632 , n29508 );
and ( n32994 , n671 , n28406 );
xor ( n32995 , n32993 , n32994 );
and ( n32996 , n715 , n27296 );
xor ( n32997 , n32995 , n32996 );
xor ( n32998 , n32992 , n32997 );
buf ( n32999 , n408 );
and ( n33000 , n599 , n32999 );
and ( n33001 , n608 , n31761 );
xor ( n33002 , n33000 , n33001 );
and ( n33003 , n611 , n30629 );
xor ( n33004 , n33002 , n33003 );
xor ( n33005 , n32998 , n33004 );
xor ( n33006 , n32988 , n33005 );
xor ( n33007 , n32968 , n33006 );
xor ( n33008 , n32937 , n33007 );
xor ( n33009 , n32885 , n33008 );
xor ( n33010 , n32800 , n33009 );
xor ( n33011 , n32675 , n33010 );
xor ( n33012 , n32598 , n33011 );
and ( n33013 , n31439 , n31443 );
and ( n33014 , n31443 , n31845 );
and ( n33015 , n31439 , n31845 );
or ( n33016 , n33013 , n33014 , n33015 );
xor ( n33017 , n33012 , n33016 );
and ( n33018 , n31846 , n31850 );
and ( n33019 , n31851 , n31854 );
or ( n33020 , n33018 , n33019 );
xor ( n33021 , n33017 , n33020 );
buf ( n33022 , n33021 );
buf ( n33023 , n33022 );
not ( n33024 , n33023 );
nor ( n33025 , n33024 , n8739 );
xor ( n33026 , n32589 , n33025 );
and ( n33027 , n31435 , n31859 );
and ( n33028 , n31860 , n31863 );
or ( n33029 , n33027 , n33028 );
xor ( n33030 , n33026 , n33029 );
buf ( n33031 , n33030 );
buf ( n33032 , n33031 );
not ( n33033 , n33032 );
buf ( n33034 , n561 );
not ( n33035 , n33034 );
nor ( n33036 , n33033 , n33035 );
xor ( n33037 , n32229 , n33036 );
xor ( n33038 , n31875 , n32226 );
nor ( n33039 , n31867 , n33035 );
and ( n33040 , n33038 , n33039 );
xor ( n33041 , n33038 , n33039 );
xor ( n33042 , n31879 , n32224 );
nor ( n33043 , n30725 , n33035 );
and ( n33044 , n33042 , n33043 );
xor ( n33045 , n33042 , n33043 );
xor ( n33046 , n31883 , n32222 );
nor ( n33047 , n29596 , n33035 );
and ( n33048 , n33046 , n33047 );
xor ( n33049 , n33046 , n33047 );
xor ( n33050 , n31887 , n32220 );
nor ( n33051 , n28487 , n33035 );
and ( n33052 , n33050 , n33051 );
xor ( n33053 , n33050 , n33051 );
xor ( n33054 , n31891 , n32218 );
nor ( n33055 , n27397 , n33035 );
and ( n33056 , n33054 , n33055 );
xor ( n33057 , n33054 , n33055 );
xor ( n33058 , n31895 , n32216 );
nor ( n33059 , n26326 , n33035 );
and ( n33060 , n33058 , n33059 );
xor ( n33061 , n33058 , n33059 );
xor ( n33062 , n31899 , n32214 );
nor ( n33063 , n25272 , n33035 );
and ( n33064 , n33062 , n33063 );
xor ( n33065 , n33062 , n33063 );
xor ( n33066 , n31903 , n32212 );
nor ( n33067 , n24242 , n33035 );
and ( n33068 , n33066 , n33067 );
xor ( n33069 , n33066 , n33067 );
xor ( n33070 , n31907 , n32210 );
nor ( n33071 , n23225 , n33035 );
and ( n33072 , n33070 , n33071 );
xor ( n33073 , n33070 , n33071 );
xor ( n33074 , n31911 , n32208 );
nor ( n33075 , n22231 , n33035 );
and ( n33076 , n33074 , n33075 );
xor ( n33077 , n33074 , n33075 );
xor ( n33078 , n31915 , n32206 );
nor ( n33079 , n21258 , n33035 );
and ( n33080 , n33078 , n33079 );
xor ( n33081 , n33078 , n33079 );
xor ( n33082 , n31919 , n32204 );
nor ( n33083 , n20303 , n33035 );
and ( n33084 , n33082 , n33083 );
xor ( n33085 , n33082 , n33083 );
xor ( n33086 , n31923 , n32202 );
nor ( n33087 , n19365 , n33035 );
and ( n33088 , n33086 , n33087 );
xor ( n33089 , n33086 , n33087 );
xor ( n33090 , n31927 , n32200 );
nor ( n33091 , n18448 , n33035 );
and ( n33092 , n33090 , n33091 );
xor ( n33093 , n33090 , n33091 );
xor ( n33094 , n31931 , n32198 );
nor ( n33095 , n17548 , n33035 );
and ( n33096 , n33094 , n33095 );
xor ( n33097 , n33094 , n33095 );
xor ( n33098 , n31935 , n32196 );
nor ( n33099 , n16669 , n33035 );
and ( n33100 , n33098 , n33099 );
xor ( n33101 , n33098 , n33099 );
xor ( n33102 , n31939 , n32194 );
nor ( n33103 , n15809 , n33035 );
and ( n33104 , n33102 , n33103 );
xor ( n33105 , n33102 , n33103 );
xor ( n33106 , n31943 , n32192 );
nor ( n33107 , n14968 , n33035 );
and ( n33108 , n33106 , n33107 );
xor ( n33109 , n33106 , n33107 );
xor ( n33110 , n31947 , n32190 );
nor ( n33111 , n14147 , n33035 );
and ( n33112 , n33110 , n33111 );
xor ( n33113 , n33110 , n33111 );
xor ( n33114 , n31951 , n32188 );
nor ( n33115 , n13349 , n33035 );
and ( n33116 , n33114 , n33115 );
xor ( n33117 , n33114 , n33115 );
xor ( n33118 , n31955 , n32186 );
nor ( n33119 , n12564 , n33035 );
and ( n33120 , n33118 , n33119 );
xor ( n33121 , n33118 , n33119 );
xor ( n33122 , n31959 , n32184 );
nor ( n33123 , n11799 , n33035 );
and ( n33124 , n33122 , n33123 );
xor ( n33125 , n33122 , n33123 );
xor ( n33126 , n31963 , n32182 );
nor ( n33127 , n11050 , n33035 );
and ( n33128 , n33126 , n33127 );
xor ( n33129 , n33126 , n33127 );
xor ( n33130 , n31967 , n32180 );
nor ( n33131 , n10321 , n33035 );
and ( n33132 , n33130 , n33131 );
xor ( n33133 , n33130 , n33131 );
xor ( n33134 , n31971 , n32178 );
nor ( n33135 , n9429 , n33035 );
and ( n33136 , n33134 , n33135 );
xor ( n33137 , n33134 , n33135 );
xor ( n33138 , n31975 , n32176 );
nor ( n33139 , n8949 , n33035 );
and ( n33140 , n33138 , n33139 );
xor ( n33141 , n33138 , n33139 );
xor ( n33142 , n31979 , n32174 );
nor ( n33143 , n9437 , n33035 );
and ( n33144 , n33142 , n33143 );
xor ( n33145 , n33142 , n33143 );
xor ( n33146 , n31983 , n32172 );
nor ( n33147 , n9446 , n33035 );
and ( n33148 , n33146 , n33147 );
xor ( n33149 , n33146 , n33147 );
xor ( n33150 , n31987 , n32170 );
nor ( n33151 , n9455 , n33035 );
and ( n33152 , n33150 , n33151 );
xor ( n33153 , n33150 , n33151 );
xor ( n33154 , n31991 , n32168 );
nor ( n33155 , n9464 , n33035 );
and ( n33156 , n33154 , n33155 );
xor ( n33157 , n33154 , n33155 );
xor ( n33158 , n31995 , n32166 );
nor ( n33159 , n9473 , n33035 );
and ( n33160 , n33158 , n33159 );
xor ( n33161 , n33158 , n33159 );
xor ( n33162 , n31999 , n32164 );
nor ( n33163 , n9482 , n33035 );
and ( n33164 , n33162 , n33163 );
xor ( n33165 , n33162 , n33163 );
xor ( n33166 , n32003 , n32162 );
nor ( n33167 , n9491 , n33035 );
and ( n33168 , n33166 , n33167 );
xor ( n33169 , n33166 , n33167 );
xor ( n33170 , n32007 , n32160 );
nor ( n33171 , n9500 , n33035 );
and ( n33172 , n33170 , n33171 );
xor ( n33173 , n33170 , n33171 );
xor ( n33174 , n32011 , n32158 );
nor ( n33175 , n9509 , n33035 );
and ( n33176 , n33174 , n33175 );
xor ( n33177 , n33174 , n33175 );
xor ( n33178 , n32015 , n32156 );
nor ( n33179 , n9518 , n33035 );
and ( n33180 , n33178 , n33179 );
xor ( n33181 , n33178 , n33179 );
xor ( n33182 , n32019 , n32154 );
nor ( n33183 , n9527 , n33035 );
and ( n33184 , n33182 , n33183 );
xor ( n33185 , n33182 , n33183 );
xor ( n33186 , n32023 , n32152 );
nor ( n33187 , n9536 , n33035 );
and ( n33188 , n33186 , n33187 );
xor ( n33189 , n33186 , n33187 );
xor ( n33190 , n32027 , n32150 );
nor ( n33191 , n9545 , n33035 );
and ( n33192 , n33190 , n33191 );
xor ( n33193 , n33190 , n33191 );
xor ( n33194 , n32031 , n32148 );
nor ( n33195 , n9554 , n33035 );
and ( n33196 , n33194 , n33195 );
xor ( n33197 , n33194 , n33195 );
xor ( n33198 , n32035 , n32146 );
nor ( n33199 , n9563 , n33035 );
and ( n33200 , n33198 , n33199 );
xor ( n33201 , n33198 , n33199 );
xor ( n33202 , n32039 , n32144 );
nor ( n33203 , n9572 , n33035 );
and ( n33204 , n33202 , n33203 );
xor ( n33205 , n33202 , n33203 );
xor ( n33206 , n32043 , n32142 );
nor ( n33207 , n9581 , n33035 );
and ( n33208 , n33206 , n33207 );
xor ( n33209 , n33206 , n33207 );
xor ( n33210 , n32047 , n32140 );
nor ( n33211 , n9590 , n33035 );
and ( n33212 , n33210 , n33211 );
xor ( n33213 , n33210 , n33211 );
xor ( n33214 , n32051 , n32138 );
nor ( n33215 , n9599 , n33035 );
and ( n33216 , n33214 , n33215 );
xor ( n33217 , n33214 , n33215 );
xor ( n33218 , n32055 , n32136 );
nor ( n33219 , n9608 , n33035 );
and ( n33220 , n33218 , n33219 );
xor ( n33221 , n33218 , n33219 );
xor ( n33222 , n32059 , n32134 );
nor ( n33223 , n9617 , n33035 );
and ( n33224 , n33222 , n33223 );
xor ( n33225 , n33222 , n33223 );
xor ( n33226 , n32063 , n32132 );
nor ( n33227 , n9626 , n33035 );
and ( n33228 , n33226 , n33227 );
xor ( n33229 , n33226 , n33227 );
xor ( n33230 , n32067 , n32130 );
nor ( n33231 , n9635 , n33035 );
and ( n33232 , n33230 , n33231 );
xor ( n33233 , n33230 , n33231 );
xor ( n33234 , n32071 , n32128 );
nor ( n33235 , n9644 , n33035 );
and ( n33236 , n33234 , n33235 );
xor ( n33237 , n33234 , n33235 );
xor ( n33238 , n32075 , n32126 );
nor ( n33239 , n9653 , n33035 );
and ( n33240 , n33238 , n33239 );
xor ( n33241 , n33238 , n33239 );
xor ( n33242 , n32079 , n32124 );
nor ( n33243 , n9662 , n33035 );
and ( n33244 , n33242 , n33243 );
xor ( n33245 , n33242 , n33243 );
xor ( n33246 , n32083 , n32122 );
nor ( n33247 , n9671 , n33035 );
and ( n33248 , n33246 , n33247 );
xor ( n33249 , n33246 , n33247 );
xor ( n33250 , n32087 , n32120 );
nor ( n33251 , n9680 , n33035 );
and ( n33252 , n33250 , n33251 );
xor ( n33253 , n33250 , n33251 );
xor ( n33254 , n32091 , n32118 );
nor ( n33255 , n9689 , n33035 );
and ( n33256 , n33254 , n33255 );
xor ( n33257 , n33254 , n33255 );
xor ( n33258 , n32095 , n32116 );
nor ( n33259 , n9698 , n33035 );
and ( n33260 , n33258 , n33259 );
xor ( n33261 , n33258 , n33259 );
xor ( n33262 , n32099 , n32114 );
nor ( n33263 , n9707 , n33035 );
and ( n33264 , n33262 , n33263 );
xor ( n33265 , n33262 , n33263 );
xor ( n33266 , n32103 , n32112 );
nor ( n33267 , n9716 , n33035 );
and ( n33268 , n33266 , n33267 );
xor ( n33269 , n33266 , n33267 );
xor ( n33270 , n32107 , n32110 );
nor ( n33271 , n9725 , n33035 );
and ( n33272 , n33270 , n33271 );
xor ( n33273 , n33270 , n33271 );
xor ( n33274 , n32108 , n32109 );
nor ( n33275 , n9734 , n33035 );
and ( n33276 , n33274 , n33275 );
xor ( n33277 , n33274 , n33275 );
nor ( n33278 , n9752 , n31869 );
nor ( n33279 , n9743 , n33035 );
and ( n33280 , n33278 , n33279 );
and ( n33281 , n33277 , n33280 );
or ( n33282 , n33276 , n33281 );
and ( n33283 , n33273 , n33282 );
or ( n33284 , n33272 , n33283 );
and ( n33285 , n33269 , n33284 );
or ( n33286 , n33268 , n33285 );
and ( n33287 , n33265 , n33286 );
or ( n33288 , n33264 , n33287 );
and ( n33289 , n33261 , n33288 );
or ( n33290 , n33260 , n33289 );
and ( n33291 , n33257 , n33290 );
or ( n33292 , n33256 , n33291 );
and ( n33293 , n33253 , n33292 );
or ( n33294 , n33252 , n33293 );
and ( n33295 , n33249 , n33294 );
or ( n33296 , n33248 , n33295 );
and ( n33297 , n33245 , n33296 );
or ( n33298 , n33244 , n33297 );
and ( n33299 , n33241 , n33298 );
or ( n33300 , n33240 , n33299 );
and ( n33301 , n33237 , n33300 );
or ( n33302 , n33236 , n33301 );
and ( n33303 , n33233 , n33302 );
or ( n33304 , n33232 , n33303 );
and ( n33305 , n33229 , n33304 );
or ( n33306 , n33228 , n33305 );
and ( n33307 , n33225 , n33306 );
or ( n33308 , n33224 , n33307 );
and ( n33309 , n33221 , n33308 );
or ( n33310 , n33220 , n33309 );
and ( n33311 , n33217 , n33310 );
or ( n33312 , n33216 , n33311 );
and ( n33313 , n33213 , n33312 );
or ( n33314 , n33212 , n33313 );
and ( n33315 , n33209 , n33314 );
or ( n33316 , n33208 , n33315 );
and ( n33317 , n33205 , n33316 );
or ( n33318 , n33204 , n33317 );
and ( n33319 , n33201 , n33318 );
or ( n33320 , n33200 , n33319 );
and ( n33321 , n33197 , n33320 );
or ( n33322 , n33196 , n33321 );
and ( n33323 , n33193 , n33322 );
or ( n33324 , n33192 , n33323 );
and ( n33325 , n33189 , n33324 );
or ( n33326 , n33188 , n33325 );
and ( n33327 , n33185 , n33326 );
or ( n33328 , n33184 , n33327 );
and ( n33329 , n33181 , n33328 );
or ( n33330 , n33180 , n33329 );
and ( n33331 , n33177 , n33330 );
or ( n33332 , n33176 , n33331 );
and ( n33333 , n33173 , n33332 );
or ( n33334 , n33172 , n33333 );
and ( n33335 , n33169 , n33334 );
or ( n33336 , n33168 , n33335 );
and ( n33337 , n33165 , n33336 );
or ( n33338 , n33164 , n33337 );
and ( n33339 , n33161 , n33338 );
or ( n33340 , n33160 , n33339 );
and ( n33341 , n33157 , n33340 );
or ( n33342 , n33156 , n33341 );
and ( n33343 , n33153 , n33342 );
or ( n33344 , n33152 , n33343 );
and ( n33345 , n33149 , n33344 );
or ( n33346 , n33148 , n33345 );
and ( n33347 , n33145 , n33346 );
or ( n33348 , n33144 , n33347 );
and ( n33349 , n33141 , n33348 );
or ( n33350 , n33140 , n33349 );
and ( n33351 , n33137 , n33350 );
or ( n33352 , n33136 , n33351 );
and ( n33353 , n33133 , n33352 );
or ( n33354 , n33132 , n33353 );
and ( n33355 , n33129 , n33354 );
or ( n33356 , n33128 , n33355 );
and ( n33357 , n33125 , n33356 );
or ( n33358 , n33124 , n33357 );
and ( n33359 , n33121 , n33358 );
or ( n33360 , n33120 , n33359 );
and ( n33361 , n33117 , n33360 );
or ( n33362 , n33116 , n33361 );
and ( n33363 , n33113 , n33362 );
or ( n33364 , n33112 , n33363 );
and ( n33365 , n33109 , n33364 );
or ( n33366 , n33108 , n33365 );
and ( n33367 , n33105 , n33366 );
or ( n33368 , n33104 , n33367 );
and ( n33369 , n33101 , n33368 );
or ( n33370 , n33100 , n33369 );
and ( n33371 , n33097 , n33370 );
or ( n33372 , n33096 , n33371 );
and ( n33373 , n33093 , n33372 );
or ( n33374 , n33092 , n33373 );
and ( n33375 , n33089 , n33374 );
or ( n33376 , n33088 , n33375 );
and ( n33377 , n33085 , n33376 );
or ( n33378 , n33084 , n33377 );
and ( n33379 , n33081 , n33378 );
or ( n33380 , n33080 , n33379 );
and ( n33381 , n33077 , n33380 );
or ( n33382 , n33076 , n33381 );
and ( n33383 , n33073 , n33382 );
or ( n33384 , n33072 , n33383 );
and ( n33385 , n33069 , n33384 );
or ( n33386 , n33068 , n33385 );
and ( n33387 , n33065 , n33386 );
or ( n33388 , n33064 , n33387 );
and ( n33389 , n33061 , n33388 );
or ( n33390 , n33060 , n33389 );
and ( n33391 , n33057 , n33390 );
or ( n33392 , n33056 , n33391 );
and ( n33393 , n33053 , n33392 );
or ( n33394 , n33052 , n33393 );
and ( n33395 , n33049 , n33394 );
or ( n33396 , n33048 , n33395 );
and ( n33397 , n33045 , n33396 );
or ( n33398 , n33044 , n33397 );
and ( n33399 , n33041 , n33398 );
or ( n33400 , n33040 , n33399 );
xor ( n33401 , n33037 , n33400 );
buf ( n33402 , n471 );
not ( n33403 , n33402 );
and ( n33404 , n33403 , n600 );
nor ( n33405 , n601 , n33404 );
buf ( n33406 , n33405 );
nor ( n33407 , n622 , n31083 );
xor ( n33408 , n33406 , n33407 );
buf ( n33409 , n33408 );
nor ( n33410 , n646 , n29948 );
xor ( n33411 , n33409 , n33410 );
and ( n33412 , n32233 , n32234 );
buf ( n33413 , n33412 );
xor ( n33414 , n33411 , n33413 );
nor ( n33415 , n684 , n28833 );
xor ( n33416 , n33414 , n33415 );
and ( n33417 , n32236 , n32237 );
and ( n33418 , n32238 , n32240 );
or ( n33419 , n33417 , n33418 );
xor ( n33420 , n33416 , n33419 );
nor ( n33421 , n733 , n27737 );
xor ( n33422 , n33420 , n33421 );
and ( n33423 , n32241 , n32242 );
and ( n33424 , n32243 , n32246 );
or ( n33425 , n33423 , n33424 );
xor ( n33426 , n33422 , n33425 );
nor ( n33427 , n796 , n26660 );
xor ( n33428 , n33426 , n33427 );
and ( n33429 , n32247 , n32248 );
and ( n33430 , n32249 , n32252 );
or ( n33431 , n33429 , n33430 );
xor ( n33432 , n33428 , n33431 );
nor ( n33433 , n868 , n25600 );
xor ( n33434 , n33432 , n33433 );
and ( n33435 , n32253 , n32254 );
and ( n33436 , n32255 , n32258 );
or ( n33437 , n33435 , n33436 );
xor ( n33438 , n33434 , n33437 );
nor ( n33439 , n958 , n24564 );
xor ( n33440 , n33438 , n33439 );
and ( n33441 , n32259 , n32260 );
and ( n33442 , n32261 , n32264 );
or ( n33443 , n33441 , n33442 );
xor ( n33444 , n33440 , n33443 );
nor ( n33445 , n1062 , n23541 );
xor ( n33446 , n33444 , n33445 );
and ( n33447 , n32265 , n32266 );
and ( n33448 , n32267 , n32270 );
or ( n33449 , n33447 , n33448 );
xor ( n33450 , n33446 , n33449 );
nor ( n33451 , n1176 , n22541 );
xor ( n33452 , n33450 , n33451 );
and ( n33453 , n32271 , n32272 );
and ( n33454 , n32273 , n32276 );
or ( n33455 , n33453 , n33454 );
xor ( n33456 , n33452 , n33455 );
nor ( n33457 , n1303 , n21562 );
xor ( n33458 , n33456 , n33457 );
and ( n33459 , n32277 , n32278 );
and ( n33460 , n32279 , n32282 );
or ( n33461 , n33459 , n33460 );
xor ( n33462 , n33458 , n33461 );
nor ( n33463 , n1445 , n20601 );
xor ( n33464 , n33462 , n33463 );
and ( n33465 , n32283 , n32284 );
and ( n33466 , n32285 , n32288 );
or ( n33467 , n33465 , n33466 );
xor ( n33468 , n33464 , n33467 );
nor ( n33469 , n1598 , n19657 );
xor ( n33470 , n33468 , n33469 );
and ( n33471 , n32289 , n32290 );
and ( n33472 , n32291 , n32294 );
or ( n33473 , n33471 , n33472 );
xor ( n33474 , n33470 , n33473 );
nor ( n33475 , n1766 , n18734 );
xor ( n33476 , n33474 , n33475 );
and ( n33477 , n32295 , n32296 );
and ( n33478 , n32297 , n32300 );
or ( n33479 , n33477 , n33478 );
xor ( n33480 , n33476 , n33479 );
nor ( n33481 , n1945 , n17828 );
xor ( n33482 , n33480 , n33481 );
and ( n33483 , n32301 , n32302 );
and ( n33484 , n32303 , n32306 );
or ( n33485 , n33483 , n33484 );
xor ( n33486 , n33482 , n33485 );
nor ( n33487 , n2137 , n16943 );
xor ( n33488 , n33486 , n33487 );
and ( n33489 , n32307 , n32308 );
and ( n33490 , n32309 , n32312 );
or ( n33491 , n33489 , n33490 );
xor ( n33492 , n33488 , n33491 );
nor ( n33493 , n2343 , n16077 );
xor ( n33494 , n33492 , n33493 );
and ( n33495 , n32313 , n32314 );
and ( n33496 , n32315 , n32318 );
or ( n33497 , n33495 , n33496 );
xor ( n33498 , n33494 , n33497 );
nor ( n33499 , n2566 , n15230 );
xor ( n33500 , n33498 , n33499 );
and ( n33501 , n32319 , n32320 );
and ( n33502 , n32321 , n32324 );
or ( n33503 , n33501 , n33502 );
xor ( n33504 , n33500 , n33503 );
nor ( n33505 , n2797 , n14403 );
xor ( n33506 , n33504 , n33505 );
and ( n33507 , n32325 , n32326 );
and ( n33508 , n32327 , n32330 );
or ( n33509 , n33507 , n33508 );
xor ( n33510 , n33506 , n33509 );
nor ( n33511 , n3043 , n13599 );
xor ( n33512 , n33510 , n33511 );
and ( n33513 , n32331 , n32332 );
and ( n33514 , n32333 , n32336 );
or ( n33515 , n33513 , n33514 );
xor ( n33516 , n33512 , n33515 );
nor ( n33517 , n3300 , n12808 );
xor ( n33518 , n33516 , n33517 );
and ( n33519 , n32337 , n32338 );
and ( n33520 , n32339 , n32342 );
or ( n33521 , n33519 , n33520 );
xor ( n33522 , n33518 , n33521 );
nor ( n33523 , n3570 , n12037 );
xor ( n33524 , n33522 , n33523 );
and ( n33525 , n32343 , n32344 );
and ( n33526 , n32345 , n32348 );
or ( n33527 , n33525 , n33526 );
xor ( n33528 , n33524 , n33527 );
nor ( n33529 , n3853 , n11282 );
xor ( n33530 , n33528 , n33529 );
and ( n33531 , n32349 , n32350 );
and ( n33532 , n32351 , n32354 );
or ( n33533 , n33531 , n33532 );
xor ( n33534 , n33530 , n33533 );
nor ( n33535 , n4151 , n10547 );
xor ( n33536 , n33534 , n33535 );
and ( n33537 , n32355 , n32356 );
and ( n33538 , n32357 , n32360 );
or ( n33539 , n33537 , n33538 );
xor ( n33540 , n33536 , n33539 );
nor ( n33541 , n4458 , n9829 );
xor ( n33542 , n33540 , n33541 );
and ( n33543 , n32361 , n32362 );
and ( n33544 , n32363 , n32366 );
or ( n33545 , n33543 , n33544 );
xor ( n33546 , n33542 , n33545 );
nor ( n33547 , n4786 , n8955 );
xor ( n33548 , n33546 , n33547 );
and ( n33549 , n32367 , n32368 );
and ( n33550 , n32369 , n32372 );
or ( n33551 , n33549 , n33550 );
xor ( n33552 , n33548 , n33551 );
nor ( n33553 , n5126 , n603 );
xor ( n33554 , n33552 , n33553 );
and ( n33555 , n32373 , n32374 );
and ( n33556 , n32375 , n32378 );
or ( n33557 , n33555 , n33556 );
xor ( n33558 , n33554 , n33557 );
nor ( n33559 , n5477 , n652 );
xor ( n33560 , n33558 , n33559 );
and ( n33561 , n32379 , n32380 );
and ( n33562 , n32381 , n32384 );
or ( n33563 , n33561 , n33562 );
xor ( n33564 , n33560 , n33563 );
nor ( n33565 , n5838 , n624 );
xor ( n33566 , n33564 , n33565 );
and ( n33567 , n32385 , n32386 );
and ( n33568 , n32387 , n32390 );
or ( n33569 , n33567 , n33568 );
xor ( n33570 , n33566 , n33569 );
nor ( n33571 , n6212 , n648 );
xor ( n33572 , n33570 , n33571 );
and ( n33573 , n32391 , n32392 );
and ( n33574 , n32393 , n32396 );
or ( n33575 , n33573 , n33574 );
xor ( n33576 , n33572 , n33575 );
nor ( n33577 , n6596 , n686 );
xor ( n33578 , n33576 , n33577 );
and ( n33579 , n32397 , n32398 );
and ( n33580 , n32399 , n32402 );
or ( n33581 , n33579 , n33580 );
xor ( n33582 , n33578 , n33581 );
nor ( n33583 , n6997 , n735 );
xor ( n33584 , n33582 , n33583 );
and ( n33585 , n32403 , n32404 );
and ( n33586 , n32405 , n32408 );
or ( n33587 , n33585 , n33586 );
xor ( n33588 , n33584 , n33587 );
nor ( n33589 , n7413 , n798 );
xor ( n33590 , n33588 , n33589 );
and ( n33591 , n32409 , n32410 );
and ( n33592 , n32411 , n32414 );
or ( n33593 , n33591 , n33592 );
xor ( n33594 , n33590 , n33593 );
nor ( n33595 , n7841 , n870 );
xor ( n33596 , n33594 , n33595 );
and ( n33597 , n32415 , n32416 );
and ( n33598 , n32417 , n32420 );
or ( n33599 , n33597 , n33598 );
xor ( n33600 , n33596 , n33599 );
nor ( n33601 , n8281 , n960 );
xor ( n33602 , n33600 , n33601 );
and ( n33603 , n32421 , n32422 );
and ( n33604 , n32423 , n32426 );
or ( n33605 , n33603 , n33604 );
xor ( n33606 , n33602 , n33605 );
nor ( n33607 , n8737 , n1064 );
xor ( n33608 , n33606 , n33607 );
and ( n33609 , n32427 , n32428 );
and ( n33610 , n32429 , n32432 );
or ( n33611 , n33609 , n33610 );
xor ( n33612 , n33608 , n33611 );
nor ( n33613 , n9420 , n1178 );
xor ( n33614 , n33612 , n33613 );
and ( n33615 , n32433 , n32434 );
and ( n33616 , n32435 , n32438 );
or ( n33617 , n33615 , n33616 );
xor ( n33618 , n33614 , n33617 );
nor ( n33619 , n10312 , n1305 );
xor ( n33620 , n33618 , n33619 );
and ( n33621 , n32439 , n32440 );
and ( n33622 , n32441 , n32444 );
or ( n33623 , n33621 , n33622 );
xor ( n33624 , n33620 , n33623 );
nor ( n33625 , n11041 , n1447 );
xor ( n33626 , n33624 , n33625 );
and ( n33627 , n32445 , n32446 );
and ( n33628 , n32447 , n32450 );
or ( n33629 , n33627 , n33628 );
xor ( n33630 , n33626 , n33629 );
nor ( n33631 , n11790 , n1600 );
xor ( n33632 , n33630 , n33631 );
and ( n33633 , n32451 , n32452 );
and ( n33634 , n32453 , n32456 );
or ( n33635 , n33633 , n33634 );
xor ( n33636 , n33632 , n33635 );
nor ( n33637 , n12555 , n1768 );
xor ( n33638 , n33636 , n33637 );
and ( n33639 , n32457 , n32458 );
and ( n33640 , n32459 , n32462 );
or ( n33641 , n33639 , n33640 );
xor ( n33642 , n33638 , n33641 );
nor ( n33643 , n13340 , n1947 );
xor ( n33644 , n33642 , n33643 );
and ( n33645 , n32463 , n32464 );
and ( n33646 , n32465 , n32468 );
or ( n33647 , n33645 , n33646 );
xor ( n33648 , n33644 , n33647 );
nor ( n33649 , n14138 , n2139 );
xor ( n33650 , n33648 , n33649 );
and ( n33651 , n32469 , n32470 );
and ( n33652 , n32471 , n32474 );
or ( n33653 , n33651 , n33652 );
xor ( n33654 , n33650 , n33653 );
nor ( n33655 , n14959 , n2345 );
xor ( n33656 , n33654 , n33655 );
and ( n33657 , n32475 , n32476 );
and ( n33658 , n32477 , n32480 );
or ( n33659 , n33657 , n33658 );
xor ( n33660 , n33656 , n33659 );
nor ( n33661 , n15800 , n2568 );
xor ( n33662 , n33660 , n33661 );
and ( n33663 , n32481 , n32482 );
and ( n33664 , n32483 , n32486 );
or ( n33665 , n33663 , n33664 );
xor ( n33666 , n33662 , n33665 );
nor ( n33667 , n16660 , n2799 );
xor ( n33668 , n33666 , n33667 );
and ( n33669 , n32487 , n32488 );
and ( n33670 , n32489 , n32492 );
or ( n33671 , n33669 , n33670 );
xor ( n33672 , n33668 , n33671 );
nor ( n33673 , n17539 , n3045 );
xor ( n33674 , n33672 , n33673 );
and ( n33675 , n32493 , n32494 );
and ( n33676 , n32495 , n32498 );
or ( n33677 , n33675 , n33676 );
xor ( n33678 , n33674 , n33677 );
nor ( n33679 , n18439 , n3302 );
xor ( n33680 , n33678 , n33679 );
and ( n33681 , n32499 , n32500 );
and ( n33682 , n32501 , n32504 );
or ( n33683 , n33681 , n33682 );
xor ( n33684 , n33680 , n33683 );
nor ( n33685 , n19356 , n3572 );
xor ( n33686 , n33684 , n33685 );
and ( n33687 , n32505 , n32506 );
and ( n33688 , n32507 , n32510 );
or ( n33689 , n33687 , n33688 );
xor ( n33690 , n33686 , n33689 );
nor ( n33691 , n20294 , n3855 );
xor ( n33692 , n33690 , n33691 );
and ( n33693 , n32511 , n32512 );
and ( n33694 , n32513 , n32516 );
or ( n33695 , n33693 , n33694 );
xor ( n33696 , n33692 , n33695 );
nor ( n33697 , n21249 , n4153 );
xor ( n33698 , n33696 , n33697 );
and ( n33699 , n32517 , n32518 );
and ( n33700 , n32519 , n32522 );
or ( n33701 , n33699 , n33700 );
xor ( n33702 , n33698 , n33701 );
nor ( n33703 , n22222 , n4460 );
xor ( n33704 , n33702 , n33703 );
and ( n33705 , n32523 , n32524 );
and ( n33706 , n32525 , n32528 );
or ( n33707 , n33705 , n33706 );
xor ( n33708 , n33704 , n33707 );
nor ( n33709 , n23216 , n4788 );
xor ( n33710 , n33708 , n33709 );
and ( n33711 , n32529 , n32530 );
and ( n33712 , n32531 , n32534 );
or ( n33713 , n33711 , n33712 );
xor ( n33714 , n33710 , n33713 );
nor ( n33715 , n24233 , n5128 );
xor ( n33716 , n33714 , n33715 );
and ( n33717 , n32535 , n32536 );
and ( n33718 , n32537 , n32540 );
or ( n33719 , n33717 , n33718 );
xor ( n33720 , n33716 , n33719 );
nor ( n33721 , n25263 , n5479 );
xor ( n33722 , n33720 , n33721 );
and ( n33723 , n32541 , n32542 );
and ( n33724 , n32543 , n32546 );
or ( n33725 , n33723 , n33724 );
xor ( n33726 , n33722 , n33725 );
nor ( n33727 , n26317 , n5840 );
xor ( n33728 , n33726 , n33727 );
and ( n33729 , n32547 , n32548 );
and ( n33730 , n32549 , n32552 );
or ( n33731 , n33729 , n33730 );
xor ( n33732 , n33728 , n33731 );
nor ( n33733 , n27388 , n6214 );
xor ( n33734 , n33732 , n33733 );
and ( n33735 , n32553 , n32554 );
and ( n33736 , n32555 , n32558 );
or ( n33737 , n33735 , n33736 );
xor ( n33738 , n33734 , n33737 );
nor ( n33739 , n28478 , n6598 );
xor ( n33740 , n33738 , n33739 );
and ( n33741 , n32559 , n32560 );
and ( n33742 , n32561 , n32564 );
or ( n33743 , n33741 , n33742 );
xor ( n33744 , n33740 , n33743 );
nor ( n33745 , n29587 , n6999 );
xor ( n33746 , n33744 , n33745 );
and ( n33747 , n32565 , n32566 );
and ( n33748 , n32567 , n32570 );
or ( n33749 , n33747 , n33748 );
xor ( n33750 , n33746 , n33749 );
nor ( n33751 , n30716 , n7415 );
xor ( n33752 , n33750 , n33751 );
and ( n33753 , n32571 , n32572 );
and ( n33754 , n32573 , n32576 );
or ( n33755 , n33753 , n33754 );
xor ( n33756 , n33752 , n33755 );
nor ( n33757 , n31858 , n7843 );
xor ( n33758 , n33756 , n33757 );
and ( n33759 , n32577 , n32578 );
and ( n33760 , n32579 , n32582 );
or ( n33761 , n33759 , n33760 );
xor ( n33762 , n33758 , n33761 );
nor ( n33763 , n33024 , n8283 );
xor ( n33764 , n33762 , n33763 );
and ( n33765 , n32583 , n32584 );
and ( n33766 , n32585 , n32588 );
or ( n33767 , n33765 , n33766 );
xor ( n33768 , n33764 , n33767 );
and ( n33769 , n32593 , n32597 );
and ( n33770 , n32597 , n33011 );
and ( n33771 , n32593 , n33011 );
or ( n33772 , n33769 , n33770 , n33771 );
buf ( n33773 , n407 );
not ( n33774 , n33773 );
and ( n33775 , n33774 , n612 );
not ( n33776 , n612 );
nor ( n33777 , n33775 , n33776 );
xor ( n33778 , n33772 , n33777 );
and ( n33779 , n32606 , n32610 );
and ( n33780 , n32610 , n32673 );
and ( n33781 , n32606 , n32673 );
or ( n33782 , n33779 , n33780 , n33781 );
and ( n33783 , n32602 , n32674 );
and ( n33784 , n32674 , n33010 );
and ( n33785 , n32602 , n33010 );
or ( n33786 , n33783 , n33784 , n33785 );
xor ( n33787 , n33782 , n33786 );
and ( n33788 , n32679 , n32799 );
and ( n33789 , n32799 , n33009 );
and ( n33790 , n32679 , n33009 );
or ( n33791 , n33788 , n33789 , n33790 );
and ( n33792 , n32612 , n32616 );
and ( n33793 , n32616 , n32672 );
and ( n33794 , n32612 , n32672 );
or ( n33795 , n33792 , n33793 , n33794 );
and ( n33796 , n32683 , n32687 );
and ( n33797 , n32687 , n32798 );
and ( n33798 , n32683 , n32798 );
or ( n33799 , n33796 , n33797 , n33798 );
xor ( n33800 , n33795 , n33799 );
and ( n33801 , n32643 , n32644 );
and ( n33802 , n32644 , n32651 );
and ( n33803 , n32643 , n32651 );
or ( n33804 , n33801 , n33802 , n33803 );
and ( n33805 , n32621 , n32625 );
and ( n33806 , n32625 , n32671 );
and ( n33807 , n32621 , n32671 );
or ( n33808 , n33805 , n33806 , n33807 );
xor ( n33809 , n33804 , n33808 );
and ( n33810 , n32630 , n32634 );
and ( n33811 , n32634 , n32670 );
and ( n33812 , n32630 , n32670 );
or ( n33813 , n33810 , n33811 , n33812 );
and ( n33814 , n32696 , n32721 );
and ( n33815 , n32721 , n32759 );
and ( n33816 , n32696 , n32759 );
or ( n33817 , n33814 , n33815 , n33816 );
xor ( n33818 , n33813 , n33817 );
and ( n33819 , n32639 , n32652 );
and ( n33820 , n32652 , n32669 );
and ( n33821 , n32639 , n32669 );
or ( n33822 , n33819 , n33820 , n33821 );
and ( n33823 , n32700 , n32704 );
and ( n33824 , n32704 , n32720 );
and ( n33825 , n32700 , n32720 );
or ( n33826 , n33823 , n33824 , n33825 );
xor ( n33827 , n33822 , n33826 );
and ( n33828 , n32657 , n32662 );
and ( n33829 , n32662 , n32668 );
and ( n33830 , n32657 , n32668 );
or ( n33831 , n33828 , n33829 , n33830 );
and ( n33832 , n32646 , n32647 );
and ( n33833 , n32647 , n32650 );
and ( n33834 , n32646 , n32650 );
or ( n33835 , n33832 , n33833 , n33834 );
and ( n33836 , n32658 , n32659 );
and ( n33837 , n32659 , n32661 );
and ( n33838 , n32658 , n32661 );
or ( n33839 , n33836 , n33837 , n33838 );
xor ( n33840 , n33835 , n33839 );
and ( n33841 , n30695 , n635 );
and ( n33842 , n31836 , n606 );
xor ( n33843 , n33841 , n33842 );
and ( n33844 , n32649 , n615 );
xor ( n33845 , n33843 , n33844 );
xor ( n33846 , n33840 , n33845 );
xor ( n33847 , n33831 , n33846 );
and ( n33848 , n32664 , n32665 );
and ( n33849 , n32665 , n32667 );
and ( n33850 , n32664 , n32667 );
or ( n33851 , n33848 , n33849 , n33850 );
and ( n33852 , n27361 , n771 );
and ( n33853 , n28456 , n719 );
xor ( n33854 , n33852 , n33853 );
and ( n33855 , n29559 , n663 );
xor ( n33856 , n33854 , n33855 );
xor ( n33857 , n33851 , n33856 );
and ( n33858 , n24214 , n1034 );
and ( n33859 , n25243 , n940 );
xor ( n33860 , n33858 , n33859 );
and ( n33861 , n26296 , n840 );
xor ( n33862 , n33860 , n33861 );
xor ( n33863 , n33857 , n33862 );
xor ( n33864 , n33847 , n33863 );
xor ( n33865 , n33827 , n33864 );
xor ( n33866 , n33818 , n33865 );
xor ( n33867 , n33809 , n33866 );
xor ( n33868 , n33800 , n33867 );
xor ( n33869 , n33791 , n33868 );
and ( n33870 , n32804 , n32884 );
and ( n33871 , n32884 , n33008 );
and ( n33872 , n32804 , n33008 );
or ( n33873 , n33870 , n33871 , n33872 );
and ( n33874 , n32692 , n32760 );
and ( n33875 , n32760 , n32797 );
and ( n33876 , n32692 , n32797 );
or ( n33877 , n33874 , n33875 , n33876 );
and ( n33878 , n32808 , n32812 );
and ( n33879 , n32812 , n32883 );
and ( n33880 , n32808 , n32883 );
or ( n33881 , n33878 , n33879 , n33880 );
xor ( n33882 , n33877 , n33881 );
and ( n33883 , n32765 , n32769 );
and ( n33884 , n32769 , n32796 );
and ( n33885 , n32765 , n32796 );
or ( n33886 , n33883 , n33884 , n33885 );
and ( n33887 , n32726 , n32742 );
and ( n33888 , n32742 , n32758 );
and ( n33889 , n32726 , n32758 );
or ( n33890 , n33887 , n33888 , n33889 );
and ( n33891 , n32709 , n32713 );
and ( n33892 , n32713 , n32719 );
and ( n33893 , n32709 , n32719 );
or ( n33894 , n33891 , n33892 , n33893 );
and ( n33895 , n32730 , n32735 );
and ( n33896 , n32735 , n32741 );
and ( n33897 , n32730 , n32741 );
or ( n33898 , n33895 , n33896 , n33897 );
xor ( n33899 , n33894 , n33898 );
and ( n33900 , n32715 , n32716 );
and ( n33901 , n32716 , n32718 );
and ( n33902 , n32715 , n32718 );
or ( n33903 , n33900 , n33901 , n33902 );
and ( n33904 , n32731 , n32732 );
and ( n33905 , n32732 , n32734 );
and ( n33906 , n32731 , n32734 );
or ( n33907 , n33904 , n33905 , n33906 );
xor ( n33908 , n33903 , n33907 );
and ( n33909 , n21216 , n1424 );
and ( n33910 , n22186 , n1254 );
xor ( n33911 , n33909 , n33910 );
and ( n33912 , n22892 , n1134 );
xor ( n33913 , n33911 , n33912 );
xor ( n33914 , n33908 , n33913 );
xor ( n33915 , n33899 , n33914 );
xor ( n33916 , n33890 , n33915 );
and ( n33917 , n32747 , n32751 );
and ( n33918 , n32751 , n32757 );
and ( n33919 , n32747 , n32757 );
or ( n33920 , n33917 , n33918 , n33919 );
and ( n33921 , n32737 , n32738 );
and ( n33922 , n32738 , n32740 );
and ( n33923 , n32737 , n32740 );
or ( n33924 , n33921 , n33922 , n33923 );
and ( n33925 , n18144 , n1882 );
and ( n33926 , n19324 , n1738 );
xor ( n33927 , n33925 , n33926 );
and ( n33928 , n20233 , n1551 );
xor ( n33929 , n33927 , n33928 );
xor ( n33930 , n33924 , n33929 );
and ( n33931 , n15758 , n2544 );
and ( n33932 , n16637 , n2298 );
xor ( n33933 , n33931 , n33932 );
and ( n33934 , n17512 , n2100 );
xor ( n33935 , n33933 , n33934 );
xor ( n33936 , n33930 , n33935 );
xor ( n33937 , n33920 , n33936 );
and ( n33938 , n32753 , n32754 );
and ( n33939 , n32754 , n32756 );
and ( n33940 , n32753 , n32756 );
or ( n33941 , n33938 , n33939 , n33940 );
and ( n33942 , n32784 , n32785 );
and ( n33943 , n32785 , n32787 );
and ( n33944 , n32784 , n32787 );
or ( n33945 , n33942 , n33943 , n33944 );
xor ( n33946 , n33941 , n33945 );
and ( n33947 , n13322 , n3271 );
and ( n33948 , n14118 , n2981 );
xor ( n33949 , n33947 , n33948 );
and ( n33950 , n14938 , n2739 );
xor ( n33951 , n33949 , n33950 );
xor ( n33952 , n33946 , n33951 );
xor ( n33953 , n33937 , n33952 );
xor ( n33954 , n33916 , n33953 );
xor ( n33955 , n33886 , n33954 );
and ( n33956 , n32774 , n32778 );
and ( n33957 , n32778 , n32795 );
and ( n33958 , n32774 , n32795 );
or ( n33959 , n33956 , n33957 , n33958 );
and ( n33960 , n32821 , n32838 );
and ( n33961 , n32838 , n32855 );
and ( n33962 , n32821 , n32855 );
or ( n33963 , n33960 , n33961 , n33962 );
xor ( n33964 , n33959 , n33963 );
and ( n33965 , n32783 , n32788 );
and ( n33966 , n32788 , n32794 );
and ( n33967 , n32783 , n32794 );
or ( n33968 , n33965 , n33966 , n33967 );
and ( n33969 , n32825 , n32831 );
and ( n33970 , n32831 , n32837 );
and ( n33971 , n32825 , n32837 );
or ( n33972 , n33969 , n33970 , n33971 );
xor ( n33973 , n33968 , n33972 );
and ( n33974 , n32790 , n32791 );
and ( n33975 , n32791 , n32793 );
and ( n33976 , n32790 , n32793 );
or ( n33977 , n33974 , n33975 , n33976 );
and ( n33978 , n11015 , n4102 );
and ( n33979 , n11769 , n3749 );
xor ( n33980 , n33978 , n33979 );
and ( n33981 , n12320 , n3495 );
xor ( n33982 , n33980 , n33981 );
xor ( n33983 , n33977 , n33982 );
and ( n33984 , n8718 , n5103 );
and ( n33985 , n9400 , n4730 );
xor ( n33986 , n33984 , n33985 );
and ( n33987 , n10291 , n4403 );
xor ( n33988 , n33986 , n33987 );
xor ( n33989 , n33983 , n33988 );
xor ( n33990 , n33973 , n33989 );
xor ( n33991 , n33964 , n33990 );
xor ( n33992 , n33955 , n33991 );
xor ( n33993 , n33882 , n33992 );
xor ( n33994 , n33873 , n33993 );
and ( n33995 , n32889 , n32936 );
and ( n33996 , n32936 , n33007 );
and ( n33997 , n32889 , n33007 );
or ( n33998 , n33995 , n33996 , n33997 );
and ( n33999 , n32817 , n32856 );
and ( n34000 , n32856 , n32882 );
and ( n34001 , n32817 , n32882 );
or ( n34002 , n33999 , n34000 , n34001 );
and ( n34003 , n32893 , n32897 );
and ( n34004 , n32897 , n32935 );
and ( n34005 , n32893 , n32935 );
or ( n34006 , n34003 , n34004 , n34005 );
xor ( n34007 , n34002 , n34006 );
and ( n34008 , n32861 , n32865 );
and ( n34009 , n32865 , n32881 );
and ( n34010 , n32861 , n32881 );
or ( n34011 , n34008 , n34009 , n34010 );
and ( n34012 , n32843 , n32848 );
and ( n34013 , n32848 , n32854 );
and ( n34014 , n32843 , n32854 );
or ( n34015 , n34012 , n34013 , n34014 );
and ( n34016 , n32833 , n32834 );
and ( n34017 , n32834 , n32836 );
and ( n34018 , n32833 , n32836 );
or ( n34019 , n34016 , n34017 , n34018 );
and ( n34020 , n32844 , n32845 );
and ( n34021 , n32845 , n32847 );
and ( n34022 , n32844 , n32847 );
or ( n34023 , n34020 , n34021 , n34022 );
xor ( n34024 , n34019 , n34023 );
and ( n34025 , n7385 , n6132 );
and ( n34026 , n7808 , n5765 );
xor ( n34027 , n34025 , n34026 );
and ( n34028 , n8079 , n5408 );
xor ( n34029 , n34027 , n34028 );
xor ( n34030 , n34024 , n34029 );
xor ( n34031 , n34015 , n34030 );
and ( n34032 , n32850 , n32851 );
and ( n34033 , n32851 , n32853 );
and ( n34034 , n32850 , n32853 );
or ( n34035 , n34032 , n34033 , n34034 );
and ( n34036 , n6187 , n7310 );
and ( n34037 , n6569 , n6971 );
xor ( n34038 , n34036 , n34037 );
and ( n34039 , n6816 , n6504 );
xor ( n34040 , n34038 , n34039 );
xor ( n34041 , n34035 , n34040 );
and ( n34042 , n4959 , n8669 );
and ( n34043 , n5459 , n8243 );
xor ( n34044 , n34042 , n34043 );
and ( n34045 , n5819 , n7662 );
xor ( n34046 , n34044 , n34045 );
xor ( n34047 , n34041 , n34046 );
xor ( n34048 , n34031 , n34047 );
xor ( n34049 , n34011 , n34048 );
and ( n34050 , n32870 , n32874 );
and ( n34051 , n32874 , n32880 );
and ( n34052 , n32870 , n32880 );
or ( n34053 , n34050 , n34051 , n34052 );
and ( n34054 , n32906 , n32911 );
and ( n34055 , n32911 , n32917 );
and ( n34056 , n32906 , n32917 );
or ( n34057 , n34054 , n34055 , n34056 );
xor ( n34058 , n34053 , n34057 );
and ( n34059 , n32876 , n32877 );
and ( n34060 , n32877 , n32879 );
and ( n34061 , n32876 , n32879 );
or ( n34062 , n34059 , n34060 , n34061 );
and ( n34063 , n32907 , n32908 );
and ( n34064 , n32908 , n32910 );
and ( n34065 , n32907 , n32910 );
or ( n34066 , n34063 , n34064 , n34065 );
xor ( n34067 , n34062 , n34066 );
and ( n34068 , n4132 , n10977 );
and ( n34069 , n4438 , n10239 );
xor ( n34070 , n34068 , n34069 );
and ( n34071 , n4766 , n9348 );
xor ( n34072 , n34070 , n34071 );
xor ( n34073 , n34067 , n34072 );
xor ( n34074 , n34058 , n34073 );
xor ( n34075 , n34049 , n34074 );
xor ( n34076 , n34007 , n34075 );
xor ( n34077 , n33998 , n34076 );
and ( n34078 , n32941 , n32967 );
and ( n34079 , n32967 , n33006 );
and ( n34080 , n32941 , n33006 );
or ( n34081 , n34078 , n34079 , n34080 );
and ( n34082 , n32902 , n32918 );
and ( n34083 , n32918 , n32934 );
and ( n34084 , n32902 , n32934 );
or ( n34085 , n34082 , n34083 , n34084 );
and ( n34086 , n32945 , n32949 );
and ( n34087 , n32949 , n32966 );
and ( n34088 , n32945 , n32966 );
or ( n34089 , n34086 , n34087 , n34088 );
xor ( n34090 , n34085 , n34089 );
and ( n34091 , n32923 , n32927 );
and ( n34092 , n32927 , n32933 );
and ( n34093 , n32923 , n32933 );
or ( n34094 , n34091 , n34092 , n34093 );
and ( n34095 , n32913 , n32914 );
and ( n34096 , n32914 , n32916 );
and ( n34097 , n32913 , n32916 );
or ( n34098 , n34095 , n34096 , n34097 );
and ( n34099 , n3182 , n13256 );
and ( n34100 , n3545 , n12531 );
xor ( n34101 , n34099 , n34100 );
and ( n34102 , n3801 , n11718 );
xor ( n34103 , n34101 , n34102 );
xor ( n34104 , n34098 , n34103 );
and ( n34105 , n2462 , n15691 );
and ( n34106 , n2779 , n14838 );
xor ( n34107 , n34105 , n34106 );
and ( n34108 , n3024 , n14044 );
xor ( n34109 , n34107 , n34108 );
xor ( n34110 , n34104 , n34109 );
xor ( n34111 , n34094 , n34110 );
and ( n34112 , n32929 , n32930 );
and ( n34113 , n32930 , n32932 );
and ( n34114 , n32929 , n32932 );
or ( n34115 , n34112 , n34113 , n34114 );
and ( n34116 , n32955 , n32956 );
and ( n34117 , n32956 , n32958 );
and ( n34118 , n32955 , n32958 );
or ( n34119 , n34116 , n34117 , n34118 );
xor ( n34120 , n34115 , n34119 );
and ( n34121 , n1933 , n18407 );
and ( n34122 , n2120 , n17422 );
xor ( n34123 , n34121 , n34122 );
and ( n34124 , n2324 , n16550 );
xor ( n34125 , n34123 , n34124 );
xor ( n34126 , n34120 , n34125 );
xor ( n34127 , n34111 , n34126 );
xor ( n34128 , n34090 , n34127 );
xor ( n34129 , n34081 , n34128 );
and ( n34130 , n32972 , n32987 );
and ( n34131 , n32987 , n33005 );
and ( n34132 , n32972 , n33005 );
or ( n34133 , n34130 , n34131 , n34132 );
and ( n34134 , n32954 , n32959 );
and ( n34135 , n32959 , n32965 );
and ( n34136 , n32954 , n32965 );
or ( n34137 , n34134 , n34135 , n34136 );
and ( n34138 , n32976 , n32980 );
and ( n34139 , n32980 , n32986 );
and ( n34140 , n32976 , n32986 );
or ( n34141 , n34138 , n34139 , n34140 );
xor ( n34142 , n34137 , n34141 );
and ( n34143 , n32961 , n32962 );
and ( n34144 , n32962 , n32964 );
and ( n34145 , n32961 , n32964 );
or ( n34146 , n34143 , n34144 , n34145 );
and ( n34147 , n1383 , n20976 );
and ( n34148 , n1580 , n20156 );
xor ( n34149 , n34147 , n34148 );
and ( n34150 , n1694 , n19222 );
xor ( n34151 , n34149 , n34150 );
xor ( n34152 , n34146 , n34151 );
and ( n34153 , n1047 , n24137 );
and ( n34154 , n1164 , n23075 );
xor ( n34155 , n34153 , n34154 );
and ( n34156 , n1287 , n22065 );
xor ( n34157 , n34155 , n34156 );
xor ( n34158 , n34152 , n34157 );
xor ( n34159 , n34142 , n34158 );
xor ( n34160 , n34133 , n34159 );
and ( n34161 , n32992 , n32997 );
and ( n34162 , n32997 , n33004 );
and ( n34163 , n32992 , n33004 );
or ( n34164 , n34161 , n34162 , n34163 );
and ( n34165 , n32982 , n32983 );
and ( n34166 , n32983 , n32985 );
and ( n34167 , n32982 , n32985 );
or ( n34168 , n34165 , n34166 , n34167 );
and ( n34169 , n32993 , n32994 );
and ( n34170 , n32994 , n32996 );
and ( n34171 , n32993 , n32996 );
or ( n34172 , n34169 , n34170 , n34171 );
xor ( n34173 , n34168 , n34172 );
and ( n34174 , n783 , n27296 );
and ( n34175 , n856 , n26216 );
xor ( n34176 , n34174 , n34175 );
and ( n34177 , n925 , n25163 );
xor ( n34178 , n34176 , n34177 );
xor ( n34179 , n34173 , n34178 );
xor ( n34180 , n34164 , n34179 );
and ( n34181 , n33000 , n33001 );
and ( n34182 , n33001 , n33003 );
and ( n34183 , n33000 , n33003 );
or ( n34184 , n34181 , n34182 , n34183 );
and ( n34185 , n632 , n30629 );
and ( n34186 , n671 , n29508 );
xor ( n34187 , n34185 , n34186 );
and ( n34188 , n715 , n28406 );
xor ( n34189 , n34187 , n34188 );
xor ( n34190 , n34184 , n34189 );
not ( n34191 , n599 );
buf ( n34192 , n407 );
not ( n34193 , n34192 );
and ( n34194 , n34193 , n599 );
nor ( n34195 , n34191 , n34194 );
and ( n34196 , n608 , n32999 );
xor ( n34197 , n34195 , n34196 );
and ( n34198 , n611 , n31761 );
xor ( n34199 , n34197 , n34198 );
xor ( n34200 , n34190 , n34199 );
xor ( n34201 , n34180 , n34200 );
xor ( n34202 , n34160 , n34201 );
xor ( n34203 , n34129 , n34202 );
xor ( n34204 , n34077 , n34203 );
xor ( n34205 , n33994 , n34204 );
xor ( n34206 , n33869 , n34205 );
xor ( n34207 , n33787 , n34206 );
xor ( n34208 , n33778 , n34207 );
and ( n34209 , n33012 , n33016 );
and ( n34210 , n33017 , n33020 );
or ( n34211 , n34209 , n34210 );
xor ( n34212 , n34208 , n34211 );
buf ( n34213 , n34212 );
buf ( n34214 , n34213 );
not ( n34215 , n34214 );
nor ( n34216 , n34215 , n8739 );
xor ( n34217 , n33768 , n34216 );
and ( n34218 , n32589 , n33025 );
and ( n34219 , n33026 , n33029 );
or ( n34220 , n34218 , n34219 );
xor ( n34221 , n34217 , n34220 );
buf ( n34222 , n34221 );
buf ( n34223 , n34222 );
not ( n34224 , n34223 );
buf ( n34225 , n562 );
not ( n34226 , n34225 );
nor ( n34227 , n34224 , n34226 );
xor ( n34228 , n33401 , n34227 );
xor ( n34229 , n33041 , n33398 );
nor ( n34230 , n33033 , n34226 );
and ( n34231 , n34229 , n34230 );
xor ( n34232 , n34229 , n34230 );
xor ( n34233 , n33045 , n33396 );
nor ( n34234 , n31867 , n34226 );
and ( n34235 , n34233 , n34234 );
xor ( n34236 , n34233 , n34234 );
xor ( n34237 , n33049 , n33394 );
nor ( n34238 , n30725 , n34226 );
and ( n34239 , n34237 , n34238 );
xor ( n34240 , n34237 , n34238 );
xor ( n34241 , n33053 , n33392 );
nor ( n34242 , n29596 , n34226 );
and ( n34243 , n34241 , n34242 );
xor ( n34244 , n34241 , n34242 );
xor ( n34245 , n33057 , n33390 );
nor ( n34246 , n28487 , n34226 );
and ( n34247 , n34245 , n34246 );
xor ( n34248 , n34245 , n34246 );
xor ( n34249 , n33061 , n33388 );
nor ( n34250 , n27397 , n34226 );
and ( n34251 , n34249 , n34250 );
xor ( n34252 , n34249 , n34250 );
xor ( n34253 , n33065 , n33386 );
nor ( n34254 , n26326 , n34226 );
and ( n34255 , n34253 , n34254 );
xor ( n34256 , n34253 , n34254 );
xor ( n34257 , n33069 , n33384 );
nor ( n34258 , n25272 , n34226 );
and ( n34259 , n34257 , n34258 );
xor ( n34260 , n34257 , n34258 );
xor ( n34261 , n33073 , n33382 );
nor ( n34262 , n24242 , n34226 );
and ( n34263 , n34261 , n34262 );
xor ( n34264 , n34261 , n34262 );
xor ( n34265 , n33077 , n33380 );
nor ( n34266 , n23225 , n34226 );
and ( n34267 , n34265 , n34266 );
xor ( n34268 , n34265 , n34266 );
xor ( n34269 , n33081 , n33378 );
nor ( n34270 , n22231 , n34226 );
and ( n34271 , n34269 , n34270 );
xor ( n34272 , n34269 , n34270 );
xor ( n34273 , n33085 , n33376 );
nor ( n34274 , n21258 , n34226 );
and ( n34275 , n34273 , n34274 );
xor ( n34276 , n34273 , n34274 );
xor ( n34277 , n33089 , n33374 );
nor ( n34278 , n20303 , n34226 );
and ( n34279 , n34277 , n34278 );
xor ( n34280 , n34277 , n34278 );
xor ( n34281 , n33093 , n33372 );
nor ( n34282 , n19365 , n34226 );
and ( n34283 , n34281 , n34282 );
xor ( n34284 , n34281 , n34282 );
xor ( n34285 , n33097 , n33370 );
nor ( n34286 , n18448 , n34226 );
and ( n34287 , n34285 , n34286 );
xor ( n34288 , n34285 , n34286 );
xor ( n34289 , n33101 , n33368 );
nor ( n34290 , n17548 , n34226 );
and ( n34291 , n34289 , n34290 );
xor ( n34292 , n34289 , n34290 );
xor ( n34293 , n33105 , n33366 );
nor ( n34294 , n16669 , n34226 );
and ( n34295 , n34293 , n34294 );
xor ( n34296 , n34293 , n34294 );
xor ( n34297 , n33109 , n33364 );
nor ( n34298 , n15809 , n34226 );
and ( n34299 , n34297 , n34298 );
xor ( n34300 , n34297 , n34298 );
xor ( n34301 , n33113 , n33362 );
nor ( n34302 , n14968 , n34226 );
and ( n34303 , n34301 , n34302 );
xor ( n34304 , n34301 , n34302 );
xor ( n34305 , n33117 , n33360 );
nor ( n34306 , n14147 , n34226 );
and ( n34307 , n34305 , n34306 );
xor ( n34308 , n34305 , n34306 );
xor ( n34309 , n33121 , n33358 );
nor ( n34310 , n13349 , n34226 );
and ( n34311 , n34309 , n34310 );
xor ( n34312 , n34309 , n34310 );
xor ( n34313 , n33125 , n33356 );
nor ( n34314 , n12564 , n34226 );
and ( n34315 , n34313 , n34314 );
xor ( n34316 , n34313 , n34314 );
xor ( n34317 , n33129 , n33354 );
nor ( n34318 , n11799 , n34226 );
and ( n34319 , n34317 , n34318 );
xor ( n34320 , n34317 , n34318 );
xor ( n34321 , n33133 , n33352 );
nor ( n34322 , n11050 , n34226 );
and ( n34323 , n34321 , n34322 );
xor ( n34324 , n34321 , n34322 );
xor ( n34325 , n33137 , n33350 );
nor ( n34326 , n10321 , n34226 );
and ( n34327 , n34325 , n34326 );
xor ( n34328 , n34325 , n34326 );
xor ( n34329 , n33141 , n33348 );
nor ( n34330 , n9429 , n34226 );
and ( n34331 , n34329 , n34330 );
xor ( n34332 , n34329 , n34330 );
xor ( n34333 , n33145 , n33346 );
nor ( n34334 , n8949 , n34226 );
and ( n34335 , n34333 , n34334 );
xor ( n34336 , n34333 , n34334 );
xor ( n34337 , n33149 , n33344 );
nor ( n34338 , n9437 , n34226 );
and ( n34339 , n34337 , n34338 );
xor ( n34340 , n34337 , n34338 );
xor ( n34341 , n33153 , n33342 );
nor ( n34342 , n9446 , n34226 );
and ( n34343 , n34341 , n34342 );
xor ( n34344 , n34341 , n34342 );
xor ( n34345 , n33157 , n33340 );
nor ( n34346 , n9455 , n34226 );
and ( n34347 , n34345 , n34346 );
xor ( n34348 , n34345 , n34346 );
xor ( n34349 , n33161 , n33338 );
nor ( n34350 , n9464 , n34226 );
and ( n34351 , n34349 , n34350 );
xor ( n34352 , n34349 , n34350 );
xor ( n34353 , n33165 , n33336 );
nor ( n34354 , n9473 , n34226 );
and ( n34355 , n34353 , n34354 );
xor ( n34356 , n34353 , n34354 );
xor ( n34357 , n33169 , n33334 );
nor ( n34358 , n9482 , n34226 );
and ( n34359 , n34357 , n34358 );
xor ( n34360 , n34357 , n34358 );
xor ( n34361 , n33173 , n33332 );
nor ( n34362 , n9491 , n34226 );
and ( n34363 , n34361 , n34362 );
xor ( n34364 , n34361 , n34362 );
xor ( n34365 , n33177 , n33330 );
nor ( n34366 , n9500 , n34226 );
and ( n34367 , n34365 , n34366 );
xor ( n34368 , n34365 , n34366 );
xor ( n34369 , n33181 , n33328 );
nor ( n34370 , n9509 , n34226 );
and ( n34371 , n34369 , n34370 );
xor ( n34372 , n34369 , n34370 );
xor ( n34373 , n33185 , n33326 );
nor ( n34374 , n9518 , n34226 );
and ( n34375 , n34373 , n34374 );
xor ( n34376 , n34373 , n34374 );
xor ( n34377 , n33189 , n33324 );
nor ( n34378 , n9527 , n34226 );
and ( n34379 , n34377 , n34378 );
xor ( n34380 , n34377 , n34378 );
xor ( n34381 , n33193 , n33322 );
nor ( n34382 , n9536 , n34226 );
and ( n34383 , n34381 , n34382 );
xor ( n34384 , n34381 , n34382 );
xor ( n34385 , n33197 , n33320 );
nor ( n34386 , n9545 , n34226 );
and ( n34387 , n34385 , n34386 );
xor ( n34388 , n34385 , n34386 );
xor ( n34389 , n33201 , n33318 );
nor ( n34390 , n9554 , n34226 );
and ( n34391 , n34389 , n34390 );
xor ( n34392 , n34389 , n34390 );
xor ( n34393 , n33205 , n33316 );
nor ( n34394 , n9563 , n34226 );
and ( n34395 , n34393 , n34394 );
xor ( n34396 , n34393 , n34394 );
xor ( n34397 , n33209 , n33314 );
nor ( n34398 , n9572 , n34226 );
and ( n34399 , n34397 , n34398 );
xor ( n34400 , n34397 , n34398 );
xor ( n34401 , n33213 , n33312 );
nor ( n34402 , n9581 , n34226 );
and ( n34403 , n34401 , n34402 );
xor ( n34404 , n34401 , n34402 );
xor ( n34405 , n33217 , n33310 );
nor ( n34406 , n9590 , n34226 );
and ( n34407 , n34405 , n34406 );
xor ( n34408 , n34405 , n34406 );
xor ( n34409 , n33221 , n33308 );
nor ( n34410 , n9599 , n34226 );
and ( n34411 , n34409 , n34410 );
xor ( n34412 , n34409 , n34410 );
xor ( n34413 , n33225 , n33306 );
nor ( n34414 , n9608 , n34226 );
and ( n34415 , n34413 , n34414 );
xor ( n34416 , n34413 , n34414 );
xor ( n34417 , n33229 , n33304 );
nor ( n34418 , n9617 , n34226 );
and ( n34419 , n34417 , n34418 );
xor ( n34420 , n34417 , n34418 );
xor ( n34421 , n33233 , n33302 );
nor ( n34422 , n9626 , n34226 );
and ( n34423 , n34421 , n34422 );
xor ( n34424 , n34421 , n34422 );
xor ( n34425 , n33237 , n33300 );
nor ( n34426 , n9635 , n34226 );
and ( n34427 , n34425 , n34426 );
xor ( n34428 , n34425 , n34426 );
xor ( n34429 , n33241 , n33298 );
nor ( n34430 , n9644 , n34226 );
and ( n34431 , n34429 , n34430 );
xor ( n34432 , n34429 , n34430 );
xor ( n34433 , n33245 , n33296 );
nor ( n34434 , n9653 , n34226 );
and ( n34435 , n34433 , n34434 );
xor ( n34436 , n34433 , n34434 );
xor ( n34437 , n33249 , n33294 );
nor ( n34438 , n9662 , n34226 );
and ( n34439 , n34437 , n34438 );
xor ( n34440 , n34437 , n34438 );
xor ( n34441 , n33253 , n33292 );
nor ( n34442 , n9671 , n34226 );
and ( n34443 , n34441 , n34442 );
xor ( n34444 , n34441 , n34442 );
xor ( n34445 , n33257 , n33290 );
nor ( n34446 , n9680 , n34226 );
and ( n34447 , n34445 , n34446 );
xor ( n34448 , n34445 , n34446 );
xor ( n34449 , n33261 , n33288 );
nor ( n34450 , n9689 , n34226 );
and ( n34451 , n34449 , n34450 );
xor ( n34452 , n34449 , n34450 );
xor ( n34453 , n33265 , n33286 );
nor ( n34454 , n9698 , n34226 );
and ( n34455 , n34453 , n34454 );
xor ( n34456 , n34453 , n34454 );
xor ( n34457 , n33269 , n33284 );
nor ( n34458 , n9707 , n34226 );
and ( n34459 , n34457 , n34458 );
xor ( n34460 , n34457 , n34458 );
xor ( n34461 , n33273 , n33282 );
nor ( n34462 , n9716 , n34226 );
and ( n34463 , n34461 , n34462 );
xor ( n34464 , n34461 , n34462 );
xor ( n34465 , n33277 , n33280 );
nor ( n34466 , n9725 , n34226 );
and ( n34467 , n34465 , n34466 );
xor ( n34468 , n34465 , n34466 );
xor ( n34469 , n33278 , n33279 );
nor ( n34470 , n9734 , n34226 );
and ( n34471 , n34469 , n34470 );
xor ( n34472 , n34469 , n34470 );
nor ( n34473 , n9752 , n33035 );
nor ( n34474 , n9743 , n34226 );
and ( n34475 , n34473 , n34474 );
and ( n34476 , n34472 , n34475 );
or ( n34477 , n34471 , n34476 );
and ( n34478 , n34468 , n34477 );
or ( n34479 , n34467 , n34478 );
and ( n34480 , n34464 , n34479 );
or ( n34481 , n34463 , n34480 );
and ( n34482 , n34460 , n34481 );
or ( n34483 , n34459 , n34482 );
and ( n34484 , n34456 , n34483 );
or ( n34485 , n34455 , n34484 );
and ( n34486 , n34452 , n34485 );
or ( n34487 , n34451 , n34486 );
and ( n34488 , n34448 , n34487 );
or ( n34489 , n34447 , n34488 );
and ( n34490 , n34444 , n34489 );
or ( n34491 , n34443 , n34490 );
and ( n34492 , n34440 , n34491 );
or ( n34493 , n34439 , n34492 );
and ( n34494 , n34436 , n34493 );
or ( n34495 , n34435 , n34494 );
and ( n34496 , n34432 , n34495 );
or ( n34497 , n34431 , n34496 );
and ( n34498 , n34428 , n34497 );
or ( n34499 , n34427 , n34498 );
and ( n34500 , n34424 , n34499 );
or ( n34501 , n34423 , n34500 );
and ( n34502 , n34420 , n34501 );
or ( n34503 , n34419 , n34502 );
and ( n34504 , n34416 , n34503 );
or ( n34505 , n34415 , n34504 );
and ( n34506 , n34412 , n34505 );
or ( n34507 , n34411 , n34506 );
and ( n34508 , n34408 , n34507 );
or ( n34509 , n34407 , n34508 );
and ( n34510 , n34404 , n34509 );
or ( n34511 , n34403 , n34510 );
and ( n34512 , n34400 , n34511 );
or ( n34513 , n34399 , n34512 );
and ( n34514 , n34396 , n34513 );
or ( n34515 , n34395 , n34514 );
and ( n34516 , n34392 , n34515 );
or ( n34517 , n34391 , n34516 );
and ( n34518 , n34388 , n34517 );
or ( n34519 , n34387 , n34518 );
and ( n34520 , n34384 , n34519 );
or ( n34521 , n34383 , n34520 );
and ( n34522 , n34380 , n34521 );
or ( n34523 , n34379 , n34522 );
and ( n34524 , n34376 , n34523 );
or ( n34525 , n34375 , n34524 );
and ( n34526 , n34372 , n34525 );
or ( n34527 , n34371 , n34526 );
and ( n34528 , n34368 , n34527 );
or ( n34529 , n34367 , n34528 );
and ( n34530 , n34364 , n34529 );
or ( n34531 , n34363 , n34530 );
and ( n34532 , n34360 , n34531 );
or ( n34533 , n34359 , n34532 );
and ( n34534 , n34356 , n34533 );
or ( n34535 , n34355 , n34534 );
and ( n34536 , n34352 , n34535 );
or ( n34537 , n34351 , n34536 );
and ( n34538 , n34348 , n34537 );
or ( n34539 , n34347 , n34538 );
and ( n34540 , n34344 , n34539 );
or ( n34541 , n34343 , n34540 );
and ( n34542 , n34340 , n34541 );
or ( n34543 , n34339 , n34542 );
and ( n34544 , n34336 , n34543 );
or ( n34545 , n34335 , n34544 );
and ( n34546 , n34332 , n34545 );
or ( n34547 , n34331 , n34546 );
and ( n34548 , n34328 , n34547 );
or ( n34549 , n34327 , n34548 );
and ( n34550 , n34324 , n34549 );
or ( n34551 , n34323 , n34550 );
and ( n34552 , n34320 , n34551 );
or ( n34553 , n34319 , n34552 );
and ( n34554 , n34316 , n34553 );
or ( n34555 , n34315 , n34554 );
and ( n34556 , n34312 , n34555 );
or ( n34557 , n34311 , n34556 );
and ( n34558 , n34308 , n34557 );
or ( n34559 , n34307 , n34558 );
and ( n34560 , n34304 , n34559 );
or ( n34561 , n34303 , n34560 );
and ( n34562 , n34300 , n34561 );
or ( n34563 , n34299 , n34562 );
and ( n34564 , n34296 , n34563 );
or ( n34565 , n34295 , n34564 );
and ( n34566 , n34292 , n34565 );
or ( n34567 , n34291 , n34566 );
and ( n34568 , n34288 , n34567 );
or ( n34569 , n34287 , n34568 );
and ( n34570 , n34284 , n34569 );
or ( n34571 , n34283 , n34570 );
and ( n34572 , n34280 , n34571 );
or ( n34573 , n34279 , n34572 );
and ( n34574 , n34276 , n34573 );
or ( n34575 , n34275 , n34574 );
and ( n34576 , n34272 , n34575 );
or ( n34577 , n34271 , n34576 );
and ( n34578 , n34268 , n34577 );
or ( n34579 , n34267 , n34578 );
and ( n34580 , n34264 , n34579 );
or ( n34581 , n34263 , n34580 );
and ( n34582 , n34260 , n34581 );
or ( n34583 , n34259 , n34582 );
and ( n34584 , n34256 , n34583 );
or ( n34585 , n34255 , n34584 );
and ( n34586 , n34252 , n34585 );
or ( n34587 , n34251 , n34586 );
and ( n34588 , n34248 , n34587 );
or ( n34589 , n34247 , n34588 );
and ( n34590 , n34244 , n34589 );
or ( n34591 , n34243 , n34590 );
and ( n34592 , n34240 , n34591 );
or ( n34593 , n34239 , n34592 );
and ( n34594 , n34236 , n34593 );
or ( n34595 , n34235 , n34594 );
and ( n34596 , n34232 , n34595 );
or ( n34597 , n34231 , n34596 );
xor ( n34598 , n34228 , n34597 );
nor ( n34599 , n622 , n32231 );
buf ( n34600 , n34599 );
buf ( n34601 , n34600 );
nor ( n34602 , n646 , n31083 );
xor ( n34603 , n34601 , n34602 );
and ( n34604 , n33406 , n33407 );
buf ( n34605 , n34604 );
xor ( n34606 , n34603 , n34605 );
nor ( n34607 , n684 , n29948 );
xor ( n34608 , n34606 , n34607 );
and ( n34609 , n33409 , n33410 );
and ( n34610 , n33411 , n33413 );
or ( n34611 , n34609 , n34610 );
xor ( n34612 , n34608 , n34611 );
nor ( n34613 , n733 , n28833 );
xor ( n34614 , n34612 , n34613 );
and ( n34615 , n33414 , n33415 );
and ( n34616 , n33416 , n33419 );
or ( n34617 , n34615 , n34616 );
xor ( n34618 , n34614 , n34617 );
nor ( n34619 , n796 , n27737 );
xor ( n34620 , n34618 , n34619 );
and ( n34621 , n33420 , n33421 );
and ( n34622 , n33422 , n33425 );
or ( n34623 , n34621 , n34622 );
xor ( n34624 , n34620 , n34623 );
nor ( n34625 , n868 , n26660 );
xor ( n34626 , n34624 , n34625 );
and ( n34627 , n33426 , n33427 );
and ( n34628 , n33428 , n33431 );
or ( n34629 , n34627 , n34628 );
xor ( n34630 , n34626 , n34629 );
nor ( n34631 , n958 , n25600 );
xor ( n34632 , n34630 , n34631 );
and ( n34633 , n33432 , n33433 );
and ( n34634 , n33434 , n33437 );
or ( n34635 , n34633 , n34634 );
xor ( n34636 , n34632 , n34635 );
nor ( n34637 , n1062 , n24564 );
xor ( n34638 , n34636 , n34637 );
and ( n34639 , n33438 , n33439 );
and ( n34640 , n33440 , n33443 );
or ( n34641 , n34639 , n34640 );
xor ( n34642 , n34638 , n34641 );
nor ( n34643 , n1176 , n23541 );
xor ( n34644 , n34642 , n34643 );
and ( n34645 , n33444 , n33445 );
and ( n34646 , n33446 , n33449 );
or ( n34647 , n34645 , n34646 );
xor ( n34648 , n34644 , n34647 );
nor ( n34649 , n1303 , n22541 );
xor ( n34650 , n34648 , n34649 );
and ( n34651 , n33450 , n33451 );
and ( n34652 , n33452 , n33455 );
or ( n34653 , n34651 , n34652 );
xor ( n34654 , n34650 , n34653 );
nor ( n34655 , n1445 , n21562 );
xor ( n34656 , n34654 , n34655 );
and ( n34657 , n33456 , n33457 );
and ( n34658 , n33458 , n33461 );
or ( n34659 , n34657 , n34658 );
xor ( n34660 , n34656 , n34659 );
nor ( n34661 , n1598 , n20601 );
xor ( n34662 , n34660 , n34661 );
and ( n34663 , n33462 , n33463 );
and ( n34664 , n33464 , n33467 );
or ( n34665 , n34663 , n34664 );
xor ( n34666 , n34662 , n34665 );
nor ( n34667 , n1766 , n19657 );
xor ( n34668 , n34666 , n34667 );
and ( n34669 , n33468 , n33469 );
and ( n34670 , n33470 , n33473 );
or ( n34671 , n34669 , n34670 );
xor ( n34672 , n34668 , n34671 );
nor ( n34673 , n1945 , n18734 );
xor ( n34674 , n34672 , n34673 );
and ( n34675 , n33474 , n33475 );
and ( n34676 , n33476 , n33479 );
or ( n34677 , n34675 , n34676 );
xor ( n34678 , n34674 , n34677 );
nor ( n34679 , n2137 , n17828 );
xor ( n34680 , n34678 , n34679 );
and ( n34681 , n33480 , n33481 );
and ( n34682 , n33482 , n33485 );
or ( n34683 , n34681 , n34682 );
xor ( n34684 , n34680 , n34683 );
nor ( n34685 , n2343 , n16943 );
xor ( n34686 , n34684 , n34685 );
and ( n34687 , n33486 , n33487 );
and ( n34688 , n33488 , n33491 );
or ( n34689 , n34687 , n34688 );
xor ( n34690 , n34686 , n34689 );
nor ( n34691 , n2566 , n16077 );
xor ( n34692 , n34690 , n34691 );
and ( n34693 , n33492 , n33493 );
and ( n34694 , n33494 , n33497 );
or ( n34695 , n34693 , n34694 );
xor ( n34696 , n34692 , n34695 );
nor ( n34697 , n2797 , n15230 );
xor ( n34698 , n34696 , n34697 );
and ( n34699 , n33498 , n33499 );
and ( n34700 , n33500 , n33503 );
or ( n34701 , n34699 , n34700 );
xor ( n34702 , n34698 , n34701 );
nor ( n34703 , n3043 , n14403 );
xor ( n34704 , n34702 , n34703 );
and ( n34705 , n33504 , n33505 );
and ( n34706 , n33506 , n33509 );
or ( n34707 , n34705 , n34706 );
xor ( n34708 , n34704 , n34707 );
nor ( n34709 , n3300 , n13599 );
xor ( n34710 , n34708 , n34709 );
and ( n34711 , n33510 , n33511 );
and ( n34712 , n33512 , n33515 );
or ( n34713 , n34711 , n34712 );
xor ( n34714 , n34710 , n34713 );
nor ( n34715 , n3570 , n12808 );
xor ( n34716 , n34714 , n34715 );
and ( n34717 , n33516 , n33517 );
and ( n34718 , n33518 , n33521 );
or ( n34719 , n34717 , n34718 );
xor ( n34720 , n34716 , n34719 );
nor ( n34721 , n3853 , n12037 );
xor ( n34722 , n34720 , n34721 );
and ( n34723 , n33522 , n33523 );
and ( n34724 , n33524 , n33527 );
or ( n34725 , n34723 , n34724 );
xor ( n34726 , n34722 , n34725 );
nor ( n34727 , n4151 , n11282 );
xor ( n34728 , n34726 , n34727 );
and ( n34729 , n33528 , n33529 );
and ( n34730 , n33530 , n33533 );
or ( n34731 , n34729 , n34730 );
xor ( n34732 , n34728 , n34731 );
nor ( n34733 , n4458 , n10547 );
xor ( n34734 , n34732 , n34733 );
and ( n34735 , n33534 , n33535 );
and ( n34736 , n33536 , n33539 );
or ( n34737 , n34735 , n34736 );
xor ( n34738 , n34734 , n34737 );
nor ( n34739 , n4786 , n9829 );
xor ( n34740 , n34738 , n34739 );
and ( n34741 , n33540 , n33541 );
and ( n34742 , n33542 , n33545 );
or ( n34743 , n34741 , n34742 );
xor ( n34744 , n34740 , n34743 );
nor ( n34745 , n5126 , n8955 );
xor ( n34746 , n34744 , n34745 );
and ( n34747 , n33546 , n33547 );
and ( n34748 , n33548 , n33551 );
or ( n34749 , n34747 , n34748 );
xor ( n34750 , n34746 , n34749 );
nor ( n34751 , n5477 , n603 );
xor ( n34752 , n34750 , n34751 );
and ( n34753 , n33552 , n33553 );
and ( n34754 , n33554 , n33557 );
or ( n34755 , n34753 , n34754 );
xor ( n34756 , n34752 , n34755 );
nor ( n34757 , n5838 , n652 );
xor ( n34758 , n34756 , n34757 );
and ( n34759 , n33558 , n33559 );
and ( n34760 , n33560 , n33563 );
or ( n34761 , n34759 , n34760 );
xor ( n34762 , n34758 , n34761 );
nor ( n34763 , n6212 , n624 );
xor ( n34764 , n34762 , n34763 );
and ( n34765 , n33564 , n33565 );
and ( n34766 , n33566 , n33569 );
or ( n34767 , n34765 , n34766 );
xor ( n34768 , n34764 , n34767 );
nor ( n34769 , n6596 , n648 );
xor ( n34770 , n34768 , n34769 );
and ( n34771 , n33570 , n33571 );
and ( n34772 , n33572 , n33575 );
or ( n34773 , n34771 , n34772 );
xor ( n34774 , n34770 , n34773 );
nor ( n34775 , n6997 , n686 );
xor ( n34776 , n34774 , n34775 );
and ( n34777 , n33576 , n33577 );
and ( n34778 , n33578 , n33581 );
or ( n34779 , n34777 , n34778 );
xor ( n34780 , n34776 , n34779 );
nor ( n34781 , n7413 , n735 );
xor ( n34782 , n34780 , n34781 );
and ( n34783 , n33582 , n33583 );
and ( n34784 , n33584 , n33587 );
or ( n34785 , n34783 , n34784 );
xor ( n34786 , n34782 , n34785 );
nor ( n34787 , n7841 , n798 );
xor ( n34788 , n34786 , n34787 );
and ( n34789 , n33588 , n33589 );
and ( n34790 , n33590 , n33593 );
or ( n34791 , n34789 , n34790 );
xor ( n34792 , n34788 , n34791 );
nor ( n34793 , n8281 , n870 );
xor ( n34794 , n34792 , n34793 );
and ( n34795 , n33594 , n33595 );
and ( n34796 , n33596 , n33599 );
or ( n34797 , n34795 , n34796 );
xor ( n34798 , n34794 , n34797 );
nor ( n34799 , n8737 , n960 );
xor ( n34800 , n34798 , n34799 );
and ( n34801 , n33600 , n33601 );
and ( n34802 , n33602 , n33605 );
or ( n34803 , n34801 , n34802 );
xor ( n34804 , n34800 , n34803 );
nor ( n34805 , n9420 , n1064 );
xor ( n34806 , n34804 , n34805 );
and ( n34807 , n33606 , n33607 );
and ( n34808 , n33608 , n33611 );
or ( n34809 , n34807 , n34808 );
xor ( n34810 , n34806 , n34809 );
nor ( n34811 , n10312 , n1178 );
xor ( n34812 , n34810 , n34811 );
and ( n34813 , n33612 , n33613 );
and ( n34814 , n33614 , n33617 );
or ( n34815 , n34813 , n34814 );
xor ( n34816 , n34812 , n34815 );
nor ( n34817 , n11041 , n1305 );
xor ( n34818 , n34816 , n34817 );
and ( n34819 , n33618 , n33619 );
and ( n34820 , n33620 , n33623 );
or ( n34821 , n34819 , n34820 );
xor ( n34822 , n34818 , n34821 );
nor ( n34823 , n11790 , n1447 );
xor ( n34824 , n34822 , n34823 );
and ( n34825 , n33624 , n33625 );
and ( n34826 , n33626 , n33629 );
or ( n34827 , n34825 , n34826 );
xor ( n34828 , n34824 , n34827 );
nor ( n34829 , n12555 , n1600 );
xor ( n34830 , n34828 , n34829 );
and ( n34831 , n33630 , n33631 );
and ( n34832 , n33632 , n33635 );
or ( n34833 , n34831 , n34832 );
xor ( n34834 , n34830 , n34833 );
nor ( n34835 , n13340 , n1768 );
xor ( n34836 , n34834 , n34835 );
and ( n34837 , n33636 , n33637 );
and ( n34838 , n33638 , n33641 );
or ( n34839 , n34837 , n34838 );
xor ( n34840 , n34836 , n34839 );
nor ( n34841 , n14138 , n1947 );
xor ( n34842 , n34840 , n34841 );
and ( n34843 , n33642 , n33643 );
and ( n34844 , n33644 , n33647 );
or ( n34845 , n34843 , n34844 );
xor ( n34846 , n34842 , n34845 );
nor ( n34847 , n14959 , n2139 );
xor ( n34848 , n34846 , n34847 );
and ( n34849 , n33648 , n33649 );
and ( n34850 , n33650 , n33653 );
or ( n34851 , n34849 , n34850 );
xor ( n34852 , n34848 , n34851 );
nor ( n34853 , n15800 , n2345 );
xor ( n34854 , n34852 , n34853 );
and ( n34855 , n33654 , n33655 );
and ( n34856 , n33656 , n33659 );
or ( n34857 , n34855 , n34856 );
xor ( n34858 , n34854 , n34857 );
nor ( n34859 , n16660 , n2568 );
xor ( n34860 , n34858 , n34859 );
and ( n34861 , n33660 , n33661 );
and ( n34862 , n33662 , n33665 );
or ( n34863 , n34861 , n34862 );
xor ( n34864 , n34860 , n34863 );
nor ( n34865 , n17539 , n2799 );
xor ( n34866 , n34864 , n34865 );
and ( n34867 , n33666 , n33667 );
and ( n34868 , n33668 , n33671 );
or ( n34869 , n34867 , n34868 );
xor ( n34870 , n34866 , n34869 );
nor ( n34871 , n18439 , n3045 );
xor ( n34872 , n34870 , n34871 );
and ( n34873 , n33672 , n33673 );
and ( n34874 , n33674 , n33677 );
or ( n34875 , n34873 , n34874 );
xor ( n34876 , n34872 , n34875 );
nor ( n34877 , n19356 , n3302 );
xor ( n34878 , n34876 , n34877 );
and ( n34879 , n33678 , n33679 );
and ( n34880 , n33680 , n33683 );
or ( n34881 , n34879 , n34880 );
xor ( n34882 , n34878 , n34881 );
nor ( n34883 , n20294 , n3572 );
xor ( n34884 , n34882 , n34883 );
and ( n34885 , n33684 , n33685 );
and ( n34886 , n33686 , n33689 );
or ( n34887 , n34885 , n34886 );
xor ( n34888 , n34884 , n34887 );
nor ( n34889 , n21249 , n3855 );
xor ( n34890 , n34888 , n34889 );
and ( n34891 , n33690 , n33691 );
and ( n34892 , n33692 , n33695 );
or ( n34893 , n34891 , n34892 );
xor ( n34894 , n34890 , n34893 );
nor ( n34895 , n22222 , n4153 );
xor ( n34896 , n34894 , n34895 );
and ( n34897 , n33696 , n33697 );
and ( n34898 , n33698 , n33701 );
or ( n34899 , n34897 , n34898 );
xor ( n34900 , n34896 , n34899 );
nor ( n34901 , n23216 , n4460 );
xor ( n34902 , n34900 , n34901 );
and ( n34903 , n33702 , n33703 );
and ( n34904 , n33704 , n33707 );
or ( n34905 , n34903 , n34904 );
xor ( n34906 , n34902 , n34905 );
nor ( n34907 , n24233 , n4788 );
xor ( n34908 , n34906 , n34907 );
and ( n34909 , n33708 , n33709 );
and ( n34910 , n33710 , n33713 );
or ( n34911 , n34909 , n34910 );
xor ( n34912 , n34908 , n34911 );
nor ( n34913 , n25263 , n5128 );
xor ( n34914 , n34912 , n34913 );
and ( n34915 , n33714 , n33715 );
and ( n34916 , n33716 , n33719 );
or ( n34917 , n34915 , n34916 );
xor ( n34918 , n34914 , n34917 );
nor ( n34919 , n26317 , n5479 );
xor ( n34920 , n34918 , n34919 );
and ( n34921 , n33720 , n33721 );
and ( n34922 , n33722 , n33725 );
or ( n34923 , n34921 , n34922 );
xor ( n34924 , n34920 , n34923 );
nor ( n34925 , n27388 , n5840 );
xor ( n34926 , n34924 , n34925 );
and ( n34927 , n33726 , n33727 );
and ( n34928 , n33728 , n33731 );
or ( n34929 , n34927 , n34928 );
xor ( n34930 , n34926 , n34929 );
nor ( n34931 , n28478 , n6214 );
xor ( n34932 , n34930 , n34931 );
and ( n34933 , n33732 , n33733 );
and ( n34934 , n33734 , n33737 );
or ( n34935 , n34933 , n34934 );
xor ( n34936 , n34932 , n34935 );
nor ( n34937 , n29587 , n6598 );
xor ( n34938 , n34936 , n34937 );
and ( n34939 , n33738 , n33739 );
and ( n34940 , n33740 , n33743 );
or ( n34941 , n34939 , n34940 );
xor ( n34942 , n34938 , n34941 );
nor ( n34943 , n30716 , n6999 );
xor ( n34944 , n34942 , n34943 );
and ( n34945 , n33744 , n33745 );
and ( n34946 , n33746 , n33749 );
or ( n34947 , n34945 , n34946 );
xor ( n34948 , n34944 , n34947 );
nor ( n34949 , n31858 , n7415 );
xor ( n34950 , n34948 , n34949 );
and ( n34951 , n33750 , n33751 );
and ( n34952 , n33752 , n33755 );
or ( n34953 , n34951 , n34952 );
xor ( n34954 , n34950 , n34953 );
nor ( n34955 , n33024 , n7843 );
xor ( n34956 , n34954 , n34955 );
and ( n34957 , n33756 , n33757 );
and ( n34958 , n33758 , n33761 );
or ( n34959 , n34957 , n34958 );
xor ( n34960 , n34956 , n34959 );
nor ( n34961 , n34215 , n8283 );
xor ( n34962 , n34960 , n34961 );
and ( n34963 , n33762 , n33763 );
and ( n34964 , n33764 , n33767 );
or ( n34965 , n34963 , n34964 );
xor ( n34966 , n34962 , n34965 );
and ( n34967 , n33782 , n33786 );
and ( n34968 , n33786 , n34206 );
and ( n34969 , n33782 , n34206 );
or ( n34970 , n34967 , n34968 , n34969 );
and ( n34971 , n33774 , n615 );
not ( n34972 , n615 );
nor ( n34973 , n34971 , n34972 );
xor ( n34974 , n34970 , n34973 );
and ( n34975 , n33795 , n33799 );
and ( n34976 , n33799 , n33867 );
and ( n34977 , n33795 , n33867 );
or ( n34978 , n34975 , n34976 , n34977 );
and ( n34979 , n33791 , n33868 );
and ( n34980 , n33868 , n34205 );
and ( n34981 , n33791 , n34205 );
or ( n34982 , n34979 , n34980 , n34981 );
xor ( n34983 , n34978 , n34982 );
and ( n34984 , n33873 , n33993 );
and ( n34985 , n33993 , n34204 );
and ( n34986 , n33873 , n34204 );
or ( n34987 , n34984 , n34985 , n34986 );
and ( n34988 , n33804 , n33808 );
and ( n34989 , n33808 , n33866 );
and ( n34990 , n33804 , n33866 );
or ( n34991 , n34988 , n34989 , n34990 );
and ( n34992 , n33877 , n33881 );
and ( n34993 , n33881 , n33992 );
and ( n34994 , n33877 , n33992 );
or ( n34995 , n34992 , n34993 , n34994 );
xor ( n34996 , n34991 , n34995 );
and ( n34997 , n33835 , n33839 );
and ( n34998 , n33839 , n33845 );
and ( n34999 , n33835 , n33845 );
or ( n35000 , n34997 , n34998 , n34999 );
and ( n35001 , n33813 , n33817 );
and ( n35002 , n33817 , n33865 );
and ( n35003 , n33813 , n33865 );
or ( n35004 , n35001 , n35002 , n35003 );
xor ( n35005 , n35000 , n35004 );
and ( n35006 , n33822 , n33826 );
and ( n35007 , n33826 , n33864 );
and ( n35008 , n33822 , n33864 );
or ( n35009 , n35006 , n35007 , n35008 );
and ( n35010 , n33890 , n33915 );
and ( n35011 , n33915 , n33953 );
and ( n35012 , n33890 , n33953 );
or ( n35013 , n35010 , n35011 , n35012 );
xor ( n35014 , n35009 , n35013 );
and ( n35015 , n33831 , n33846 );
and ( n35016 , n33846 , n33863 );
and ( n35017 , n33831 , n33863 );
or ( n35018 , n35015 , n35016 , n35017 );
and ( n35019 , n33894 , n33898 );
and ( n35020 , n33898 , n33914 );
and ( n35021 , n33894 , n33914 );
or ( n35022 , n35019 , n35020 , n35021 );
xor ( n35023 , n35018 , n35022 );
and ( n35024 , n33851 , n33856 );
and ( n35025 , n33856 , n33862 );
and ( n35026 , n33851 , n33862 );
or ( n35027 , n35024 , n35025 , n35026 );
and ( n35028 , n33841 , n33842 );
and ( n35029 , n33842 , n33844 );
and ( n35030 , n33841 , n33844 );
or ( n35031 , n35028 , n35029 , n35030 );
and ( n35032 , n33852 , n33853 );
and ( n35033 , n33853 , n33855 );
and ( n35034 , n33852 , n33855 );
or ( n35035 , n35032 , n35033 , n35034 );
xor ( n35036 , n35031 , n35035 );
and ( n35037 , n30695 , n663 );
and ( n35038 , n31836 , n635 );
xor ( n35039 , n35037 , n35038 );
and ( n35040 , n32649 , n606 );
xor ( n35041 , n35039 , n35040 );
xor ( n35042 , n35036 , n35041 );
xor ( n35043 , n35027 , n35042 );
and ( n35044 , n33858 , n33859 );
and ( n35045 , n33859 , n33861 );
and ( n35046 , n33858 , n33861 );
or ( n35047 , n35044 , n35045 , n35046 );
and ( n35048 , n27361 , n840 );
and ( n35049 , n28456 , n771 );
xor ( n35050 , n35048 , n35049 );
and ( n35051 , n29559 , n719 );
xor ( n35052 , n35050 , n35051 );
xor ( n35053 , n35047 , n35052 );
and ( n35054 , n24214 , n1134 );
and ( n35055 , n25243 , n1034 );
xor ( n35056 , n35054 , n35055 );
and ( n35057 , n26296 , n940 );
xor ( n35058 , n35056 , n35057 );
xor ( n35059 , n35053 , n35058 );
xor ( n35060 , n35043 , n35059 );
xor ( n35061 , n35023 , n35060 );
xor ( n35062 , n35014 , n35061 );
xor ( n35063 , n35005 , n35062 );
xor ( n35064 , n34996 , n35063 );
xor ( n35065 , n34987 , n35064 );
and ( n35066 , n33998 , n34076 );
and ( n35067 , n34076 , n34203 );
and ( n35068 , n33998 , n34203 );
or ( n35069 , n35066 , n35067 , n35068 );
and ( n35070 , n33886 , n33954 );
and ( n35071 , n33954 , n33991 );
and ( n35072 , n33886 , n33991 );
or ( n35073 , n35070 , n35071 , n35072 );
and ( n35074 , n34002 , n34006 );
and ( n35075 , n34006 , n34075 );
and ( n35076 , n34002 , n34075 );
or ( n35077 , n35074 , n35075 , n35076 );
xor ( n35078 , n35073 , n35077 );
and ( n35079 , n33959 , n33963 );
and ( n35080 , n33963 , n33990 );
and ( n35081 , n33959 , n33990 );
or ( n35082 , n35079 , n35080 , n35081 );
and ( n35083 , n33920 , n33936 );
and ( n35084 , n33936 , n33952 );
and ( n35085 , n33920 , n33952 );
or ( n35086 , n35083 , n35084 , n35085 );
and ( n35087 , n33903 , n33907 );
and ( n35088 , n33907 , n33913 );
and ( n35089 , n33903 , n33913 );
or ( n35090 , n35087 , n35088 , n35089 );
and ( n35091 , n33924 , n33929 );
and ( n35092 , n33929 , n33935 );
and ( n35093 , n33924 , n33935 );
or ( n35094 , n35091 , n35092 , n35093 );
xor ( n35095 , n35090 , n35094 );
and ( n35096 , n33909 , n33910 );
and ( n35097 , n33910 , n33912 );
and ( n35098 , n33909 , n33912 );
or ( n35099 , n35096 , n35097 , n35098 );
and ( n35100 , n33925 , n33926 );
and ( n35101 , n33926 , n33928 );
and ( n35102 , n33925 , n33928 );
or ( n35103 , n35100 , n35101 , n35102 );
xor ( n35104 , n35099 , n35103 );
and ( n35105 , n21216 , n1551 );
and ( n35106 , n22186 , n1424 );
xor ( n35107 , n35105 , n35106 );
and ( n35108 , n22892 , n1254 );
xor ( n35109 , n35107 , n35108 );
xor ( n35110 , n35104 , n35109 );
xor ( n35111 , n35095 , n35110 );
xor ( n35112 , n35086 , n35111 );
and ( n35113 , n33941 , n33945 );
and ( n35114 , n33945 , n33951 );
and ( n35115 , n33941 , n33951 );
or ( n35116 , n35113 , n35114 , n35115 );
and ( n35117 , n33931 , n33932 );
and ( n35118 , n33932 , n33934 );
and ( n35119 , n33931 , n33934 );
or ( n35120 , n35117 , n35118 , n35119 );
and ( n35121 , n18144 , n2100 );
and ( n35122 , n19324 , n1882 );
xor ( n35123 , n35121 , n35122 );
and ( n35124 , n20233 , n1738 );
xor ( n35125 , n35123 , n35124 );
xor ( n35126 , n35120 , n35125 );
and ( n35127 , n15758 , n2739 );
and ( n35128 , n16637 , n2544 );
xor ( n35129 , n35127 , n35128 );
and ( n35130 , n17512 , n2298 );
xor ( n35131 , n35129 , n35130 );
xor ( n35132 , n35126 , n35131 );
xor ( n35133 , n35116 , n35132 );
and ( n35134 , n33947 , n33948 );
and ( n35135 , n33948 , n33950 );
and ( n35136 , n33947 , n33950 );
or ( n35137 , n35134 , n35135 , n35136 );
and ( n35138 , n33978 , n33979 );
and ( n35139 , n33979 , n33981 );
and ( n35140 , n33978 , n33981 );
or ( n35141 , n35138 , n35139 , n35140 );
xor ( n35142 , n35137 , n35141 );
and ( n35143 , n13322 , n3495 );
and ( n35144 , n14118 , n3271 );
xor ( n35145 , n35143 , n35144 );
and ( n35146 , n14938 , n2981 );
xor ( n35147 , n35145 , n35146 );
xor ( n35148 , n35142 , n35147 );
xor ( n35149 , n35133 , n35148 );
xor ( n35150 , n35112 , n35149 );
xor ( n35151 , n35082 , n35150 );
and ( n35152 , n33968 , n33972 );
and ( n35153 , n33972 , n33989 );
and ( n35154 , n33968 , n33989 );
or ( n35155 , n35152 , n35153 , n35154 );
and ( n35156 , n34015 , n34030 );
and ( n35157 , n34030 , n34047 );
and ( n35158 , n34015 , n34047 );
or ( n35159 , n35156 , n35157 , n35158 );
xor ( n35160 , n35155 , n35159 );
and ( n35161 , n33977 , n33982 );
and ( n35162 , n33982 , n33988 );
and ( n35163 , n33977 , n33988 );
or ( n35164 , n35161 , n35162 , n35163 );
and ( n35165 , n34019 , n34023 );
and ( n35166 , n34023 , n34029 );
and ( n35167 , n34019 , n34029 );
or ( n35168 , n35165 , n35166 , n35167 );
xor ( n35169 , n35164 , n35168 );
and ( n35170 , n33984 , n33985 );
and ( n35171 , n33985 , n33987 );
and ( n35172 , n33984 , n33987 );
or ( n35173 , n35170 , n35171 , n35172 );
and ( n35174 , n11015 , n4403 );
and ( n35175 , n11769 , n4102 );
xor ( n35176 , n35174 , n35175 );
and ( n35177 , n12320 , n3749 );
xor ( n35178 , n35176 , n35177 );
xor ( n35179 , n35173 , n35178 );
and ( n35180 , n8718 , n5408 );
and ( n35181 , n9400 , n5103 );
xor ( n35182 , n35180 , n35181 );
and ( n35183 , n10291 , n4730 );
xor ( n35184 , n35182 , n35183 );
xor ( n35185 , n35179 , n35184 );
xor ( n35186 , n35169 , n35185 );
xor ( n35187 , n35160 , n35186 );
xor ( n35188 , n35151 , n35187 );
xor ( n35189 , n35078 , n35188 );
xor ( n35190 , n35069 , n35189 );
and ( n35191 , n34081 , n34128 );
and ( n35192 , n34128 , n34202 );
and ( n35193 , n34081 , n34202 );
or ( n35194 , n35191 , n35192 , n35193 );
and ( n35195 , n34011 , n34048 );
and ( n35196 , n34048 , n34074 );
and ( n35197 , n34011 , n34074 );
or ( n35198 , n35195 , n35196 , n35197 );
and ( n35199 , n34085 , n34089 );
and ( n35200 , n34089 , n34127 );
and ( n35201 , n34085 , n34127 );
or ( n35202 , n35199 , n35200 , n35201 );
xor ( n35203 , n35198 , n35202 );
and ( n35204 , n34053 , n34057 );
and ( n35205 , n34057 , n34073 );
and ( n35206 , n34053 , n34073 );
or ( n35207 , n35204 , n35205 , n35206 );
and ( n35208 , n34035 , n34040 );
and ( n35209 , n34040 , n34046 );
and ( n35210 , n34035 , n34046 );
or ( n35211 , n35208 , n35209 , n35210 );
and ( n35212 , n34025 , n34026 );
and ( n35213 , n34026 , n34028 );
and ( n35214 , n34025 , n34028 );
or ( n35215 , n35212 , n35213 , n35214 );
and ( n35216 , n34036 , n34037 );
and ( n35217 , n34037 , n34039 );
and ( n35218 , n34036 , n34039 );
or ( n35219 , n35216 , n35217 , n35218 );
xor ( n35220 , n35215 , n35219 );
and ( n35221 , n7385 , n6504 );
and ( n35222 , n7808 , n6132 );
xor ( n35223 , n35221 , n35222 );
and ( n35224 , n8079 , n5765 );
xor ( n35225 , n35223 , n35224 );
xor ( n35226 , n35220 , n35225 );
xor ( n35227 , n35211 , n35226 );
and ( n35228 , n34042 , n34043 );
and ( n35229 , n34043 , n34045 );
and ( n35230 , n34042 , n34045 );
or ( n35231 , n35228 , n35229 , n35230 );
and ( n35232 , n6187 , n7662 );
and ( n35233 , n6569 , n7310 );
xor ( n35234 , n35232 , n35233 );
buf ( n35235 , n6816 );
xor ( n35236 , n35234 , n35235 );
xor ( n35237 , n35231 , n35236 );
and ( n35238 , n4959 , n9348 );
and ( n35239 , n5459 , n8669 );
xor ( n35240 , n35238 , n35239 );
and ( n35241 , n5819 , n8243 );
xor ( n35242 , n35240 , n35241 );
xor ( n35243 , n35237 , n35242 );
xor ( n35244 , n35227 , n35243 );
xor ( n35245 , n35207 , n35244 );
and ( n35246 , n34062 , n34066 );
and ( n35247 , n34066 , n34072 );
and ( n35248 , n34062 , n34072 );
or ( n35249 , n35246 , n35247 , n35248 );
and ( n35250 , n34098 , n34103 );
and ( n35251 , n34103 , n34109 );
and ( n35252 , n34098 , n34109 );
or ( n35253 , n35250 , n35251 , n35252 );
xor ( n35254 , n35249 , n35253 );
and ( n35255 , n34068 , n34069 );
and ( n35256 , n34069 , n34071 );
and ( n35257 , n34068 , n34071 );
or ( n35258 , n35255 , n35256 , n35257 );
and ( n35259 , n34099 , n34100 );
and ( n35260 , n34100 , n34102 );
and ( n35261 , n34099 , n34102 );
or ( n35262 , n35259 , n35260 , n35261 );
xor ( n35263 , n35258 , n35262 );
and ( n35264 , n4132 , n11718 );
and ( n35265 , n4438 , n10977 );
xor ( n35266 , n35264 , n35265 );
and ( n35267 , n4766 , n10239 );
xor ( n35268 , n35266 , n35267 );
xor ( n35269 , n35263 , n35268 );
xor ( n35270 , n35254 , n35269 );
xor ( n35271 , n35245 , n35270 );
xor ( n35272 , n35203 , n35271 );
xor ( n35273 , n35194 , n35272 );
and ( n35274 , n34133 , n34159 );
and ( n35275 , n34159 , n34201 );
and ( n35276 , n34133 , n34201 );
or ( n35277 , n35274 , n35275 , n35276 );
and ( n35278 , n34094 , n34110 );
and ( n35279 , n34110 , n34126 );
and ( n35280 , n34094 , n34126 );
or ( n35281 , n35278 , n35279 , n35280 );
and ( n35282 , n34137 , n34141 );
and ( n35283 , n34141 , n34158 );
and ( n35284 , n34137 , n34158 );
or ( n35285 , n35282 , n35283 , n35284 );
xor ( n35286 , n35281 , n35285 );
and ( n35287 , n34115 , n34119 );
and ( n35288 , n34119 , n34125 );
and ( n35289 , n34115 , n34125 );
or ( n35290 , n35287 , n35288 , n35289 );
and ( n35291 , n34105 , n34106 );
and ( n35292 , n34106 , n34108 );
and ( n35293 , n34105 , n34108 );
or ( n35294 , n35291 , n35292 , n35293 );
and ( n35295 , n3182 , n14044 );
and ( n35296 , n3545 , n13256 );
xor ( n35297 , n35295 , n35296 );
and ( n35298 , n3801 , n12531 );
xor ( n35299 , n35297 , n35298 );
xor ( n35300 , n35294 , n35299 );
and ( n35301 , n2462 , n16550 );
and ( n35302 , n2779 , n15691 );
xor ( n35303 , n35301 , n35302 );
and ( n35304 , n3024 , n14838 );
xor ( n35305 , n35303 , n35304 );
xor ( n35306 , n35300 , n35305 );
xor ( n35307 , n35290 , n35306 );
and ( n35308 , n34121 , n34122 );
and ( n35309 , n34122 , n34124 );
and ( n35310 , n34121 , n34124 );
or ( n35311 , n35308 , n35309 , n35310 );
and ( n35312 , n34147 , n34148 );
and ( n35313 , n34148 , n34150 );
and ( n35314 , n34147 , n34150 );
or ( n35315 , n35312 , n35313 , n35314 );
xor ( n35316 , n35311 , n35315 );
and ( n35317 , n1933 , n19222 );
and ( n35318 , n2120 , n18407 );
xor ( n35319 , n35317 , n35318 );
and ( n35320 , n2324 , n17422 );
xor ( n35321 , n35319 , n35320 );
xor ( n35322 , n35316 , n35321 );
xor ( n35323 , n35307 , n35322 );
xor ( n35324 , n35286 , n35323 );
xor ( n35325 , n35277 , n35324 );
and ( n35326 , n34164 , n34179 );
and ( n35327 , n34179 , n34200 );
and ( n35328 , n34164 , n34200 );
or ( n35329 , n35326 , n35327 , n35328 );
and ( n35330 , n34146 , n34151 );
and ( n35331 , n34151 , n34157 );
and ( n35332 , n34146 , n34157 );
or ( n35333 , n35330 , n35331 , n35332 );
and ( n35334 , n34168 , n34172 );
and ( n35335 , n34172 , n34178 );
and ( n35336 , n34168 , n34178 );
or ( n35337 , n35334 , n35335 , n35336 );
xor ( n35338 , n35333 , n35337 );
and ( n35339 , n34153 , n34154 );
and ( n35340 , n34154 , n34156 );
and ( n35341 , n34153 , n34156 );
or ( n35342 , n35339 , n35340 , n35341 );
and ( n35343 , n1383 , n22065 );
and ( n35344 , n1580 , n20976 );
xor ( n35345 , n35343 , n35344 );
and ( n35346 , n1694 , n20156 );
xor ( n35347 , n35345 , n35346 );
xor ( n35348 , n35342 , n35347 );
and ( n35349 , n1047 , n25163 );
and ( n35350 , n1164 , n24137 );
xor ( n35351 , n35349 , n35350 );
and ( n35352 , n1287 , n23075 );
xor ( n35353 , n35351 , n35352 );
xor ( n35354 , n35348 , n35353 );
xor ( n35355 , n35338 , n35354 );
xor ( n35356 , n35329 , n35355 );
and ( n35357 , n34184 , n34189 );
and ( n35358 , n34189 , n34199 );
and ( n35359 , n34184 , n34199 );
or ( n35360 , n35357 , n35358 , n35359 );
and ( n35361 , n34174 , n34175 );
and ( n35362 , n34175 , n34177 );
and ( n35363 , n34174 , n34177 );
or ( n35364 , n35361 , n35362 , n35363 );
and ( n35365 , n34185 , n34186 );
and ( n35366 , n34186 , n34188 );
and ( n35367 , n34185 , n34188 );
or ( n35368 , n35365 , n35366 , n35367 );
xor ( n35369 , n35364 , n35368 );
and ( n35370 , n783 , n28406 );
and ( n35371 , n856 , n27296 );
xor ( n35372 , n35370 , n35371 );
and ( n35373 , n925 , n26216 );
xor ( n35374 , n35372 , n35373 );
xor ( n35375 , n35369 , n35374 );
xor ( n35376 , n35360 , n35375 );
and ( n35377 , n34195 , n34196 );
and ( n35378 , n34196 , n34198 );
and ( n35379 , n34195 , n34198 );
or ( n35380 , n35377 , n35378 , n35379 );
and ( n35381 , n632 , n31761 );
and ( n35382 , n671 , n30629 );
xor ( n35383 , n35381 , n35382 );
and ( n35384 , n715 , n29508 );
xor ( n35385 , n35383 , n35384 );
xor ( n35386 , n35380 , n35385 );
not ( n35387 , n608 );
and ( n35388 , n34193 , n608 );
nor ( n35389 , n35387 , n35388 );
and ( n35390 , n611 , n32999 );
xor ( n35391 , n35389 , n35390 );
xor ( n35392 , n35386 , n35391 );
xor ( n35393 , n35376 , n35392 );
xor ( n35394 , n35356 , n35393 );
xor ( n35395 , n35325 , n35394 );
xor ( n35396 , n35273 , n35395 );
xor ( n35397 , n35190 , n35396 );
xor ( n35398 , n35065 , n35397 );
xor ( n35399 , n34983 , n35398 );
xor ( n35400 , n34974 , n35399 );
and ( n35401 , n33772 , n33777 );
and ( n35402 , n33777 , n34207 );
and ( n35403 , n33772 , n34207 );
or ( n35404 , n35401 , n35402 , n35403 );
xor ( n35405 , n35400 , n35404 );
and ( n35406 , n34208 , n34211 );
xor ( n35407 , n35405 , n35406 );
buf ( n35408 , n35407 );
buf ( n35409 , n35408 );
not ( n35410 , n35409 );
nor ( n35411 , n35410 , n8739 );
xor ( n35412 , n34966 , n35411 );
and ( n35413 , n33768 , n34216 );
and ( n35414 , n34217 , n34220 );
or ( n35415 , n35413 , n35414 );
xor ( n35416 , n35412 , n35415 );
buf ( n35417 , n35416 );
buf ( n35418 , n35417 );
not ( n35419 , n35418 );
buf ( n35420 , n563 );
not ( n35421 , n35420 );
nor ( n35422 , n35419 , n35421 );
xor ( n35423 , n34598 , n35422 );
xor ( n35424 , n34232 , n34595 );
nor ( n35425 , n34224 , n35421 );
and ( n35426 , n35424 , n35425 );
xor ( n35427 , n35424 , n35425 );
xor ( n35428 , n34236 , n34593 );
nor ( n35429 , n33033 , n35421 );
and ( n35430 , n35428 , n35429 );
xor ( n35431 , n35428 , n35429 );
xor ( n35432 , n34240 , n34591 );
nor ( n35433 , n31867 , n35421 );
and ( n35434 , n35432 , n35433 );
xor ( n35435 , n35432 , n35433 );
xor ( n35436 , n34244 , n34589 );
nor ( n35437 , n30725 , n35421 );
and ( n35438 , n35436 , n35437 );
xor ( n35439 , n35436 , n35437 );
xor ( n35440 , n34248 , n34587 );
nor ( n35441 , n29596 , n35421 );
and ( n35442 , n35440 , n35441 );
xor ( n35443 , n35440 , n35441 );
xor ( n35444 , n34252 , n34585 );
nor ( n35445 , n28487 , n35421 );
and ( n35446 , n35444 , n35445 );
xor ( n35447 , n35444 , n35445 );
xor ( n35448 , n34256 , n34583 );
nor ( n35449 , n27397 , n35421 );
and ( n35450 , n35448 , n35449 );
xor ( n35451 , n35448 , n35449 );
xor ( n35452 , n34260 , n34581 );
nor ( n35453 , n26326 , n35421 );
and ( n35454 , n35452 , n35453 );
xor ( n35455 , n35452 , n35453 );
xor ( n35456 , n34264 , n34579 );
nor ( n35457 , n25272 , n35421 );
and ( n35458 , n35456 , n35457 );
xor ( n35459 , n35456 , n35457 );
xor ( n35460 , n34268 , n34577 );
nor ( n35461 , n24242 , n35421 );
and ( n35462 , n35460 , n35461 );
xor ( n35463 , n35460 , n35461 );
xor ( n35464 , n34272 , n34575 );
nor ( n35465 , n23225 , n35421 );
and ( n35466 , n35464 , n35465 );
xor ( n35467 , n35464 , n35465 );
xor ( n35468 , n34276 , n34573 );
nor ( n35469 , n22231 , n35421 );
and ( n35470 , n35468 , n35469 );
xor ( n35471 , n35468 , n35469 );
xor ( n35472 , n34280 , n34571 );
nor ( n35473 , n21258 , n35421 );
and ( n35474 , n35472 , n35473 );
xor ( n35475 , n35472 , n35473 );
xor ( n35476 , n34284 , n34569 );
nor ( n35477 , n20303 , n35421 );
and ( n35478 , n35476 , n35477 );
xor ( n35479 , n35476 , n35477 );
xor ( n35480 , n34288 , n34567 );
nor ( n35481 , n19365 , n35421 );
and ( n35482 , n35480 , n35481 );
xor ( n35483 , n35480 , n35481 );
xor ( n35484 , n34292 , n34565 );
nor ( n35485 , n18448 , n35421 );
and ( n35486 , n35484 , n35485 );
xor ( n35487 , n35484 , n35485 );
xor ( n35488 , n34296 , n34563 );
nor ( n35489 , n17548 , n35421 );
and ( n35490 , n35488 , n35489 );
xor ( n35491 , n35488 , n35489 );
xor ( n35492 , n34300 , n34561 );
nor ( n35493 , n16669 , n35421 );
and ( n35494 , n35492 , n35493 );
xor ( n35495 , n35492 , n35493 );
xor ( n35496 , n34304 , n34559 );
nor ( n35497 , n15809 , n35421 );
and ( n35498 , n35496 , n35497 );
xor ( n35499 , n35496 , n35497 );
xor ( n35500 , n34308 , n34557 );
nor ( n35501 , n14968 , n35421 );
and ( n35502 , n35500 , n35501 );
xor ( n35503 , n35500 , n35501 );
xor ( n35504 , n34312 , n34555 );
nor ( n35505 , n14147 , n35421 );
and ( n35506 , n35504 , n35505 );
xor ( n35507 , n35504 , n35505 );
xor ( n35508 , n34316 , n34553 );
nor ( n35509 , n13349 , n35421 );
and ( n35510 , n35508 , n35509 );
xor ( n35511 , n35508 , n35509 );
xor ( n35512 , n34320 , n34551 );
nor ( n35513 , n12564 , n35421 );
and ( n35514 , n35512 , n35513 );
xor ( n35515 , n35512 , n35513 );
xor ( n35516 , n34324 , n34549 );
nor ( n35517 , n11799 , n35421 );
and ( n35518 , n35516 , n35517 );
xor ( n35519 , n35516 , n35517 );
xor ( n35520 , n34328 , n34547 );
nor ( n35521 , n11050 , n35421 );
and ( n35522 , n35520 , n35521 );
xor ( n35523 , n35520 , n35521 );
xor ( n35524 , n34332 , n34545 );
nor ( n35525 , n10321 , n35421 );
and ( n35526 , n35524 , n35525 );
xor ( n35527 , n35524 , n35525 );
xor ( n35528 , n34336 , n34543 );
nor ( n35529 , n9429 , n35421 );
and ( n35530 , n35528 , n35529 );
xor ( n35531 , n35528 , n35529 );
xor ( n35532 , n34340 , n34541 );
nor ( n35533 , n8949 , n35421 );
and ( n35534 , n35532 , n35533 );
xor ( n35535 , n35532 , n35533 );
xor ( n35536 , n34344 , n34539 );
nor ( n35537 , n9437 , n35421 );
and ( n35538 , n35536 , n35537 );
xor ( n35539 , n35536 , n35537 );
xor ( n35540 , n34348 , n34537 );
nor ( n35541 , n9446 , n35421 );
and ( n35542 , n35540 , n35541 );
xor ( n35543 , n35540 , n35541 );
xor ( n35544 , n34352 , n34535 );
nor ( n35545 , n9455 , n35421 );
and ( n35546 , n35544 , n35545 );
xor ( n35547 , n35544 , n35545 );
xor ( n35548 , n34356 , n34533 );
nor ( n35549 , n9464 , n35421 );
and ( n35550 , n35548 , n35549 );
xor ( n35551 , n35548 , n35549 );
xor ( n35552 , n34360 , n34531 );
nor ( n35553 , n9473 , n35421 );
and ( n35554 , n35552 , n35553 );
xor ( n35555 , n35552 , n35553 );
xor ( n35556 , n34364 , n34529 );
nor ( n35557 , n9482 , n35421 );
and ( n35558 , n35556 , n35557 );
xor ( n35559 , n35556 , n35557 );
xor ( n35560 , n34368 , n34527 );
nor ( n35561 , n9491 , n35421 );
and ( n35562 , n35560 , n35561 );
xor ( n35563 , n35560 , n35561 );
xor ( n35564 , n34372 , n34525 );
nor ( n35565 , n9500 , n35421 );
and ( n35566 , n35564 , n35565 );
xor ( n35567 , n35564 , n35565 );
xor ( n35568 , n34376 , n34523 );
nor ( n35569 , n9509 , n35421 );
and ( n35570 , n35568 , n35569 );
xor ( n35571 , n35568 , n35569 );
xor ( n35572 , n34380 , n34521 );
nor ( n35573 , n9518 , n35421 );
and ( n35574 , n35572 , n35573 );
xor ( n35575 , n35572 , n35573 );
xor ( n35576 , n34384 , n34519 );
nor ( n35577 , n9527 , n35421 );
and ( n35578 , n35576 , n35577 );
xor ( n35579 , n35576 , n35577 );
xor ( n35580 , n34388 , n34517 );
nor ( n35581 , n9536 , n35421 );
and ( n35582 , n35580 , n35581 );
xor ( n35583 , n35580 , n35581 );
xor ( n35584 , n34392 , n34515 );
nor ( n35585 , n9545 , n35421 );
and ( n35586 , n35584 , n35585 );
xor ( n35587 , n35584 , n35585 );
xor ( n35588 , n34396 , n34513 );
nor ( n35589 , n9554 , n35421 );
and ( n35590 , n35588 , n35589 );
xor ( n35591 , n35588 , n35589 );
xor ( n35592 , n34400 , n34511 );
nor ( n35593 , n9563 , n35421 );
and ( n35594 , n35592 , n35593 );
xor ( n35595 , n35592 , n35593 );
xor ( n35596 , n34404 , n34509 );
nor ( n35597 , n9572 , n35421 );
and ( n35598 , n35596 , n35597 );
xor ( n35599 , n35596 , n35597 );
xor ( n35600 , n34408 , n34507 );
nor ( n35601 , n9581 , n35421 );
and ( n35602 , n35600 , n35601 );
xor ( n35603 , n35600 , n35601 );
xor ( n35604 , n34412 , n34505 );
nor ( n35605 , n9590 , n35421 );
and ( n35606 , n35604 , n35605 );
xor ( n35607 , n35604 , n35605 );
xor ( n35608 , n34416 , n34503 );
nor ( n35609 , n9599 , n35421 );
and ( n35610 , n35608 , n35609 );
xor ( n35611 , n35608 , n35609 );
xor ( n35612 , n34420 , n34501 );
nor ( n35613 , n9608 , n35421 );
and ( n35614 , n35612 , n35613 );
xor ( n35615 , n35612 , n35613 );
xor ( n35616 , n34424 , n34499 );
nor ( n35617 , n9617 , n35421 );
and ( n35618 , n35616 , n35617 );
xor ( n35619 , n35616 , n35617 );
xor ( n35620 , n34428 , n34497 );
nor ( n35621 , n9626 , n35421 );
and ( n35622 , n35620 , n35621 );
xor ( n35623 , n35620 , n35621 );
xor ( n35624 , n34432 , n34495 );
nor ( n35625 , n9635 , n35421 );
and ( n35626 , n35624 , n35625 );
xor ( n35627 , n35624 , n35625 );
xor ( n35628 , n34436 , n34493 );
nor ( n35629 , n9644 , n35421 );
and ( n35630 , n35628 , n35629 );
xor ( n35631 , n35628 , n35629 );
xor ( n35632 , n34440 , n34491 );
nor ( n35633 , n9653 , n35421 );
and ( n35634 , n35632 , n35633 );
xor ( n35635 , n35632 , n35633 );
xor ( n35636 , n34444 , n34489 );
nor ( n35637 , n9662 , n35421 );
and ( n35638 , n35636 , n35637 );
xor ( n35639 , n35636 , n35637 );
xor ( n35640 , n34448 , n34487 );
nor ( n35641 , n9671 , n35421 );
and ( n35642 , n35640 , n35641 );
xor ( n35643 , n35640 , n35641 );
xor ( n35644 , n34452 , n34485 );
nor ( n35645 , n9680 , n35421 );
and ( n35646 , n35644 , n35645 );
xor ( n35647 , n35644 , n35645 );
xor ( n35648 , n34456 , n34483 );
nor ( n35649 , n9689 , n35421 );
and ( n35650 , n35648 , n35649 );
xor ( n35651 , n35648 , n35649 );
xor ( n35652 , n34460 , n34481 );
nor ( n35653 , n9698 , n35421 );
and ( n35654 , n35652 , n35653 );
xor ( n35655 , n35652 , n35653 );
xor ( n35656 , n34464 , n34479 );
nor ( n35657 , n9707 , n35421 );
and ( n35658 , n35656 , n35657 );
xor ( n35659 , n35656 , n35657 );
xor ( n35660 , n34468 , n34477 );
nor ( n35661 , n9716 , n35421 );
and ( n35662 , n35660 , n35661 );
xor ( n35663 , n35660 , n35661 );
xor ( n35664 , n34472 , n34475 );
nor ( n35665 , n9725 , n35421 );
and ( n35666 , n35664 , n35665 );
xor ( n35667 , n35664 , n35665 );
xor ( n35668 , n34473 , n34474 );
nor ( n35669 , n9734 , n35421 );
and ( n35670 , n35668 , n35669 );
xor ( n35671 , n35668 , n35669 );
nor ( n35672 , n9752 , n34226 );
nor ( n35673 , n9743 , n35421 );
and ( n35674 , n35672 , n35673 );
and ( n35675 , n35671 , n35674 );
or ( n35676 , n35670 , n35675 );
and ( n35677 , n35667 , n35676 );
or ( n35678 , n35666 , n35677 );
and ( n35679 , n35663 , n35678 );
or ( n35680 , n35662 , n35679 );
and ( n35681 , n35659 , n35680 );
or ( n35682 , n35658 , n35681 );
and ( n35683 , n35655 , n35682 );
or ( n35684 , n35654 , n35683 );
and ( n35685 , n35651 , n35684 );
or ( n35686 , n35650 , n35685 );
and ( n35687 , n35647 , n35686 );
or ( n35688 , n35646 , n35687 );
and ( n35689 , n35643 , n35688 );
or ( n35690 , n35642 , n35689 );
and ( n35691 , n35639 , n35690 );
or ( n35692 , n35638 , n35691 );
and ( n35693 , n35635 , n35692 );
or ( n35694 , n35634 , n35693 );
and ( n35695 , n35631 , n35694 );
or ( n35696 , n35630 , n35695 );
and ( n35697 , n35627 , n35696 );
or ( n35698 , n35626 , n35697 );
and ( n35699 , n35623 , n35698 );
or ( n35700 , n35622 , n35699 );
and ( n35701 , n35619 , n35700 );
or ( n35702 , n35618 , n35701 );
and ( n35703 , n35615 , n35702 );
or ( n35704 , n35614 , n35703 );
and ( n35705 , n35611 , n35704 );
or ( n35706 , n35610 , n35705 );
and ( n35707 , n35607 , n35706 );
or ( n35708 , n35606 , n35707 );
and ( n35709 , n35603 , n35708 );
or ( n35710 , n35602 , n35709 );
and ( n35711 , n35599 , n35710 );
or ( n35712 , n35598 , n35711 );
and ( n35713 , n35595 , n35712 );
or ( n35714 , n35594 , n35713 );
and ( n35715 , n35591 , n35714 );
or ( n35716 , n35590 , n35715 );
and ( n35717 , n35587 , n35716 );
or ( n35718 , n35586 , n35717 );
and ( n35719 , n35583 , n35718 );
or ( n35720 , n35582 , n35719 );
and ( n35721 , n35579 , n35720 );
or ( n35722 , n35578 , n35721 );
and ( n35723 , n35575 , n35722 );
or ( n35724 , n35574 , n35723 );
and ( n35725 , n35571 , n35724 );
or ( n35726 , n35570 , n35725 );
and ( n35727 , n35567 , n35726 );
or ( n35728 , n35566 , n35727 );
and ( n35729 , n35563 , n35728 );
or ( n35730 , n35562 , n35729 );
and ( n35731 , n35559 , n35730 );
or ( n35732 , n35558 , n35731 );
and ( n35733 , n35555 , n35732 );
or ( n35734 , n35554 , n35733 );
and ( n35735 , n35551 , n35734 );
or ( n35736 , n35550 , n35735 );
and ( n35737 , n35547 , n35736 );
or ( n35738 , n35546 , n35737 );
and ( n35739 , n35543 , n35738 );
or ( n35740 , n35542 , n35739 );
and ( n35741 , n35539 , n35740 );
or ( n35742 , n35538 , n35741 );
and ( n35743 , n35535 , n35742 );
or ( n35744 , n35534 , n35743 );
and ( n35745 , n35531 , n35744 );
or ( n35746 , n35530 , n35745 );
and ( n35747 , n35527 , n35746 );
or ( n35748 , n35526 , n35747 );
and ( n35749 , n35523 , n35748 );
or ( n35750 , n35522 , n35749 );
and ( n35751 , n35519 , n35750 );
or ( n35752 , n35518 , n35751 );
and ( n35753 , n35515 , n35752 );
or ( n35754 , n35514 , n35753 );
and ( n35755 , n35511 , n35754 );
or ( n35756 , n35510 , n35755 );
and ( n35757 , n35507 , n35756 );
or ( n35758 , n35506 , n35757 );
and ( n35759 , n35503 , n35758 );
or ( n35760 , n35502 , n35759 );
and ( n35761 , n35499 , n35760 );
or ( n35762 , n35498 , n35761 );
and ( n35763 , n35495 , n35762 );
or ( n35764 , n35494 , n35763 );
and ( n35765 , n35491 , n35764 );
or ( n35766 , n35490 , n35765 );
and ( n35767 , n35487 , n35766 );
or ( n35768 , n35486 , n35767 );
and ( n35769 , n35483 , n35768 );
or ( n35770 , n35482 , n35769 );
and ( n35771 , n35479 , n35770 );
or ( n35772 , n35478 , n35771 );
and ( n35773 , n35475 , n35772 );
or ( n35774 , n35474 , n35773 );
and ( n35775 , n35471 , n35774 );
or ( n35776 , n35470 , n35775 );
and ( n35777 , n35467 , n35776 );
or ( n35778 , n35466 , n35777 );
and ( n35779 , n35463 , n35778 );
or ( n35780 , n35462 , n35779 );
and ( n35781 , n35459 , n35780 );
or ( n35782 , n35458 , n35781 );
and ( n35783 , n35455 , n35782 );
or ( n35784 , n35454 , n35783 );
and ( n35785 , n35451 , n35784 );
or ( n35786 , n35450 , n35785 );
and ( n35787 , n35447 , n35786 );
or ( n35788 , n35446 , n35787 );
and ( n35789 , n35443 , n35788 );
or ( n35790 , n35442 , n35789 );
and ( n35791 , n35439 , n35790 );
or ( n35792 , n35438 , n35791 );
and ( n35793 , n35435 , n35792 );
or ( n35794 , n35434 , n35793 );
and ( n35795 , n35431 , n35794 );
or ( n35796 , n35430 , n35795 );
and ( n35797 , n35427 , n35796 );
or ( n35798 , n35426 , n35797 );
xor ( n35799 , n35423 , n35798 );
and ( n35800 , n33403 , n621 );
nor ( n35801 , n622 , n35800 );
nor ( n35802 , n646 , n32231 );
xor ( n35803 , n35801 , n35802 );
buf ( n35804 , n35803 );
nor ( n35805 , n684 , n31083 );
xor ( n35806 , n35804 , n35805 );
and ( n35807 , n34601 , n34602 );
and ( n35808 , n34603 , n34605 );
or ( n35809 , n35807 , n35808 );
xor ( n35810 , n35806 , n35809 );
nor ( n35811 , n733 , n29948 );
xor ( n35812 , n35810 , n35811 );
and ( n35813 , n34606 , n34607 );
and ( n35814 , n34608 , n34611 );
or ( n35815 , n35813 , n35814 );
xor ( n35816 , n35812 , n35815 );
nor ( n35817 , n796 , n28833 );
xor ( n35818 , n35816 , n35817 );
and ( n35819 , n34612 , n34613 );
and ( n35820 , n34614 , n34617 );
or ( n35821 , n35819 , n35820 );
xor ( n35822 , n35818 , n35821 );
nor ( n35823 , n868 , n27737 );
xor ( n35824 , n35822 , n35823 );
and ( n35825 , n34618 , n34619 );
and ( n35826 , n34620 , n34623 );
or ( n35827 , n35825 , n35826 );
xor ( n35828 , n35824 , n35827 );
nor ( n35829 , n958 , n26660 );
xor ( n35830 , n35828 , n35829 );
and ( n35831 , n34624 , n34625 );
and ( n35832 , n34626 , n34629 );
or ( n35833 , n35831 , n35832 );
xor ( n35834 , n35830 , n35833 );
nor ( n35835 , n1062 , n25600 );
xor ( n35836 , n35834 , n35835 );
and ( n35837 , n34630 , n34631 );
and ( n35838 , n34632 , n34635 );
or ( n35839 , n35837 , n35838 );
xor ( n35840 , n35836 , n35839 );
nor ( n35841 , n1176 , n24564 );
xor ( n35842 , n35840 , n35841 );
and ( n35843 , n34636 , n34637 );
and ( n35844 , n34638 , n34641 );
or ( n35845 , n35843 , n35844 );
xor ( n35846 , n35842 , n35845 );
nor ( n35847 , n1303 , n23541 );
xor ( n35848 , n35846 , n35847 );
and ( n35849 , n34642 , n34643 );
and ( n35850 , n34644 , n34647 );
or ( n35851 , n35849 , n35850 );
xor ( n35852 , n35848 , n35851 );
nor ( n35853 , n1445 , n22541 );
xor ( n35854 , n35852 , n35853 );
and ( n35855 , n34648 , n34649 );
and ( n35856 , n34650 , n34653 );
or ( n35857 , n35855 , n35856 );
xor ( n35858 , n35854 , n35857 );
nor ( n35859 , n1598 , n21562 );
xor ( n35860 , n35858 , n35859 );
and ( n35861 , n34654 , n34655 );
and ( n35862 , n34656 , n34659 );
or ( n35863 , n35861 , n35862 );
xor ( n35864 , n35860 , n35863 );
nor ( n35865 , n1766 , n20601 );
xor ( n35866 , n35864 , n35865 );
and ( n35867 , n34660 , n34661 );
and ( n35868 , n34662 , n34665 );
or ( n35869 , n35867 , n35868 );
xor ( n35870 , n35866 , n35869 );
nor ( n35871 , n1945 , n19657 );
xor ( n35872 , n35870 , n35871 );
and ( n35873 , n34666 , n34667 );
and ( n35874 , n34668 , n34671 );
or ( n35875 , n35873 , n35874 );
xor ( n35876 , n35872 , n35875 );
nor ( n35877 , n2137 , n18734 );
xor ( n35878 , n35876 , n35877 );
and ( n35879 , n34672 , n34673 );
and ( n35880 , n34674 , n34677 );
or ( n35881 , n35879 , n35880 );
xor ( n35882 , n35878 , n35881 );
nor ( n35883 , n2343 , n17828 );
xor ( n35884 , n35882 , n35883 );
and ( n35885 , n34678 , n34679 );
and ( n35886 , n34680 , n34683 );
or ( n35887 , n35885 , n35886 );
xor ( n35888 , n35884 , n35887 );
nor ( n35889 , n2566 , n16943 );
xor ( n35890 , n35888 , n35889 );
and ( n35891 , n34684 , n34685 );
and ( n35892 , n34686 , n34689 );
or ( n35893 , n35891 , n35892 );
xor ( n35894 , n35890 , n35893 );
nor ( n35895 , n2797 , n16077 );
xor ( n35896 , n35894 , n35895 );
and ( n35897 , n34690 , n34691 );
and ( n35898 , n34692 , n34695 );
or ( n35899 , n35897 , n35898 );
xor ( n35900 , n35896 , n35899 );
nor ( n35901 , n3043 , n15230 );
xor ( n35902 , n35900 , n35901 );
and ( n35903 , n34696 , n34697 );
and ( n35904 , n34698 , n34701 );
or ( n35905 , n35903 , n35904 );
xor ( n35906 , n35902 , n35905 );
nor ( n35907 , n3300 , n14403 );
xor ( n35908 , n35906 , n35907 );
and ( n35909 , n34702 , n34703 );
and ( n35910 , n34704 , n34707 );
or ( n35911 , n35909 , n35910 );
xor ( n35912 , n35908 , n35911 );
nor ( n35913 , n3570 , n13599 );
xor ( n35914 , n35912 , n35913 );
and ( n35915 , n34708 , n34709 );
and ( n35916 , n34710 , n34713 );
or ( n35917 , n35915 , n35916 );
xor ( n35918 , n35914 , n35917 );
nor ( n35919 , n3853 , n12808 );
xor ( n35920 , n35918 , n35919 );
and ( n35921 , n34714 , n34715 );
and ( n35922 , n34716 , n34719 );
or ( n35923 , n35921 , n35922 );
xor ( n35924 , n35920 , n35923 );
nor ( n35925 , n4151 , n12037 );
xor ( n35926 , n35924 , n35925 );
and ( n35927 , n34720 , n34721 );
and ( n35928 , n34722 , n34725 );
or ( n35929 , n35927 , n35928 );
xor ( n35930 , n35926 , n35929 );
nor ( n35931 , n4458 , n11282 );
xor ( n35932 , n35930 , n35931 );
and ( n35933 , n34726 , n34727 );
and ( n35934 , n34728 , n34731 );
or ( n35935 , n35933 , n35934 );
xor ( n35936 , n35932 , n35935 );
nor ( n35937 , n4786 , n10547 );
xor ( n35938 , n35936 , n35937 );
and ( n35939 , n34732 , n34733 );
and ( n35940 , n34734 , n34737 );
or ( n35941 , n35939 , n35940 );
xor ( n35942 , n35938 , n35941 );
nor ( n35943 , n5126 , n9829 );
xor ( n35944 , n35942 , n35943 );
and ( n35945 , n34738 , n34739 );
and ( n35946 , n34740 , n34743 );
or ( n35947 , n35945 , n35946 );
xor ( n35948 , n35944 , n35947 );
nor ( n35949 , n5477 , n8955 );
xor ( n35950 , n35948 , n35949 );
and ( n35951 , n34744 , n34745 );
and ( n35952 , n34746 , n34749 );
or ( n35953 , n35951 , n35952 );
xor ( n35954 , n35950 , n35953 );
nor ( n35955 , n5838 , n603 );
xor ( n35956 , n35954 , n35955 );
and ( n35957 , n34750 , n34751 );
and ( n35958 , n34752 , n34755 );
or ( n35959 , n35957 , n35958 );
xor ( n35960 , n35956 , n35959 );
nor ( n35961 , n6212 , n652 );
xor ( n35962 , n35960 , n35961 );
and ( n35963 , n34756 , n34757 );
and ( n35964 , n34758 , n34761 );
or ( n35965 , n35963 , n35964 );
xor ( n35966 , n35962 , n35965 );
nor ( n35967 , n6596 , n624 );
xor ( n35968 , n35966 , n35967 );
and ( n35969 , n34762 , n34763 );
and ( n35970 , n34764 , n34767 );
or ( n35971 , n35969 , n35970 );
xor ( n35972 , n35968 , n35971 );
nor ( n35973 , n6997 , n648 );
xor ( n35974 , n35972 , n35973 );
and ( n35975 , n34768 , n34769 );
and ( n35976 , n34770 , n34773 );
or ( n35977 , n35975 , n35976 );
xor ( n35978 , n35974 , n35977 );
nor ( n35979 , n7413 , n686 );
xor ( n35980 , n35978 , n35979 );
and ( n35981 , n34774 , n34775 );
and ( n35982 , n34776 , n34779 );
or ( n35983 , n35981 , n35982 );
xor ( n35984 , n35980 , n35983 );
nor ( n35985 , n7841 , n735 );
xor ( n35986 , n35984 , n35985 );
and ( n35987 , n34780 , n34781 );
and ( n35988 , n34782 , n34785 );
or ( n35989 , n35987 , n35988 );
xor ( n35990 , n35986 , n35989 );
nor ( n35991 , n8281 , n798 );
xor ( n35992 , n35990 , n35991 );
and ( n35993 , n34786 , n34787 );
and ( n35994 , n34788 , n34791 );
or ( n35995 , n35993 , n35994 );
xor ( n35996 , n35992 , n35995 );
nor ( n35997 , n8737 , n870 );
xor ( n35998 , n35996 , n35997 );
and ( n35999 , n34792 , n34793 );
and ( n36000 , n34794 , n34797 );
or ( n36001 , n35999 , n36000 );
xor ( n36002 , n35998 , n36001 );
nor ( n36003 , n9420 , n960 );
xor ( n36004 , n36002 , n36003 );
and ( n36005 , n34798 , n34799 );
and ( n36006 , n34800 , n34803 );
or ( n36007 , n36005 , n36006 );
xor ( n36008 , n36004 , n36007 );
nor ( n36009 , n10312 , n1064 );
xor ( n36010 , n36008 , n36009 );
and ( n36011 , n34804 , n34805 );
and ( n36012 , n34806 , n34809 );
or ( n36013 , n36011 , n36012 );
xor ( n36014 , n36010 , n36013 );
nor ( n36015 , n11041 , n1178 );
xor ( n36016 , n36014 , n36015 );
and ( n36017 , n34810 , n34811 );
and ( n36018 , n34812 , n34815 );
or ( n36019 , n36017 , n36018 );
xor ( n36020 , n36016 , n36019 );
nor ( n36021 , n11790 , n1305 );
xor ( n36022 , n36020 , n36021 );
and ( n36023 , n34816 , n34817 );
and ( n36024 , n34818 , n34821 );
or ( n36025 , n36023 , n36024 );
xor ( n36026 , n36022 , n36025 );
nor ( n36027 , n12555 , n1447 );
xor ( n36028 , n36026 , n36027 );
and ( n36029 , n34822 , n34823 );
and ( n36030 , n34824 , n34827 );
or ( n36031 , n36029 , n36030 );
xor ( n36032 , n36028 , n36031 );
nor ( n36033 , n13340 , n1600 );
xor ( n36034 , n36032 , n36033 );
and ( n36035 , n34828 , n34829 );
and ( n36036 , n34830 , n34833 );
or ( n36037 , n36035 , n36036 );
xor ( n36038 , n36034 , n36037 );
nor ( n36039 , n14138 , n1768 );
xor ( n36040 , n36038 , n36039 );
and ( n36041 , n34834 , n34835 );
and ( n36042 , n34836 , n34839 );
or ( n36043 , n36041 , n36042 );
xor ( n36044 , n36040 , n36043 );
nor ( n36045 , n14959 , n1947 );
xor ( n36046 , n36044 , n36045 );
and ( n36047 , n34840 , n34841 );
and ( n36048 , n34842 , n34845 );
or ( n36049 , n36047 , n36048 );
xor ( n36050 , n36046 , n36049 );
nor ( n36051 , n15800 , n2139 );
xor ( n36052 , n36050 , n36051 );
and ( n36053 , n34846 , n34847 );
and ( n36054 , n34848 , n34851 );
or ( n36055 , n36053 , n36054 );
xor ( n36056 , n36052 , n36055 );
nor ( n36057 , n16660 , n2345 );
xor ( n36058 , n36056 , n36057 );
and ( n36059 , n34852 , n34853 );
and ( n36060 , n34854 , n34857 );
or ( n36061 , n36059 , n36060 );
xor ( n36062 , n36058 , n36061 );
nor ( n36063 , n17539 , n2568 );
xor ( n36064 , n36062 , n36063 );
and ( n36065 , n34858 , n34859 );
and ( n36066 , n34860 , n34863 );
or ( n36067 , n36065 , n36066 );
xor ( n36068 , n36064 , n36067 );
nor ( n36069 , n18439 , n2799 );
xor ( n36070 , n36068 , n36069 );
and ( n36071 , n34864 , n34865 );
and ( n36072 , n34866 , n34869 );
or ( n36073 , n36071 , n36072 );
xor ( n36074 , n36070 , n36073 );
nor ( n36075 , n19356 , n3045 );
xor ( n36076 , n36074 , n36075 );
and ( n36077 , n34870 , n34871 );
and ( n36078 , n34872 , n34875 );
or ( n36079 , n36077 , n36078 );
xor ( n36080 , n36076 , n36079 );
nor ( n36081 , n20294 , n3302 );
xor ( n36082 , n36080 , n36081 );
and ( n36083 , n34876 , n34877 );
and ( n36084 , n34878 , n34881 );
or ( n36085 , n36083 , n36084 );
xor ( n36086 , n36082 , n36085 );
nor ( n36087 , n21249 , n3572 );
xor ( n36088 , n36086 , n36087 );
and ( n36089 , n34882 , n34883 );
and ( n36090 , n34884 , n34887 );
or ( n36091 , n36089 , n36090 );
xor ( n36092 , n36088 , n36091 );
nor ( n36093 , n22222 , n3855 );
xor ( n36094 , n36092 , n36093 );
and ( n36095 , n34888 , n34889 );
and ( n36096 , n34890 , n34893 );
or ( n36097 , n36095 , n36096 );
xor ( n36098 , n36094 , n36097 );
nor ( n36099 , n23216 , n4153 );
xor ( n36100 , n36098 , n36099 );
and ( n36101 , n34894 , n34895 );
and ( n36102 , n34896 , n34899 );
or ( n36103 , n36101 , n36102 );
xor ( n36104 , n36100 , n36103 );
nor ( n36105 , n24233 , n4460 );
xor ( n36106 , n36104 , n36105 );
and ( n36107 , n34900 , n34901 );
and ( n36108 , n34902 , n34905 );
or ( n36109 , n36107 , n36108 );
xor ( n36110 , n36106 , n36109 );
nor ( n36111 , n25263 , n4788 );
xor ( n36112 , n36110 , n36111 );
and ( n36113 , n34906 , n34907 );
and ( n36114 , n34908 , n34911 );
or ( n36115 , n36113 , n36114 );
xor ( n36116 , n36112 , n36115 );
nor ( n36117 , n26317 , n5128 );
xor ( n36118 , n36116 , n36117 );
and ( n36119 , n34912 , n34913 );
and ( n36120 , n34914 , n34917 );
or ( n36121 , n36119 , n36120 );
xor ( n36122 , n36118 , n36121 );
nor ( n36123 , n27388 , n5479 );
xor ( n36124 , n36122 , n36123 );
and ( n36125 , n34918 , n34919 );
and ( n36126 , n34920 , n34923 );
or ( n36127 , n36125 , n36126 );
xor ( n36128 , n36124 , n36127 );
nor ( n36129 , n28478 , n5840 );
xor ( n36130 , n36128 , n36129 );
and ( n36131 , n34924 , n34925 );
and ( n36132 , n34926 , n34929 );
or ( n36133 , n36131 , n36132 );
xor ( n36134 , n36130 , n36133 );
nor ( n36135 , n29587 , n6214 );
xor ( n36136 , n36134 , n36135 );
and ( n36137 , n34930 , n34931 );
and ( n36138 , n34932 , n34935 );
or ( n36139 , n36137 , n36138 );
xor ( n36140 , n36136 , n36139 );
nor ( n36141 , n30716 , n6598 );
xor ( n36142 , n36140 , n36141 );
and ( n36143 , n34936 , n34937 );
and ( n36144 , n34938 , n34941 );
or ( n36145 , n36143 , n36144 );
xor ( n36146 , n36142 , n36145 );
nor ( n36147 , n31858 , n6999 );
xor ( n36148 , n36146 , n36147 );
and ( n36149 , n34942 , n34943 );
and ( n36150 , n34944 , n34947 );
or ( n36151 , n36149 , n36150 );
xor ( n36152 , n36148 , n36151 );
nor ( n36153 , n33024 , n7415 );
xor ( n36154 , n36152 , n36153 );
and ( n36155 , n34948 , n34949 );
and ( n36156 , n34950 , n34953 );
or ( n36157 , n36155 , n36156 );
xor ( n36158 , n36154 , n36157 );
nor ( n36159 , n34215 , n7843 );
xor ( n36160 , n36158 , n36159 );
and ( n36161 , n34954 , n34955 );
and ( n36162 , n34956 , n34959 );
or ( n36163 , n36161 , n36162 );
xor ( n36164 , n36160 , n36163 );
nor ( n36165 , n35410 , n8283 );
xor ( n36166 , n36164 , n36165 );
and ( n36167 , n34960 , n34961 );
and ( n36168 , n34962 , n34965 );
or ( n36169 , n36167 , n36168 );
xor ( n36170 , n36166 , n36169 );
and ( n36171 , n34978 , n34982 );
and ( n36172 , n34982 , n35398 );
and ( n36173 , n34978 , n35398 );
or ( n36174 , n36171 , n36172 , n36173 );
and ( n36175 , n33774 , n606 );
not ( n36176 , n606 );
nor ( n36177 , n36175 , n36176 );
xor ( n36178 , n36174 , n36177 );
and ( n36179 , n34991 , n34995 );
and ( n36180 , n34995 , n35063 );
and ( n36181 , n34991 , n35063 );
or ( n36182 , n36179 , n36180 , n36181 );
and ( n36183 , n34987 , n35064 );
and ( n36184 , n35064 , n35397 );
and ( n36185 , n34987 , n35397 );
or ( n36186 , n36183 , n36184 , n36185 );
xor ( n36187 , n36182 , n36186 );
and ( n36188 , n35069 , n35189 );
and ( n36189 , n35189 , n35396 );
and ( n36190 , n35069 , n35396 );
or ( n36191 , n36188 , n36189 , n36190 );
and ( n36192 , n35000 , n35004 );
and ( n36193 , n35004 , n35062 );
and ( n36194 , n35000 , n35062 );
or ( n36195 , n36192 , n36193 , n36194 );
and ( n36196 , n35073 , n35077 );
and ( n36197 , n35077 , n35188 );
and ( n36198 , n35073 , n35188 );
or ( n36199 , n36196 , n36197 , n36198 );
xor ( n36200 , n36195 , n36199 );
and ( n36201 , n35031 , n35035 );
and ( n36202 , n35035 , n35041 );
and ( n36203 , n35031 , n35041 );
or ( n36204 , n36201 , n36202 , n36203 );
and ( n36205 , n35009 , n35013 );
and ( n36206 , n35013 , n35061 );
and ( n36207 , n35009 , n35061 );
or ( n36208 , n36205 , n36206 , n36207 );
xor ( n36209 , n36204 , n36208 );
and ( n36210 , n35018 , n35022 );
and ( n36211 , n35022 , n35060 );
and ( n36212 , n35018 , n35060 );
or ( n36213 , n36210 , n36211 , n36212 );
and ( n36214 , n35086 , n35111 );
and ( n36215 , n35111 , n35149 );
and ( n36216 , n35086 , n35149 );
or ( n36217 , n36214 , n36215 , n36216 );
xor ( n36218 , n36213 , n36217 );
and ( n36219 , n35027 , n35042 );
and ( n36220 , n35042 , n35059 );
and ( n36221 , n35027 , n35059 );
or ( n36222 , n36219 , n36220 , n36221 );
and ( n36223 , n35090 , n35094 );
and ( n36224 , n35094 , n35110 );
and ( n36225 , n35090 , n35110 );
or ( n36226 , n36223 , n36224 , n36225 );
xor ( n36227 , n36222 , n36226 );
and ( n36228 , n35047 , n35052 );
and ( n36229 , n35052 , n35058 );
and ( n36230 , n35047 , n35058 );
or ( n36231 , n36228 , n36229 , n36230 );
and ( n36232 , n35037 , n35038 );
and ( n36233 , n35038 , n35040 );
and ( n36234 , n35037 , n35040 );
or ( n36235 , n36232 , n36233 , n36234 );
and ( n36236 , n35048 , n35049 );
and ( n36237 , n35049 , n35051 );
and ( n36238 , n35048 , n35051 );
or ( n36239 , n36236 , n36237 , n36238 );
xor ( n36240 , n36235 , n36239 );
and ( n36241 , n30695 , n719 );
and ( n36242 , n31836 , n663 );
xor ( n36243 , n36241 , n36242 );
and ( n36244 , n32649 , n635 );
xor ( n36245 , n36243 , n36244 );
xor ( n36246 , n36240 , n36245 );
xor ( n36247 , n36231 , n36246 );
and ( n36248 , n35054 , n35055 );
and ( n36249 , n35055 , n35057 );
and ( n36250 , n35054 , n35057 );
or ( n36251 , n36248 , n36249 , n36250 );
and ( n36252 , n27361 , n940 );
and ( n36253 , n28456 , n840 );
xor ( n36254 , n36252 , n36253 );
and ( n36255 , n29559 , n771 );
xor ( n36256 , n36254 , n36255 );
xor ( n36257 , n36251 , n36256 );
and ( n36258 , n24214 , n1254 );
and ( n36259 , n25243 , n1134 );
xor ( n36260 , n36258 , n36259 );
and ( n36261 , n26296 , n1034 );
xor ( n36262 , n36260 , n36261 );
xor ( n36263 , n36257 , n36262 );
xor ( n36264 , n36247 , n36263 );
xor ( n36265 , n36227 , n36264 );
xor ( n36266 , n36218 , n36265 );
xor ( n36267 , n36209 , n36266 );
xor ( n36268 , n36200 , n36267 );
xor ( n36269 , n36191 , n36268 );
and ( n36270 , n35194 , n35272 );
and ( n36271 , n35272 , n35395 );
and ( n36272 , n35194 , n35395 );
or ( n36273 , n36270 , n36271 , n36272 );
and ( n36274 , n35082 , n35150 );
and ( n36275 , n35150 , n35187 );
and ( n36276 , n35082 , n35187 );
or ( n36277 , n36274 , n36275 , n36276 );
and ( n36278 , n35198 , n35202 );
and ( n36279 , n35202 , n35271 );
and ( n36280 , n35198 , n35271 );
or ( n36281 , n36278 , n36279 , n36280 );
xor ( n36282 , n36277 , n36281 );
and ( n36283 , n35155 , n35159 );
and ( n36284 , n35159 , n35186 );
and ( n36285 , n35155 , n35186 );
or ( n36286 , n36283 , n36284 , n36285 );
and ( n36287 , n35116 , n35132 );
and ( n36288 , n35132 , n35148 );
and ( n36289 , n35116 , n35148 );
or ( n36290 , n36287 , n36288 , n36289 );
and ( n36291 , n35099 , n35103 );
and ( n36292 , n35103 , n35109 );
and ( n36293 , n35099 , n35109 );
or ( n36294 , n36291 , n36292 , n36293 );
and ( n36295 , n35120 , n35125 );
and ( n36296 , n35125 , n35131 );
and ( n36297 , n35120 , n35131 );
or ( n36298 , n36295 , n36296 , n36297 );
xor ( n36299 , n36294 , n36298 );
and ( n36300 , n35105 , n35106 );
and ( n36301 , n35106 , n35108 );
and ( n36302 , n35105 , n35108 );
or ( n36303 , n36300 , n36301 , n36302 );
and ( n36304 , n35121 , n35122 );
and ( n36305 , n35122 , n35124 );
and ( n36306 , n35121 , n35124 );
or ( n36307 , n36304 , n36305 , n36306 );
xor ( n36308 , n36303 , n36307 );
and ( n36309 , n21216 , n1738 );
and ( n36310 , n22186 , n1551 );
xor ( n36311 , n36309 , n36310 );
and ( n36312 , n22892 , n1424 );
xor ( n36313 , n36311 , n36312 );
xor ( n36314 , n36308 , n36313 );
xor ( n36315 , n36299 , n36314 );
xor ( n36316 , n36290 , n36315 );
and ( n36317 , n35137 , n35141 );
and ( n36318 , n35141 , n35147 );
and ( n36319 , n35137 , n35147 );
or ( n36320 , n36317 , n36318 , n36319 );
and ( n36321 , n35127 , n35128 );
and ( n36322 , n35128 , n35130 );
and ( n36323 , n35127 , n35130 );
or ( n36324 , n36321 , n36322 , n36323 );
and ( n36325 , n18144 , n2298 );
and ( n36326 , n19324 , n2100 );
xor ( n36327 , n36325 , n36326 );
and ( n36328 , n20233 , n1882 );
xor ( n36329 , n36327 , n36328 );
xor ( n36330 , n36324 , n36329 );
and ( n36331 , n15758 , n2981 );
and ( n36332 , n16637 , n2739 );
xor ( n36333 , n36331 , n36332 );
and ( n36334 , n17512 , n2544 );
xor ( n36335 , n36333 , n36334 );
xor ( n36336 , n36330 , n36335 );
xor ( n36337 , n36320 , n36336 );
and ( n36338 , n35143 , n35144 );
and ( n36339 , n35144 , n35146 );
and ( n36340 , n35143 , n35146 );
or ( n36341 , n36338 , n36339 , n36340 );
and ( n36342 , n35174 , n35175 );
and ( n36343 , n35175 , n35177 );
and ( n36344 , n35174 , n35177 );
or ( n36345 , n36342 , n36343 , n36344 );
xor ( n36346 , n36341 , n36345 );
and ( n36347 , n13322 , n3749 );
and ( n36348 , n14118 , n3495 );
xor ( n36349 , n36347 , n36348 );
and ( n36350 , n14938 , n3271 );
xor ( n36351 , n36349 , n36350 );
xor ( n36352 , n36346 , n36351 );
xor ( n36353 , n36337 , n36352 );
xor ( n36354 , n36316 , n36353 );
xor ( n36355 , n36286 , n36354 );
and ( n36356 , n35164 , n35168 );
and ( n36357 , n35168 , n35185 );
and ( n36358 , n35164 , n35185 );
or ( n36359 , n36356 , n36357 , n36358 );
and ( n36360 , n35211 , n35226 );
and ( n36361 , n35226 , n35243 );
and ( n36362 , n35211 , n35243 );
or ( n36363 , n36360 , n36361 , n36362 );
xor ( n36364 , n36359 , n36363 );
and ( n36365 , n35173 , n35178 );
and ( n36366 , n35178 , n35184 );
and ( n36367 , n35173 , n35184 );
or ( n36368 , n36365 , n36366 , n36367 );
and ( n36369 , n35215 , n35219 );
and ( n36370 , n35219 , n35225 );
and ( n36371 , n35215 , n35225 );
or ( n36372 , n36369 , n36370 , n36371 );
xor ( n36373 , n36368 , n36372 );
and ( n36374 , n35180 , n35181 );
and ( n36375 , n35181 , n35183 );
and ( n36376 , n35180 , n35183 );
or ( n36377 , n36374 , n36375 , n36376 );
and ( n36378 , n11015 , n4730 );
and ( n36379 , n11769 , n4403 );
xor ( n36380 , n36378 , n36379 );
and ( n36381 , n12320 , n4102 );
xor ( n36382 , n36380 , n36381 );
xor ( n36383 , n36377 , n36382 );
and ( n36384 , n8718 , n5765 );
and ( n36385 , n9400 , n5408 );
xor ( n36386 , n36384 , n36385 );
and ( n36387 , n10291 , n5103 );
xor ( n36388 , n36386 , n36387 );
xor ( n36389 , n36383 , n36388 );
xor ( n36390 , n36373 , n36389 );
xor ( n36391 , n36364 , n36390 );
xor ( n36392 , n36355 , n36391 );
xor ( n36393 , n36282 , n36392 );
xor ( n36394 , n36273 , n36393 );
and ( n36395 , n35277 , n35324 );
and ( n36396 , n35324 , n35394 );
and ( n36397 , n35277 , n35394 );
or ( n36398 , n36395 , n36396 , n36397 );
and ( n36399 , n35207 , n35244 );
and ( n36400 , n35244 , n35270 );
and ( n36401 , n35207 , n35270 );
or ( n36402 , n36399 , n36400 , n36401 );
and ( n36403 , n35281 , n35285 );
and ( n36404 , n35285 , n35323 );
and ( n36405 , n35281 , n35323 );
or ( n36406 , n36403 , n36404 , n36405 );
xor ( n36407 , n36402 , n36406 );
and ( n36408 , n35249 , n35253 );
and ( n36409 , n35253 , n35269 );
and ( n36410 , n35249 , n35269 );
or ( n36411 , n36408 , n36409 , n36410 );
and ( n36412 , n35231 , n35236 );
and ( n36413 , n35236 , n35242 );
and ( n36414 , n35231 , n35242 );
or ( n36415 , n36412 , n36413 , n36414 );
and ( n36416 , n35221 , n35222 );
and ( n36417 , n35222 , n35224 );
and ( n36418 , n35221 , n35224 );
or ( n36419 , n36416 , n36417 , n36418 );
and ( n36420 , n35232 , n35233 );
and ( n36421 , n35233 , n35235 );
and ( n36422 , n35232 , n35235 );
or ( n36423 , n36420 , n36421 , n36422 );
xor ( n36424 , n36419 , n36423 );
and ( n36425 , n7385 , n6971 );
and ( n36426 , n7808 , n6504 );
xor ( n36427 , n36425 , n36426 );
and ( n36428 , n8079 , n6132 );
xor ( n36429 , n36427 , n36428 );
xor ( n36430 , n36424 , n36429 );
xor ( n36431 , n36415 , n36430 );
and ( n36432 , n35238 , n35239 );
and ( n36433 , n35239 , n35241 );
and ( n36434 , n35238 , n35241 );
or ( n36435 , n36432 , n36433 , n36434 );
and ( n36436 , n6187 , n8243 );
and ( n36437 , n6569 , n7662 );
xor ( n36438 , n36436 , n36437 );
and ( n36439 , n6816 , n7310 );
xor ( n36440 , n36438 , n36439 );
xor ( n36441 , n36435 , n36440 );
and ( n36442 , n4959 , n10239 );
and ( n36443 , n5459 , n9348 );
xor ( n36444 , n36442 , n36443 );
and ( n36445 , n5819 , n8669 );
xor ( n36446 , n36444 , n36445 );
xor ( n36447 , n36441 , n36446 );
xor ( n36448 , n36431 , n36447 );
xor ( n36449 , n36411 , n36448 );
and ( n36450 , n35258 , n35262 );
and ( n36451 , n35262 , n35268 );
and ( n36452 , n35258 , n35268 );
or ( n36453 , n36450 , n36451 , n36452 );
and ( n36454 , n35294 , n35299 );
and ( n36455 , n35299 , n35305 );
and ( n36456 , n35294 , n35305 );
or ( n36457 , n36454 , n36455 , n36456 );
xor ( n36458 , n36453 , n36457 );
and ( n36459 , n35264 , n35265 );
and ( n36460 , n35265 , n35267 );
and ( n36461 , n35264 , n35267 );
or ( n36462 , n36459 , n36460 , n36461 );
and ( n36463 , n35295 , n35296 );
and ( n36464 , n35296 , n35298 );
and ( n36465 , n35295 , n35298 );
or ( n36466 , n36463 , n36464 , n36465 );
xor ( n36467 , n36462 , n36466 );
and ( n36468 , n4132 , n12531 );
and ( n36469 , n4438 , n11718 );
xor ( n36470 , n36468 , n36469 );
and ( n36471 , n4766 , n10977 );
xor ( n36472 , n36470 , n36471 );
xor ( n36473 , n36467 , n36472 );
xor ( n36474 , n36458 , n36473 );
xor ( n36475 , n36449 , n36474 );
xor ( n36476 , n36407 , n36475 );
xor ( n36477 , n36398 , n36476 );
and ( n36478 , n35329 , n35355 );
and ( n36479 , n35355 , n35393 );
and ( n36480 , n35329 , n35393 );
or ( n36481 , n36478 , n36479 , n36480 );
and ( n36482 , n35290 , n35306 );
and ( n36483 , n35306 , n35322 );
and ( n36484 , n35290 , n35322 );
or ( n36485 , n36482 , n36483 , n36484 );
and ( n36486 , n35333 , n35337 );
and ( n36487 , n35337 , n35354 );
and ( n36488 , n35333 , n35354 );
or ( n36489 , n36486 , n36487 , n36488 );
xor ( n36490 , n36485 , n36489 );
and ( n36491 , n35311 , n35315 );
and ( n36492 , n35315 , n35321 );
and ( n36493 , n35311 , n35321 );
or ( n36494 , n36491 , n36492 , n36493 );
and ( n36495 , n35301 , n35302 );
and ( n36496 , n35302 , n35304 );
and ( n36497 , n35301 , n35304 );
or ( n36498 , n36495 , n36496 , n36497 );
and ( n36499 , n3182 , n14838 );
and ( n36500 , n3545 , n14044 );
xor ( n36501 , n36499 , n36500 );
and ( n36502 , n3801 , n13256 );
xor ( n36503 , n36501 , n36502 );
xor ( n36504 , n36498 , n36503 );
and ( n36505 , n2462 , n17422 );
and ( n36506 , n2779 , n16550 );
xor ( n36507 , n36505 , n36506 );
and ( n36508 , n3024 , n15691 );
xor ( n36509 , n36507 , n36508 );
xor ( n36510 , n36504 , n36509 );
xor ( n36511 , n36494 , n36510 );
and ( n36512 , n35317 , n35318 );
and ( n36513 , n35318 , n35320 );
and ( n36514 , n35317 , n35320 );
or ( n36515 , n36512 , n36513 , n36514 );
and ( n36516 , n35343 , n35344 );
and ( n36517 , n35344 , n35346 );
and ( n36518 , n35343 , n35346 );
or ( n36519 , n36516 , n36517 , n36518 );
xor ( n36520 , n36515 , n36519 );
and ( n36521 , n1933 , n20156 );
and ( n36522 , n2120 , n19222 );
xor ( n36523 , n36521 , n36522 );
and ( n36524 , n2324 , n18407 );
xor ( n36525 , n36523 , n36524 );
xor ( n36526 , n36520 , n36525 );
xor ( n36527 , n36511 , n36526 );
xor ( n36528 , n36490 , n36527 );
xor ( n36529 , n36481 , n36528 );
and ( n36530 , n35360 , n35375 );
and ( n36531 , n35375 , n35392 );
and ( n36532 , n35360 , n35392 );
or ( n36533 , n36530 , n36531 , n36532 );
and ( n36534 , n35342 , n35347 );
and ( n36535 , n35347 , n35353 );
and ( n36536 , n35342 , n35353 );
or ( n36537 , n36534 , n36535 , n36536 );
and ( n36538 , n35364 , n35368 );
and ( n36539 , n35368 , n35374 );
and ( n36540 , n35364 , n35374 );
or ( n36541 , n36538 , n36539 , n36540 );
xor ( n36542 , n36537 , n36541 );
and ( n36543 , n35349 , n35350 );
and ( n36544 , n35350 , n35352 );
and ( n36545 , n35349 , n35352 );
or ( n36546 , n36543 , n36544 , n36545 );
and ( n36547 , n1383 , n23075 );
and ( n36548 , n1580 , n22065 );
xor ( n36549 , n36547 , n36548 );
and ( n36550 , n1694 , n20976 );
xor ( n36551 , n36549 , n36550 );
xor ( n36552 , n36546 , n36551 );
and ( n36553 , n1047 , n26216 );
and ( n36554 , n1164 , n25163 );
xor ( n36555 , n36553 , n36554 );
and ( n36556 , n1287 , n24137 );
xor ( n36557 , n36555 , n36556 );
xor ( n36558 , n36552 , n36557 );
xor ( n36559 , n36542 , n36558 );
xor ( n36560 , n36533 , n36559 );
and ( n36561 , n35380 , n35385 );
and ( n36562 , n35385 , n35391 );
and ( n36563 , n35380 , n35391 );
or ( n36564 , n36561 , n36562 , n36563 );
and ( n36565 , n35370 , n35371 );
and ( n36566 , n35371 , n35373 );
and ( n36567 , n35370 , n35373 );
or ( n36568 , n36565 , n36566 , n36567 );
and ( n36569 , n35381 , n35382 );
and ( n36570 , n35382 , n35384 );
and ( n36571 , n35381 , n35384 );
or ( n36572 , n36569 , n36570 , n36571 );
xor ( n36573 , n36568 , n36572 );
and ( n36574 , n783 , n29508 );
and ( n36575 , n856 , n28406 );
xor ( n36576 , n36574 , n36575 );
and ( n36577 , n925 , n27296 );
xor ( n36578 , n36576 , n36577 );
xor ( n36579 , n36573 , n36578 );
xor ( n36580 , n36564 , n36579 );
and ( n36581 , n35389 , n35390 );
not ( n36582 , n611 );
and ( n36583 , n34193 , n611 );
nor ( n36584 , n36582 , n36583 );
xor ( n36585 , n36581 , n36584 );
and ( n36586 , n632 , n32999 );
and ( n36587 , n671 , n31761 );
xor ( n36588 , n36586 , n36587 );
and ( n36589 , n715 , n30629 );
xor ( n36590 , n36588 , n36589 );
xor ( n36591 , n36585 , n36590 );
xor ( n36592 , n36580 , n36591 );
xor ( n36593 , n36560 , n36592 );
xor ( n36594 , n36529 , n36593 );
xor ( n36595 , n36477 , n36594 );
xor ( n36596 , n36394 , n36595 );
xor ( n36597 , n36269 , n36596 );
xor ( n36598 , n36187 , n36597 );
xor ( n36599 , n36178 , n36598 );
and ( n36600 , n34970 , n34973 );
and ( n36601 , n34973 , n35399 );
and ( n36602 , n34970 , n35399 );
or ( n36603 , n36600 , n36601 , n36602 );
xor ( n36604 , n36599 , n36603 );
and ( n36605 , n35400 , n35404 );
and ( n36606 , n35405 , n35406 );
or ( n36607 , n36605 , n36606 );
xor ( n36608 , n36604 , n36607 );
buf ( n36609 , n36608 );
buf ( n36610 , n36609 );
not ( n36611 , n36610 );
nor ( n36612 , n36611 , n8739 );
xor ( n36613 , n36170 , n36612 );
and ( n36614 , n34966 , n35411 );
and ( n36615 , n35412 , n35415 );
or ( n36616 , n36614 , n36615 );
xor ( n36617 , n36613 , n36616 );
buf ( n36618 , n36617 );
buf ( n36619 , n36618 );
not ( n36620 , n36619 );
buf ( n36621 , n564 );
not ( n36622 , n36621 );
nor ( n36623 , n36620 , n36622 );
xor ( n36624 , n35799 , n36623 );
xor ( n36625 , n35427 , n35796 );
nor ( n36626 , n35419 , n36622 );
and ( n36627 , n36625 , n36626 );
xor ( n36628 , n36625 , n36626 );
xor ( n36629 , n35431 , n35794 );
nor ( n36630 , n34224 , n36622 );
and ( n36631 , n36629 , n36630 );
xor ( n36632 , n36629 , n36630 );
xor ( n36633 , n35435 , n35792 );
nor ( n36634 , n33033 , n36622 );
and ( n36635 , n36633 , n36634 );
xor ( n36636 , n36633 , n36634 );
xor ( n36637 , n35439 , n35790 );
nor ( n36638 , n31867 , n36622 );
and ( n36639 , n36637 , n36638 );
xor ( n36640 , n36637 , n36638 );
xor ( n36641 , n35443 , n35788 );
nor ( n36642 , n30725 , n36622 );
and ( n36643 , n36641 , n36642 );
xor ( n36644 , n36641 , n36642 );
xor ( n36645 , n35447 , n35786 );
nor ( n36646 , n29596 , n36622 );
and ( n36647 , n36645 , n36646 );
xor ( n36648 , n36645 , n36646 );
xor ( n36649 , n35451 , n35784 );
nor ( n36650 , n28487 , n36622 );
and ( n36651 , n36649 , n36650 );
xor ( n36652 , n36649 , n36650 );
xor ( n36653 , n35455 , n35782 );
nor ( n36654 , n27397 , n36622 );
and ( n36655 , n36653 , n36654 );
xor ( n36656 , n36653 , n36654 );
xor ( n36657 , n35459 , n35780 );
nor ( n36658 , n26326 , n36622 );
and ( n36659 , n36657 , n36658 );
xor ( n36660 , n36657 , n36658 );
xor ( n36661 , n35463 , n35778 );
nor ( n36662 , n25272 , n36622 );
and ( n36663 , n36661 , n36662 );
xor ( n36664 , n36661 , n36662 );
xor ( n36665 , n35467 , n35776 );
nor ( n36666 , n24242 , n36622 );
and ( n36667 , n36665 , n36666 );
xor ( n36668 , n36665 , n36666 );
xor ( n36669 , n35471 , n35774 );
nor ( n36670 , n23225 , n36622 );
and ( n36671 , n36669 , n36670 );
xor ( n36672 , n36669 , n36670 );
xor ( n36673 , n35475 , n35772 );
nor ( n36674 , n22231 , n36622 );
and ( n36675 , n36673 , n36674 );
xor ( n36676 , n36673 , n36674 );
xor ( n36677 , n35479 , n35770 );
nor ( n36678 , n21258 , n36622 );
and ( n36679 , n36677 , n36678 );
xor ( n36680 , n36677 , n36678 );
xor ( n36681 , n35483 , n35768 );
nor ( n36682 , n20303 , n36622 );
and ( n36683 , n36681 , n36682 );
xor ( n36684 , n36681 , n36682 );
xor ( n36685 , n35487 , n35766 );
nor ( n36686 , n19365 , n36622 );
and ( n36687 , n36685 , n36686 );
xor ( n36688 , n36685 , n36686 );
xor ( n36689 , n35491 , n35764 );
nor ( n36690 , n18448 , n36622 );
and ( n36691 , n36689 , n36690 );
xor ( n36692 , n36689 , n36690 );
xor ( n36693 , n35495 , n35762 );
nor ( n36694 , n17548 , n36622 );
and ( n36695 , n36693 , n36694 );
xor ( n36696 , n36693 , n36694 );
xor ( n36697 , n35499 , n35760 );
nor ( n36698 , n16669 , n36622 );
and ( n36699 , n36697 , n36698 );
xor ( n36700 , n36697 , n36698 );
xor ( n36701 , n35503 , n35758 );
nor ( n36702 , n15809 , n36622 );
and ( n36703 , n36701 , n36702 );
xor ( n36704 , n36701 , n36702 );
xor ( n36705 , n35507 , n35756 );
nor ( n36706 , n14968 , n36622 );
and ( n36707 , n36705 , n36706 );
xor ( n36708 , n36705 , n36706 );
xor ( n36709 , n35511 , n35754 );
nor ( n36710 , n14147 , n36622 );
and ( n36711 , n36709 , n36710 );
xor ( n36712 , n36709 , n36710 );
xor ( n36713 , n35515 , n35752 );
nor ( n36714 , n13349 , n36622 );
and ( n36715 , n36713 , n36714 );
xor ( n36716 , n36713 , n36714 );
xor ( n36717 , n35519 , n35750 );
nor ( n36718 , n12564 , n36622 );
and ( n36719 , n36717 , n36718 );
xor ( n36720 , n36717 , n36718 );
xor ( n36721 , n35523 , n35748 );
nor ( n36722 , n11799 , n36622 );
and ( n36723 , n36721 , n36722 );
xor ( n36724 , n36721 , n36722 );
xor ( n36725 , n35527 , n35746 );
nor ( n36726 , n11050 , n36622 );
and ( n36727 , n36725 , n36726 );
xor ( n36728 , n36725 , n36726 );
xor ( n36729 , n35531 , n35744 );
nor ( n36730 , n10321 , n36622 );
and ( n36731 , n36729 , n36730 );
xor ( n36732 , n36729 , n36730 );
xor ( n36733 , n35535 , n35742 );
nor ( n36734 , n9429 , n36622 );
and ( n36735 , n36733 , n36734 );
xor ( n36736 , n36733 , n36734 );
xor ( n36737 , n35539 , n35740 );
nor ( n36738 , n8949 , n36622 );
and ( n36739 , n36737 , n36738 );
xor ( n36740 , n36737 , n36738 );
xor ( n36741 , n35543 , n35738 );
nor ( n36742 , n9437 , n36622 );
and ( n36743 , n36741 , n36742 );
xor ( n36744 , n36741 , n36742 );
xor ( n36745 , n35547 , n35736 );
nor ( n36746 , n9446 , n36622 );
and ( n36747 , n36745 , n36746 );
xor ( n36748 , n36745 , n36746 );
xor ( n36749 , n35551 , n35734 );
nor ( n36750 , n9455 , n36622 );
and ( n36751 , n36749 , n36750 );
xor ( n36752 , n36749 , n36750 );
xor ( n36753 , n35555 , n35732 );
nor ( n36754 , n9464 , n36622 );
and ( n36755 , n36753 , n36754 );
xor ( n36756 , n36753 , n36754 );
xor ( n36757 , n35559 , n35730 );
nor ( n36758 , n9473 , n36622 );
and ( n36759 , n36757 , n36758 );
xor ( n36760 , n36757 , n36758 );
xor ( n36761 , n35563 , n35728 );
nor ( n36762 , n9482 , n36622 );
and ( n36763 , n36761 , n36762 );
xor ( n36764 , n36761 , n36762 );
xor ( n36765 , n35567 , n35726 );
nor ( n36766 , n9491 , n36622 );
and ( n36767 , n36765 , n36766 );
xor ( n36768 , n36765 , n36766 );
xor ( n36769 , n35571 , n35724 );
nor ( n36770 , n9500 , n36622 );
and ( n36771 , n36769 , n36770 );
xor ( n36772 , n36769 , n36770 );
xor ( n36773 , n35575 , n35722 );
nor ( n36774 , n9509 , n36622 );
and ( n36775 , n36773 , n36774 );
xor ( n36776 , n36773 , n36774 );
xor ( n36777 , n35579 , n35720 );
nor ( n36778 , n9518 , n36622 );
and ( n36779 , n36777 , n36778 );
xor ( n36780 , n36777 , n36778 );
xor ( n36781 , n35583 , n35718 );
nor ( n36782 , n9527 , n36622 );
and ( n36783 , n36781 , n36782 );
xor ( n36784 , n36781 , n36782 );
xor ( n36785 , n35587 , n35716 );
nor ( n36786 , n9536 , n36622 );
and ( n36787 , n36785 , n36786 );
xor ( n36788 , n36785 , n36786 );
xor ( n36789 , n35591 , n35714 );
nor ( n36790 , n9545 , n36622 );
and ( n36791 , n36789 , n36790 );
xor ( n36792 , n36789 , n36790 );
xor ( n36793 , n35595 , n35712 );
nor ( n36794 , n9554 , n36622 );
and ( n36795 , n36793 , n36794 );
xor ( n36796 , n36793 , n36794 );
xor ( n36797 , n35599 , n35710 );
nor ( n36798 , n9563 , n36622 );
and ( n36799 , n36797 , n36798 );
xor ( n36800 , n36797 , n36798 );
xor ( n36801 , n35603 , n35708 );
nor ( n36802 , n9572 , n36622 );
and ( n36803 , n36801 , n36802 );
xor ( n36804 , n36801 , n36802 );
xor ( n36805 , n35607 , n35706 );
nor ( n36806 , n9581 , n36622 );
and ( n36807 , n36805 , n36806 );
xor ( n36808 , n36805 , n36806 );
xor ( n36809 , n35611 , n35704 );
nor ( n36810 , n9590 , n36622 );
and ( n36811 , n36809 , n36810 );
xor ( n36812 , n36809 , n36810 );
xor ( n36813 , n35615 , n35702 );
nor ( n36814 , n9599 , n36622 );
and ( n36815 , n36813 , n36814 );
xor ( n36816 , n36813 , n36814 );
xor ( n36817 , n35619 , n35700 );
nor ( n36818 , n9608 , n36622 );
and ( n36819 , n36817 , n36818 );
xor ( n36820 , n36817 , n36818 );
xor ( n36821 , n35623 , n35698 );
nor ( n36822 , n9617 , n36622 );
and ( n36823 , n36821 , n36822 );
xor ( n36824 , n36821 , n36822 );
xor ( n36825 , n35627 , n35696 );
nor ( n36826 , n9626 , n36622 );
and ( n36827 , n36825 , n36826 );
xor ( n36828 , n36825 , n36826 );
xor ( n36829 , n35631 , n35694 );
nor ( n36830 , n9635 , n36622 );
and ( n36831 , n36829 , n36830 );
xor ( n36832 , n36829 , n36830 );
xor ( n36833 , n35635 , n35692 );
nor ( n36834 , n9644 , n36622 );
and ( n36835 , n36833 , n36834 );
xor ( n36836 , n36833 , n36834 );
xor ( n36837 , n35639 , n35690 );
nor ( n36838 , n9653 , n36622 );
and ( n36839 , n36837 , n36838 );
xor ( n36840 , n36837 , n36838 );
xor ( n36841 , n35643 , n35688 );
nor ( n36842 , n9662 , n36622 );
and ( n36843 , n36841 , n36842 );
xor ( n36844 , n36841 , n36842 );
xor ( n36845 , n35647 , n35686 );
nor ( n36846 , n9671 , n36622 );
and ( n36847 , n36845 , n36846 );
xor ( n36848 , n36845 , n36846 );
xor ( n36849 , n35651 , n35684 );
nor ( n36850 , n9680 , n36622 );
and ( n36851 , n36849 , n36850 );
xor ( n36852 , n36849 , n36850 );
xor ( n36853 , n35655 , n35682 );
nor ( n36854 , n9689 , n36622 );
and ( n36855 , n36853 , n36854 );
xor ( n36856 , n36853 , n36854 );
xor ( n36857 , n35659 , n35680 );
nor ( n36858 , n9698 , n36622 );
and ( n36859 , n36857 , n36858 );
xor ( n36860 , n36857 , n36858 );
xor ( n36861 , n35663 , n35678 );
nor ( n36862 , n9707 , n36622 );
and ( n36863 , n36861 , n36862 );
xor ( n36864 , n36861 , n36862 );
xor ( n36865 , n35667 , n35676 );
nor ( n36866 , n9716 , n36622 );
and ( n36867 , n36865 , n36866 );
xor ( n36868 , n36865 , n36866 );
xor ( n36869 , n35671 , n35674 );
nor ( n36870 , n9725 , n36622 );
and ( n36871 , n36869 , n36870 );
xor ( n36872 , n36869 , n36870 );
xor ( n36873 , n35672 , n35673 );
nor ( n36874 , n9734 , n36622 );
and ( n36875 , n36873 , n36874 );
xor ( n36876 , n36873 , n36874 );
nor ( n36877 , n9752 , n35421 );
nor ( n36878 , n9743 , n36622 );
and ( n36879 , n36877 , n36878 );
and ( n36880 , n36876 , n36879 );
or ( n36881 , n36875 , n36880 );
and ( n36882 , n36872 , n36881 );
or ( n36883 , n36871 , n36882 );
and ( n36884 , n36868 , n36883 );
or ( n36885 , n36867 , n36884 );
and ( n36886 , n36864 , n36885 );
or ( n36887 , n36863 , n36886 );
and ( n36888 , n36860 , n36887 );
or ( n36889 , n36859 , n36888 );
and ( n36890 , n36856 , n36889 );
or ( n36891 , n36855 , n36890 );
and ( n36892 , n36852 , n36891 );
or ( n36893 , n36851 , n36892 );
and ( n36894 , n36848 , n36893 );
or ( n36895 , n36847 , n36894 );
and ( n36896 , n36844 , n36895 );
or ( n36897 , n36843 , n36896 );
and ( n36898 , n36840 , n36897 );
or ( n36899 , n36839 , n36898 );
and ( n36900 , n36836 , n36899 );
or ( n36901 , n36835 , n36900 );
and ( n36902 , n36832 , n36901 );
or ( n36903 , n36831 , n36902 );
and ( n36904 , n36828 , n36903 );
or ( n36905 , n36827 , n36904 );
and ( n36906 , n36824 , n36905 );
or ( n36907 , n36823 , n36906 );
and ( n36908 , n36820 , n36907 );
or ( n36909 , n36819 , n36908 );
and ( n36910 , n36816 , n36909 );
or ( n36911 , n36815 , n36910 );
and ( n36912 , n36812 , n36911 );
or ( n36913 , n36811 , n36912 );
and ( n36914 , n36808 , n36913 );
or ( n36915 , n36807 , n36914 );
and ( n36916 , n36804 , n36915 );
or ( n36917 , n36803 , n36916 );
and ( n36918 , n36800 , n36917 );
or ( n36919 , n36799 , n36918 );
and ( n36920 , n36796 , n36919 );
or ( n36921 , n36795 , n36920 );
and ( n36922 , n36792 , n36921 );
or ( n36923 , n36791 , n36922 );
and ( n36924 , n36788 , n36923 );
or ( n36925 , n36787 , n36924 );
and ( n36926 , n36784 , n36925 );
or ( n36927 , n36783 , n36926 );
and ( n36928 , n36780 , n36927 );
or ( n36929 , n36779 , n36928 );
and ( n36930 , n36776 , n36929 );
or ( n36931 , n36775 , n36930 );
and ( n36932 , n36772 , n36931 );
or ( n36933 , n36771 , n36932 );
and ( n36934 , n36768 , n36933 );
or ( n36935 , n36767 , n36934 );
and ( n36936 , n36764 , n36935 );
or ( n36937 , n36763 , n36936 );
and ( n36938 , n36760 , n36937 );
or ( n36939 , n36759 , n36938 );
and ( n36940 , n36756 , n36939 );
or ( n36941 , n36755 , n36940 );
and ( n36942 , n36752 , n36941 );
or ( n36943 , n36751 , n36942 );
and ( n36944 , n36748 , n36943 );
or ( n36945 , n36747 , n36944 );
and ( n36946 , n36744 , n36945 );
or ( n36947 , n36743 , n36946 );
and ( n36948 , n36740 , n36947 );
or ( n36949 , n36739 , n36948 );
and ( n36950 , n36736 , n36949 );
or ( n36951 , n36735 , n36950 );
and ( n36952 , n36732 , n36951 );
or ( n36953 , n36731 , n36952 );
and ( n36954 , n36728 , n36953 );
or ( n36955 , n36727 , n36954 );
and ( n36956 , n36724 , n36955 );
or ( n36957 , n36723 , n36956 );
and ( n36958 , n36720 , n36957 );
or ( n36959 , n36719 , n36958 );
and ( n36960 , n36716 , n36959 );
or ( n36961 , n36715 , n36960 );
and ( n36962 , n36712 , n36961 );
or ( n36963 , n36711 , n36962 );
and ( n36964 , n36708 , n36963 );
or ( n36965 , n36707 , n36964 );
and ( n36966 , n36704 , n36965 );
or ( n36967 , n36703 , n36966 );
and ( n36968 , n36700 , n36967 );
or ( n36969 , n36699 , n36968 );
and ( n36970 , n36696 , n36969 );
or ( n36971 , n36695 , n36970 );
and ( n36972 , n36692 , n36971 );
or ( n36973 , n36691 , n36972 );
and ( n36974 , n36688 , n36973 );
or ( n36975 , n36687 , n36974 );
and ( n36976 , n36684 , n36975 );
or ( n36977 , n36683 , n36976 );
and ( n36978 , n36680 , n36977 );
or ( n36979 , n36679 , n36978 );
and ( n36980 , n36676 , n36979 );
or ( n36981 , n36675 , n36980 );
and ( n36982 , n36672 , n36981 );
or ( n36983 , n36671 , n36982 );
and ( n36984 , n36668 , n36983 );
or ( n36985 , n36667 , n36984 );
and ( n36986 , n36664 , n36985 );
or ( n36987 , n36663 , n36986 );
and ( n36988 , n36660 , n36987 );
or ( n36989 , n36659 , n36988 );
and ( n36990 , n36656 , n36989 );
or ( n36991 , n36655 , n36990 );
and ( n36992 , n36652 , n36991 );
or ( n36993 , n36651 , n36992 );
and ( n36994 , n36648 , n36993 );
or ( n36995 , n36647 , n36994 );
and ( n36996 , n36644 , n36995 );
or ( n36997 , n36643 , n36996 );
and ( n36998 , n36640 , n36997 );
or ( n36999 , n36639 , n36998 );
and ( n37000 , n36636 , n36999 );
or ( n37001 , n36635 , n37000 );
and ( n37002 , n36632 , n37001 );
or ( n37003 , n36631 , n37002 );
and ( n37004 , n36628 , n37003 );
or ( n37005 , n36627 , n37004 );
xor ( n37006 , n36624 , n37005 );
and ( n37007 , n33403 , n645 );
nor ( n37008 , n646 , n37007 );
nor ( n37009 , n684 , n32231 );
xor ( n37010 , n37008 , n37009 );
and ( n37011 , n35801 , n35802 );
buf ( n37012 , n37011 );
xor ( n37013 , n37010 , n37012 );
nor ( n37014 , n733 , n31083 );
xor ( n37015 , n37013 , n37014 );
and ( n37016 , n35804 , n35805 );
and ( n37017 , n35806 , n35809 );
or ( n37018 , n37016 , n37017 );
xor ( n37019 , n37015 , n37018 );
nor ( n37020 , n796 , n29948 );
xor ( n37021 , n37019 , n37020 );
and ( n37022 , n35810 , n35811 );
and ( n37023 , n35812 , n35815 );
or ( n37024 , n37022 , n37023 );
xor ( n37025 , n37021 , n37024 );
nor ( n37026 , n868 , n28833 );
xor ( n37027 , n37025 , n37026 );
and ( n37028 , n35816 , n35817 );
and ( n37029 , n35818 , n35821 );
or ( n37030 , n37028 , n37029 );
xor ( n37031 , n37027 , n37030 );
nor ( n37032 , n958 , n27737 );
xor ( n37033 , n37031 , n37032 );
and ( n37034 , n35822 , n35823 );
and ( n37035 , n35824 , n35827 );
or ( n37036 , n37034 , n37035 );
xor ( n37037 , n37033 , n37036 );
nor ( n37038 , n1062 , n26660 );
xor ( n37039 , n37037 , n37038 );
and ( n37040 , n35828 , n35829 );
and ( n37041 , n35830 , n35833 );
or ( n37042 , n37040 , n37041 );
xor ( n37043 , n37039 , n37042 );
nor ( n37044 , n1176 , n25600 );
xor ( n37045 , n37043 , n37044 );
and ( n37046 , n35834 , n35835 );
and ( n37047 , n35836 , n35839 );
or ( n37048 , n37046 , n37047 );
xor ( n37049 , n37045 , n37048 );
nor ( n37050 , n1303 , n24564 );
xor ( n37051 , n37049 , n37050 );
and ( n37052 , n35840 , n35841 );
and ( n37053 , n35842 , n35845 );
or ( n37054 , n37052 , n37053 );
xor ( n37055 , n37051 , n37054 );
nor ( n37056 , n1445 , n23541 );
xor ( n37057 , n37055 , n37056 );
and ( n37058 , n35846 , n35847 );
and ( n37059 , n35848 , n35851 );
or ( n37060 , n37058 , n37059 );
xor ( n37061 , n37057 , n37060 );
nor ( n37062 , n1598 , n22541 );
xor ( n37063 , n37061 , n37062 );
and ( n37064 , n35852 , n35853 );
and ( n37065 , n35854 , n35857 );
or ( n37066 , n37064 , n37065 );
xor ( n37067 , n37063 , n37066 );
nor ( n37068 , n1766 , n21562 );
xor ( n37069 , n37067 , n37068 );
and ( n37070 , n35858 , n35859 );
and ( n37071 , n35860 , n35863 );
or ( n37072 , n37070 , n37071 );
xor ( n37073 , n37069 , n37072 );
nor ( n37074 , n1945 , n20601 );
xor ( n37075 , n37073 , n37074 );
and ( n37076 , n35864 , n35865 );
and ( n37077 , n35866 , n35869 );
or ( n37078 , n37076 , n37077 );
xor ( n37079 , n37075 , n37078 );
nor ( n37080 , n2137 , n19657 );
xor ( n37081 , n37079 , n37080 );
and ( n37082 , n35870 , n35871 );
and ( n37083 , n35872 , n35875 );
or ( n37084 , n37082 , n37083 );
xor ( n37085 , n37081 , n37084 );
nor ( n37086 , n2343 , n18734 );
xor ( n37087 , n37085 , n37086 );
and ( n37088 , n35876 , n35877 );
and ( n37089 , n35878 , n35881 );
or ( n37090 , n37088 , n37089 );
xor ( n37091 , n37087 , n37090 );
nor ( n37092 , n2566 , n17828 );
xor ( n37093 , n37091 , n37092 );
and ( n37094 , n35882 , n35883 );
and ( n37095 , n35884 , n35887 );
or ( n37096 , n37094 , n37095 );
xor ( n37097 , n37093 , n37096 );
nor ( n37098 , n2797 , n16943 );
xor ( n37099 , n37097 , n37098 );
and ( n37100 , n35888 , n35889 );
and ( n37101 , n35890 , n35893 );
or ( n37102 , n37100 , n37101 );
xor ( n37103 , n37099 , n37102 );
nor ( n37104 , n3043 , n16077 );
xor ( n37105 , n37103 , n37104 );
and ( n37106 , n35894 , n35895 );
and ( n37107 , n35896 , n35899 );
or ( n37108 , n37106 , n37107 );
xor ( n37109 , n37105 , n37108 );
nor ( n37110 , n3300 , n15230 );
xor ( n37111 , n37109 , n37110 );
and ( n37112 , n35900 , n35901 );
and ( n37113 , n35902 , n35905 );
or ( n37114 , n37112 , n37113 );
xor ( n37115 , n37111 , n37114 );
nor ( n37116 , n3570 , n14403 );
xor ( n37117 , n37115 , n37116 );
and ( n37118 , n35906 , n35907 );
and ( n37119 , n35908 , n35911 );
or ( n37120 , n37118 , n37119 );
xor ( n37121 , n37117 , n37120 );
nor ( n37122 , n3853 , n13599 );
xor ( n37123 , n37121 , n37122 );
and ( n37124 , n35912 , n35913 );
and ( n37125 , n35914 , n35917 );
or ( n37126 , n37124 , n37125 );
xor ( n37127 , n37123 , n37126 );
nor ( n37128 , n4151 , n12808 );
xor ( n37129 , n37127 , n37128 );
and ( n37130 , n35918 , n35919 );
and ( n37131 , n35920 , n35923 );
or ( n37132 , n37130 , n37131 );
xor ( n37133 , n37129 , n37132 );
nor ( n37134 , n4458 , n12037 );
xor ( n37135 , n37133 , n37134 );
and ( n37136 , n35924 , n35925 );
and ( n37137 , n35926 , n35929 );
or ( n37138 , n37136 , n37137 );
xor ( n37139 , n37135 , n37138 );
nor ( n37140 , n4786 , n11282 );
xor ( n37141 , n37139 , n37140 );
and ( n37142 , n35930 , n35931 );
and ( n37143 , n35932 , n35935 );
or ( n37144 , n37142 , n37143 );
xor ( n37145 , n37141 , n37144 );
nor ( n37146 , n5126 , n10547 );
xor ( n37147 , n37145 , n37146 );
and ( n37148 , n35936 , n35937 );
and ( n37149 , n35938 , n35941 );
or ( n37150 , n37148 , n37149 );
xor ( n37151 , n37147 , n37150 );
nor ( n37152 , n5477 , n9829 );
xor ( n37153 , n37151 , n37152 );
and ( n37154 , n35942 , n35943 );
and ( n37155 , n35944 , n35947 );
or ( n37156 , n37154 , n37155 );
xor ( n37157 , n37153 , n37156 );
nor ( n37158 , n5838 , n8955 );
xor ( n37159 , n37157 , n37158 );
and ( n37160 , n35948 , n35949 );
and ( n37161 , n35950 , n35953 );
or ( n37162 , n37160 , n37161 );
xor ( n37163 , n37159 , n37162 );
nor ( n37164 , n6212 , n603 );
xor ( n37165 , n37163 , n37164 );
and ( n37166 , n35954 , n35955 );
and ( n37167 , n35956 , n35959 );
or ( n37168 , n37166 , n37167 );
xor ( n37169 , n37165 , n37168 );
nor ( n37170 , n6596 , n652 );
xor ( n37171 , n37169 , n37170 );
and ( n37172 , n35960 , n35961 );
and ( n37173 , n35962 , n35965 );
or ( n37174 , n37172 , n37173 );
xor ( n37175 , n37171 , n37174 );
nor ( n37176 , n6997 , n624 );
xor ( n37177 , n37175 , n37176 );
and ( n37178 , n35966 , n35967 );
and ( n37179 , n35968 , n35971 );
or ( n37180 , n37178 , n37179 );
xor ( n37181 , n37177 , n37180 );
nor ( n37182 , n7413 , n648 );
xor ( n37183 , n37181 , n37182 );
and ( n37184 , n35972 , n35973 );
and ( n37185 , n35974 , n35977 );
or ( n37186 , n37184 , n37185 );
xor ( n37187 , n37183 , n37186 );
nor ( n37188 , n7841 , n686 );
xor ( n37189 , n37187 , n37188 );
and ( n37190 , n35978 , n35979 );
and ( n37191 , n35980 , n35983 );
or ( n37192 , n37190 , n37191 );
xor ( n37193 , n37189 , n37192 );
nor ( n37194 , n8281 , n735 );
xor ( n37195 , n37193 , n37194 );
and ( n37196 , n35984 , n35985 );
and ( n37197 , n35986 , n35989 );
or ( n37198 , n37196 , n37197 );
xor ( n37199 , n37195 , n37198 );
nor ( n37200 , n8737 , n798 );
xor ( n37201 , n37199 , n37200 );
and ( n37202 , n35990 , n35991 );
and ( n37203 , n35992 , n35995 );
or ( n37204 , n37202 , n37203 );
xor ( n37205 , n37201 , n37204 );
nor ( n37206 , n9420 , n870 );
xor ( n37207 , n37205 , n37206 );
and ( n37208 , n35996 , n35997 );
and ( n37209 , n35998 , n36001 );
or ( n37210 , n37208 , n37209 );
xor ( n37211 , n37207 , n37210 );
nor ( n37212 , n10312 , n960 );
xor ( n37213 , n37211 , n37212 );
and ( n37214 , n36002 , n36003 );
and ( n37215 , n36004 , n36007 );
or ( n37216 , n37214 , n37215 );
xor ( n37217 , n37213 , n37216 );
nor ( n37218 , n11041 , n1064 );
xor ( n37219 , n37217 , n37218 );
and ( n37220 , n36008 , n36009 );
and ( n37221 , n36010 , n36013 );
or ( n37222 , n37220 , n37221 );
xor ( n37223 , n37219 , n37222 );
nor ( n37224 , n11790 , n1178 );
xor ( n37225 , n37223 , n37224 );
and ( n37226 , n36014 , n36015 );
and ( n37227 , n36016 , n36019 );
or ( n37228 , n37226 , n37227 );
xor ( n37229 , n37225 , n37228 );
nor ( n37230 , n12555 , n1305 );
xor ( n37231 , n37229 , n37230 );
and ( n37232 , n36020 , n36021 );
and ( n37233 , n36022 , n36025 );
or ( n37234 , n37232 , n37233 );
xor ( n37235 , n37231 , n37234 );
nor ( n37236 , n13340 , n1447 );
xor ( n37237 , n37235 , n37236 );
and ( n37238 , n36026 , n36027 );
and ( n37239 , n36028 , n36031 );
or ( n37240 , n37238 , n37239 );
xor ( n37241 , n37237 , n37240 );
nor ( n37242 , n14138 , n1600 );
xor ( n37243 , n37241 , n37242 );
and ( n37244 , n36032 , n36033 );
and ( n37245 , n36034 , n36037 );
or ( n37246 , n37244 , n37245 );
xor ( n37247 , n37243 , n37246 );
nor ( n37248 , n14959 , n1768 );
xor ( n37249 , n37247 , n37248 );
and ( n37250 , n36038 , n36039 );
and ( n37251 , n36040 , n36043 );
or ( n37252 , n37250 , n37251 );
xor ( n37253 , n37249 , n37252 );
nor ( n37254 , n15800 , n1947 );
xor ( n37255 , n37253 , n37254 );
and ( n37256 , n36044 , n36045 );
and ( n37257 , n36046 , n36049 );
or ( n37258 , n37256 , n37257 );
xor ( n37259 , n37255 , n37258 );
nor ( n37260 , n16660 , n2139 );
xor ( n37261 , n37259 , n37260 );
and ( n37262 , n36050 , n36051 );
and ( n37263 , n36052 , n36055 );
or ( n37264 , n37262 , n37263 );
xor ( n37265 , n37261 , n37264 );
nor ( n37266 , n17539 , n2345 );
xor ( n37267 , n37265 , n37266 );
and ( n37268 , n36056 , n36057 );
and ( n37269 , n36058 , n36061 );
or ( n37270 , n37268 , n37269 );
xor ( n37271 , n37267 , n37270 );
nor ( n37272 , n18439 , n2568 );
xor ( n37273 , n37271 , n37272 );
and ( n37274 , n36062 , n36063 );
and ( n37275 , n36064 , n36067 );
or ( n37276 , n37274 , n37275 );
xor ( n37277 , n37273 , n37276 );
nor ( n37278 , n19356 , n2799 );
xor ( n37279 , n37277 , n37278 );
and ( n37280 , n36068 , n36069 );
and ( n37281 , n36070 , n36073 );
or ( n37282 , n37280 , n37281 );
xor ( n37283 , n37279 , n37282 );
nor ( n37284 , n20294 , n3045 );
xor ( n37285 , n37283 , n37284 );
and ( n37286 , n36074 , n36075 );
and ( n37287 , n36076 , n36079 );
or ( n37288 , n37286 , n37287 );
xor ( n37289 , n37285 , n37288 );
nor ( n37290 , n21249 , n3302 );
xor ( n37291 , n37289 , n37290 );
and ( n37292 , n36080 , n36081 );
and ( n37293 , n36082 , n36085 );
or ( n37294 , n37292 , n37293 );
xor ( n37295 , n37291 , n37294 );
nor ( n37296 , n22222 , n3572 );
xor ( n37297 , n37295 , n37296 );
and ( n37298 , n36086 , n36087 );
and ( n37299 , n36088 , n36091 );
or ( n37300 , n37298 , n37299 );
xor ( n37301 , n37297 , n37300 );
nor ( n37302 , n23216 , n3855 );
xor ( n37303 , n37301 , n37302 );
and ( n37304 , n36092 , n36093 );
and ( n37305 , n36094 , n36097 );
or ( n37306 , n37304 , n37305 );
xor ( n37307 , n37303 , n37306 );
nor ( n37308 , n24233 , n4153 );
xor ( n37309 , n37307 , n37308 );
and ( n37310 , n36098 , n36099 );
and ( n37311 , n36100 , n36103 );
or ( n37312 , n37310 , n37311 );
xor ( n37313 , n37309 , n37312 );
nor ( n37314 , n25263 , n4460 );
xor ( n37315 , n37313 , n37314 );
and ( n37316 , n36104 , n36105 );
and ( n37317 , n36106 , n36109 );
or ( n37318 , n37316 , n37317 );
xor ( n37319 , n37315 , n37318 );
nor ( n37320 , n26317 , n4788 );
xor ( n37321 , n37319 , n37320 );
and ( n37322 , n36110 , n36111 );
and ( n37323 , n36112 , n36115 );
or ( n37324 , n37322 , n37323 );
xor ( n37325 , n37321 , n37324 );
nor ( n37326 , n27388 , n5128 );
xor ( n37327 , n37325 , n37326 );
and ( n37328 , n36116 , n36117 );
and ( n37329 , n36118 , n36121 );
or ( n37330 , n37328 , n37329 );
xor ( n37331 , n37327 , n37330 );
nor ( n37332 , n28478 , n5479 );
xor ( n37333 , n37331 , n37332 );
and ( n37334 , n36122 , n36123 );
and ( n37335 , n36124 , n36127 );
or ( n37336 , n37334 , n37335 );
xor ( n37337 , n37333 , n37336 );
nor ( n37338 , n29587 , n5840 );
xor ( n37339 , n37337 , n37338 );
and ( n37340 , n36128 , n36129 );
and ( n37341 , n36130 , n36133 );
or ( n37342 , n37340 , n37341 );
xor ( n37343 , n37339 , n37342 );
nor ( n37344 , n30716 , n6214 );
xor ( n37345 , n37343 , n37344 );
and ( n37346 , n36134 , n36135 );
and ( n37347 , n36136 , n36139 );
or ( n37348 , n37346 , n37347 );
xor ( n37349 , n37345 , n37348 );
nor ( n37350 , n31858 , n6598 );
xor ( n37351 , n37349 , n37350 );
and ( n37352 , n36140 , n36141 );
and ( n37353 , n36142 , n36145 );
or ( n37354 , n37352 , n37353 );
xor ( n37355 , n37351 , n37354 );
nor ( n37356 , n33024 , n6999 );
xor ( n37357 , n37355 , n37356 );
and ( n37358 , n36146 , n36147 );
and ( n37359 , n36148 , n36151 );
or ( n37360 , n37358 , n37359 );
xor ( n37361 , n37357 , n37360 );
nor ( n37362 , n34215 , n7415 );
xor ( n37363 , n37361 , n37362 );
and ( n37364 , n36152 , n36153 );
and ( n37365 , n36154 , n36157 );
or ( n37366 , n37364 , n37365 );
xor ( n37367 , n37363 , n37366 );
nor ( n37368 , n35410 , n7843 );
xor ( n37369 , n37367 , n37368 );
and ( n37370 , n36158 , n36159 );
and ( n37371 , n36160 , n36163 );
or ( n37372 , n37370 , n37371 );
xor ( n37373 , n37369 , n37372 );
nor ( n37374 , n36611 , n8283 );
xor ( n37375 , n37373 , n37374 );
and ( n37376 , n36164 , n36165 );
and ( n37377 , n36166 , n36169 );
or ( n37378 , n37376 , n37377 );
xor ( n37379 , n37375 , n37378 );
and ( n37380 , n36182 , n36186 );
and ( n37381 , n36186 , n36597 );
and ( n37382 , n36182 , n36597 );
or ( n37383 , n37380 , n37381 , n37382 );
and ( n37384 , n33774 , n635 );
not ( n37385 , n635 );
nor ( n37386 , n37384 , n37385 );
xor ( n37387 , n37383 , n37386 );
and ( n37388 , n36195 , n36199 );
and ( n37389 , n36199 , n36267 );
and ( n37390 , n36195 , n36267 );
or ( n37391 , n37388 , n37389 , n37390 );
and ( n37392 , n36191 , n36268 );
and ( n37393 , n36268 , n36596 );
and ( n37394 , n36191 , n36596 );
or ( n37395 , n37392 , n37393 , n37394 );
xor ( n37396 , n37391 , n37395 );
and ( n37397 , n36273 , n36393 );
and ( n37398 , n36393 , n36595 );
and ( n37399 , n36273 , n36595 );
or ( n37400 , n37397 , n37398 , n37399 );
and ( n37401 , n36204 , n36208 );
and ( n37402 , n36208 , n36266 );
and ( n37403 , n36204 , n36266 );
or ( n37404 , n37401 , n37402 , n37403 );
and ( n37405 , n36277 , n36281 );
and ( n37406 , n36281 , n36392 );
and ( n37407 , n36277 , n36392 );
or ( n37408 , n37405 , n37406 , n37407 );
xor ( n37409 , n37404 , n37408 );
and ( n37410 , n36235 , n36239 );
and ( n37411 , n36239 , n36245 );
and ( n37412 , n36235 , n36245 );
or ( n37413 , n37410 , n37411 , n37412 );
and ( n37414 , n36213 , n36217 );
and ( n37415 , n36217 , n36265 );
and ( n37416 , n36213 , n36265 );
or ( n37417 , n37414 , n37415 , n37416 );
xor ( n37418 , n37413 , n37417 );
and ( n37419 , n36222 , n36226 );
and ( n37420 , n36226 , n36264 );
and ( n37421 , n36222 , n36264 );
or ( n37422 , n37419 , n37420 , n37421 );
and ( n37423 , n36290 , n36315 );
and ( n37424 , n36315 , n36353 );
and ( n37425 , n36290 , n36353 );
or ( n37426 , n37423 , n37424 , n37425 );
xor ( n37427 , n37422 , n37426 );
and ( n37428 , n36231 , n36246 );
and ( n37429 , n36246 , n36263 );
and ( n37430 , n36231 , n36263 );
or ( n37431 , n37428 , n37429 , n37430 );
and ( n37432 , n36294 , n36298 );
and ( n37433 , n36298 , n36314 );
and ( n37434 , n36294 , n36314 );
or ( n37435 , n37432 , n37433 , n37434 );
xor ( n37436 , n37431 , n37435 );
and ( n37437 , n36251 , n36256 );
and ( n37438 , n36256 , n36262 );
and ( n37439 , n36251 , n36262 );
or ( n37440 , n37437 , n37438 , n37439 );
and ( n37441 , n36241 , n36242 );
and ( n37442 , n36242 , n36244 );
and ( n37443 , n36241 , n36244 );
or ( n37444 , n37441 , n37442 , n37443 );
and ( n37445 , n36252 , n36253 );
and ( n37446 , n36253 , n36255 );
and ( n37447 , n36252 , n36255 );
or ( n37448 , n37445 , n37446 , n37447 );
xor ( n37449 , n37444 , n37448 );
and ( n37450 , n30695 , n771 );
and ( n37451 , n31836 , n719 );
xor ( n37452 , n37450 , n37451 );
and ( n37453 , n32649 , n663 );
xor ( n37454 , n37452 , n37453 );
xor ( n37455 , n37449 , n37454 );
xor ( n37456 , n37440 , n37455 );
and ( n37457 , n36258 , n36259 );
and ( n37458 , n36259 , n36261 );
and ( n37459 , n36258 , n36261 );
or ( n37460 , n37457 , n37458 , n37459 );
and ( n37461 , n27361 , n1034 );
and ( n37462 , n28456 , n940 );
xor ( n37463 , n37461 , n37462 );
and ( n37464 , n29559 , n840 );
xor ( n37465 , n37463 , n37464 );
xor ( n37466 , n37460 , n37465 );
and ( n37467 , n24214 , n1424 );
and ( n37468 , n25243 , n1254 );
xor ( n37469 , n37467 , n37468 );
and ( n37470 , n26296 , n1134 );
xor ( n37471 , n37469 , n37470 );
xor ( n37472 , n37466 , n37471 );
xor ( n37473 , n37456 , n37472 );
xor ( n37474 , n37436 , n37473 );
xor ( n37475 , n37427 , n37474 );
xor ( n37476 , n37418 , n37475 );
xor ( n37477 , n37409 , n37476 );
xor ( n37478 , n37400 , n37477 );
and ( n37479 , n36398 , n36476 );
and ( n37480 , n36476 , n36594 );
and ( n37481 , n36398 , n36594 );
or ( n37482 , n37479 , n37480 , n37481 );
and ( n37483 , n36286 , n36354 );
and ( n37484 , n36354 , n36391 );
and ( n37485 , n36286 , n36391 );
or ( n37486 , n37483 , n37484 , n37485 );
and ( n37487 , n36402 , n36406 );
and ( n37488 , n36406 , n36475 );
and ( n37489 , n36402 , n36475 );
or ( n37490 , n37487 , n37488 , n37489 );
xor ( n37491 , n37486 , n37490 );
and ( n37492 , n36359 , n36363 );
and ( n37493 , n36363 , n36390 );
and ( n37494 , n36359 , n36390 );
or ( n37495 , n37492 , n37493 , n37494 );
and ( n37496 , n36320 , n36336 );
and ( n37497 , n36336 , n36352 );
and ( n37498 , n36320 , n36352 );
or ( n37499 , n37496 , n37497 , n37498 );
and ( n37500 , n36303 , n36307 );
and ( n37501 , n36307 , n36313 );
and ( n37502 , n36303 , n36313 );
or ( n37503 , n37500 , n37501 , n37502 );
and ( n37504 , n36324 , n36329 );
and ( n37505 , n36329 , n36335 );
and ( n37506 , n36324 , n36335 );
or ( n37507 , n37504 , n37505 , n37506 );
xor ( n37508 , n37503 , n37507 );
and ( n37509 , n36309 , n36310 );
and ( n37510 , n36310 , n36312 );
and ( n37511 , n36309 , n36312 );
or ( n37512 , n37509 , n37510 , n37511 );
and ( n37513 , n36325 , n36326 );
and ( n37514 , n36326 , n36328 );
and ( n37515 , n36325 , n36328 );
or ( n37516 , n37513 , n37514 , n37515 );
xor ( n37517 , n37512 , n37516 );
and ( n37518 , n21216 , n1882 );
and ( n37519 , n22186 , n1738 );
xor ( n37520 , n37518 , n37519 );
and ( n37521 , n22892 , n1551 );
xor ( n37522 , n37520 , n37521 );
xor ( n37523 , n37517 , n37522 );
xor ( n37524 , n37508 , n37523 );
xor ( n37525 , n37499 , n37524 );
and ( n37526 , n36341 , n36345 );
and ( n37527 , n36345 , n36351 );
and ( n37528 , n36341 , n36351 );
or ( n37529 , n37526 , n37527 , n37528 );
and ( n37530 , n36331 , n36332 );
and ( n37531 , n36332 , n36334 );
and ( n37532 , n36331 , n36334 );
or ( n37533 , n37530 , n37531 , n37532 );
and ( n37534 , n18144 , n2544 );
and ( n37535 , n19324 , n2298 );
xor ( n37536 , n37534 , n37535 );
and ( n37537 , n20233 , n2100 );
xor ( n37538 , n37536 , n37537 );
xor ( n37539 , n37533 , n37538 );
and ( n37540 , n15758 , n3271 );
and ( n37541 , n16637 , n2981 );
xor ( n37542 , n37540 , n37541 );
and ( n37543 , n17512 , n2739 );
xor ( n37544 , n37542 , n37543 );
xor ( n37545 , n37539 , n37544 );
xor ( n37546 , n37529 , n37545 );
and ( n37547 , n36347 , n36348 );
and ( n37548 , n36348 , n36350 );
and ( n37549 , n36347 , n36350 );
or ( n37550 , n37547 , n37548 , n37549 );
and ( n37551 , n36378 , n36379 );
and ( n37552 , n36379 , n36381 );
and ( n37553 , n36378 , n36381 );
or ( n37554 , n37551 , n37552 , n37553 );
xor ( n37555 , n37550 , n37554 );
and ( n37556 , n13322 , n4102 );
and ( n37557 , n14118 , n3749 );
xor ( n37558 , n37556 , n37557 );
and ( n37559 , n14938 , n3495 );
xor ( n37560 , n37558 , n37559 );
xor ( n37561 , n37555 , n37560 );
xor ( n37562 , n37546 , n37561 );
xor ( n37563 , n37525 , n37562 );
xor ( n37564 , n37495 , n37563 );
and ( n37565 , n36368 , n36372 );
and ( n37566 , n36372 , n36389 );
and ( n37567 , n36368 , n36389 );
or ( n37568 , n37565 , n37566 , n37567 );
and ( n37569 , n36415 , n36430 );
and ( n37570 , n36430 , n36447 );
and ( n37571 , n36415 , n36447 );
or ( n37572 , n37569 , n37570 , n37571 );
xor ( n37573 , n37568 , n37572 );
and ( n37574 , n36377 , n36382 );
and ( n37575 , n36382 , n36388 );
and ( n37576 , n36377 , n36388 );
or ( n37577 , n37574 , n37575 , n37576 );
and ( n37578 , n36419 , n36423 );
and ( n37579 , n36423 , n36429 );
and ( n37580 , n36419 , n36429 );
or ( n37581 , n37578 , n37579 , n37580 );
xor ( n37582 , n37577 , n37581 );
and ( n37583 , n36384 , n36385 );
and ( n37584 , n36385 , n36387 );
and ( n37585 , n36384 , n36387 );
or ( n37586 , n37583 , n37584 , n37585 );
and ( n37587 , n11015 , n5103 );
and ( n37588 , n11769 , n4730 );
xor ( n37589 , n37587 , n37588 );
and ( n37590 , n12320 , n4403 );
xor ( n37591 , n37589 , n37590 );
xor ( n37592 , n37586 , n37591 );
and ( n37593 , n8718 , n6132 );
and ( n37594 , n9400 , n5765 );
xor ( n37595 , n37593 , n37594 );
and ( n37596 , n10291 , n5408 );
xor ( n37597 , n37595 , n37596 );
xor ( n37598 , n37592 , n37597 );
xor ( n37599 , n37582 , n37598 );
xor ( n37600 , n37573 , n37599 );
xor ( n37601 , n37564 , n37600 );
xor ( n37602 , n37491 , n37601 );
xor ( n37603 , n37482 , n37602 );
and ( n37604 , n36481 , n36528 );
and ( n37605 , n36528 , n36593 );
and ( n37606 , n36481 , n36593 );
or ( n37607 , n37604 , n37605 , n37606 );
and ( n37608 , n36411 , n36448 );
and ( n37609 , n36448 , n36474 );
and ( n37610 , n36411 , n36474 );
or ( n37611 , n37608 , n37609 , n37610 );
and ( n37612 , n36485 , n36489 );
and ( n37613 , n36489 , n36527 );
and ( n37614 , n36485 , n36527 );
or ( n37615 , n37612 , n37613 , n37614 );
xor ( n37616 , n37611 , n37615 );
and ( n37617 , n36453 , n36457 );
and ( n37618 , n36457 , n36473 );
and ( n37619 , n36453 , n36473 );
or ( n37620 , n37617 , n37618 , n37619 );
and ( n37621 , n36435 , n36440 );
and ( n37622 , n36440 , n36446 );
and ( n37623 , n36435 , n36446 );
or ( n37624 , n37621 , n37622 , n37623 );
and ( n37625 , n36425 , n36426 );
and ( n37626 , n36426 , n36428 );
and ( n37627 , n36425 , n36428 );
or ( n37628 , n37625 , n37626 , n37627 );
and ( n37629 , n36436 , n36437 );
and ( n37630 , n36437 , n36439 );
and ( n37631 , n36436 , n36439 );
or ( n37632 , n37629 , n37630 , n37631 );
xor ( n37633 , n37628 , n37632 );
buf ( n37634 , n7385 );
and ( n37635 , n7808 , n6971 );
xor ( n37636 , n37634 , n37635 );
and ( n37637 , n8079 , n6504 );
xor ( n37638 , n37636 , n37637 );
xor ( n37639 , n37633 , n37638 );
xor ( n37640 , n37624 , n37639 );
and ( n37641 , n36442 , n36443 );
and ( n37642 , n36443 , n36445 );
and ( n37643 , n36442 , n36445 );
or ( n37644 , n37641 , n37642 , n37643 );
and ( n37645 , n6187 , n8669 );
and ( n37646 , n6569 , n8243 );
xor ( n37647 , n37645 , n37646 );
and ( n37648 , n6816 , n7662 );
xor ( n37649 , n37647 , n37648 );
xor ( n37650 , n37644 , n37649 );
and ( n37651 , n4959 , n10977 );
and ( n37652 , n5459 , n10239 );
xor ( n37653 , n37651 , n37652 );
and ( n37654 , n5819 , n9348 );
xor ( n37655 , n37653 , n37654 );
xor ( n37656 , n37650 , n37655 );
xor ( n37657 , n37640 , n37656 );
xor ( n37658 , n37620 , n37657 );
and ( n37659 , n36462 , n36466 );
and ( n37660 , n36466 , n36472 );
and ( n37661 , n36462 , n36472 );
or ( n37662 , n37659 , n37660 , n37661 );
and ( n37663 , n36498 , n36503 );
and ( n37664 , n36503 , n36509 );
and ( n37665 , n36498 , n36509 );
or ( n37666 , n37663 , n37664 , n37665 );
xor ( n37667 , n37662 , n37666 );
and ( n37668 , n36468 , n36469 );
and ( n37669 , n36469 , n36471 );
and ( n37670 , n36468 , n36471 );
or ( n37671 , n37668 , n37669 , n37670 );
and ( n37672 , n36499 , n36500 );
and ( n37673 , n36500 , n36502 );
and ( n37674 , n36499 , n36502 );
or ( n37675 , n37672 , n37673 , n37674 );
xor ( n37676 , n37671 , n37675 );
and ( n37677 , n4132 , n13256 );
and ( n37678 , n4438 , n12531 );
xor ( n37679 , n37677 , n37678 );
and ( n37680 , n4766 , n11718 );
xor ( n37681 , n37679 , n37680 );
xor ( n37682 , n37676 , n37681 );
xor ( n37683 , n37667 , n37682 );
xor ( n37684 , n37658 , n37683 );
xor ( n37685 , n37616 , n37684 );
xor ( n37686 , n37607 , n37685 );
and ( n37687 , n36533 , n36559 );
and ( n37688 , n36559 , n36592 );
and ( n37689 , n36533 , n36592 );
or ( n37690 , n37687 , n37688 , n37689 );
and ( n37691 , n36494 , n36510 );
and ( n37692 , n36510 , n36526 );
and ( n37693 , n36494 , n36526 );
or ( n37694 , n37691 , n37692 , n37693 );
and ( n37695 , n36537 , n36541 );
and ( n37696 , n36541 , n36558 );
and ( n37697 , n36537 , n36558 );
or ( n37698 , n37695 , n37696 , n37697 );
xor ( n37699 , n37694 , n37698 );
and ( n37700 , n36515 , n36519 );
and ( n37701 , n36519 , n36525 );
and ( n37702 , n36515 , n36525 );
or ( n37703 , n37700 , n37701 , n37702 );
and ( n37704 , n36505 , n36506 );
and ( n37705 , n36506 , n36508 );
and ( n37706 , n36505 , n36508 );
or ( n37707 , n37704 , n37705 , n37706 );
and ( n37708 , n3182 , n15691 );
and ( n37709 , n3545 , n14838 );
xor ( n37710 , n37708 , n37709 );
and ( n37711 , n3801 , n14044 );
xor ( n37712 , n37710 , n37711 );
xor ( n37713 , n37707 , n37712 );
and ( n37714 , n2462 , n18407 );
and ( n37715 , n2779 , n17422 );
xor ( n37716 , n37714 , n37715 );
and ( n37717 , n3024 , n16550 );
xor ( n37718 , n37716 , n37717 );
xor ( n37719 , n37713 , n37718 );
xor ( n37720 , n37703 , n37719 );
and ( n37721 , n36521 , n36522 );
and ( n37722 , n36522 , n36524 );
and ( n37723 , n36521 , n36524 );
or ( n37724 , n37721 , n37722 , n37723 );
and ( n37725 , n36547 , n36548 );
and ( n37726 , n36548 , n36550 );
and ( n37727 , n36547 , n36550 );
or ( n37728 , n37725 , n37726 , n37727 );
xor ( n37729 , n37724 , n37728 );
and ( n37730 , n1933 , n20976 );
and ( n37731 , n2120 , n20156 );
xor ( n37732 , n37730 , n37731 );
and ( n37733 , n2324 , n19222 );
xor ( n37734 , n37732 , n37733 );
xor ( n37735 , n37729 , n37734 );
xor ( n37736 , n37720 , n37735 );
xor ( n37737 , n37699 , n37736 );
xor ( n37738 , n37690 , n37737 );
and ( n37739 , n36564 , n36579 );
and ( n37740 , n36579 , n36591 );
and ( n37741 , n36564 , n36591 );
or ( n37742 , n37739 , n37740 , n37741 );
and ( n37743 , n36546 , n36551 );
and ( n37744 , n36551 , n36557 );
and ( n37745 , n36546 , n36557 );
or ( n37746 , n37743 , n37744 , n37745 );
and ( n37747 , n36568 , n36572 );
and ( n37748 , n36572 , n36578 );
and ( n37749 , n36568 , n36578 );
or ( n37750 , n37747 , n37748 , n37749 );
xor ( n37751 , n37746 , n37750 );
and ( n37752 , n36553 , n36554 );
and ( n37753 , n36554 , n36556 );
and ( n37754 , n36553 , n36556 );
or ( n37755 , n37752 , n37753 , n37754 );
and ( n37756 , n1383 , n24137 );
and ( n37757 , n1580 , n23075 );
xor ( n37758 , n37756 , n37757 );
and ( n37759 , n1694 , n22065 );
xor ( n37760 , n37758 , n37759 );
xor ( n37761 , n37755 , n37760 );
and ( n37762 , n1047 , n27296 );
and ( n37763 , n1164 , n26216 );
xor ( n37764 , n37762 , n37763 );
and ( n37765 , n1287 , n25163 );
xor ( n37766 , n37764 , n37765 );
xor ( n37767 , n37761 , n37766 );
xor ( n37768 , n37751 , n37767 );
xor ( n37769 , n37742 , n37768 );
and ( n37770 , n36581 , n36584 );
and ( n37771 , n36584 , n36590 );
and ( n37772 , n36581 , n36590 );
or ( n37773 , n37770 , n37771 , n37772 );
not ( n37774 , n632 );
and ( n37775 , n34193 , n632 );
nor ( n37776 , n37774 , n37775 );
and ( n37777 , n671 , n32999 );
xor ( n37778 , n37776 , n37777 );
and ( n37779 , n715 , n31761 );
xor ( n37780 , n37778 , n37779 );
xor ( n37781 , n37773 , n37780 );
and ( n37782 , n36574 , n36575 );
and ( n37783 , n36575 , n36577 );
and ( n37784 , n36574 , n36577 );
or ( n37785 , n37782 , n37783 , n37784 );
and ( n37786 , n36586 , n36587 );
and ( n37787 , n36587 , n36589 );
and ( n37788 , n36586 , n36589 );
or ( n37789 , n37786 , n37787 , n37788 );
xor ( n37790 , n37785 , n37789 );
and ( n37791 , n783 , n30629 );
and ( n37792 , n856 , n29508 );
xor ( n37793 , n37791 , n37792 );
and ( n37794 , n925 , n28406 );
xor ( n37795 , n37793 , n37794 );
xor ( n37796 , n37790 , n37795 );
xor ( n37797 , n37781 , n37796 );
xor ( n37798 , n37769 , n37797 );
xor ( n37799 , n37738 , n37798 );
xor ( n37800 , n37686 , n37799 );
xor ( n37801 , n37603 , n37800 );
xor ( n37802 , n37478 , n37801 );
xor ( n37803 , n37396 , n37802 );
xor ( n37804 , n37387 , n37803 );
and ( n37805 , n36174 , n36177 );
and ( n37806 , n36177 , n36598 );
and ( n37807 , n36174 , n36598 );
or ( n37808 , n37805 , n37806 , n37807 );
xor ( n37809 , n37804 , n37808 );
and ( n37810 , n36599 , n36603 );
and ( n37811 , n36604 , n36607 );
or ( n37812 , n37810 , n37811 );
xor ( n37813 , n37809 , n37812 );
buf ( n37814 , n37813 );
buf ( n37815 , n37814 );
not ( n37816 , n37815 );
nor ( n37817 , n37816 , n8739 );
xor ( n37818 , n37379 , n37817 );
and ( n37819 , n36170 , n36612 );
and ( n37820 , n36613 , n36616 );
or ( n37821 , n37819 , n37820 );
xor ( n37822 , n37818 , n37821 );
buf ( n37823 , n37822 );
buf ( n37824 , n37823 );
not ( n37825 , n37824 );
buf ( n37826 , n565 );
not ( n37827 , n37826 );
nor ( n37828 , n37825 , n37827 );
xor ( n37829 , n37006 , n37828 );
xor ( n37830 , n36628 , n37003 );
nor ( n37831 , n36620 , n37827 );
and ( n37832 , n37830 , n37831 );
xor ( n37833 , n37830 , n37831 );
xor ( n37834 , n36632 , n37001 );
nor ( n37835 , n35419 , n37827 );
and ( n37836 , n37834 , n37835 );
xor ( n37837 , n37834 , n37835 );
xor ( n37838 , n36636 , n36999 );
nor ( n37839 , n34224 , n37827 );
and ( n37840 , n37838 , n37839 );
xor ( n37841 , n37838 , n37839 );
xor ( n37842 , n36640 , n36997 );
nor ( n37843 , n33033 , n37827 );
and ( n37844 , n37842 , n37843 );
xor ( n37845 , n37842 , n37843 );
xor ( n37846 , n36644 , n36995 );
nor ( n37847 , n31867 , n37827 );
and ( n37848 , n37846 , n37847 );
xor ( n37849 , n37846 , n37847 );
xor ( n37850 , n36648 , n36993 );
nor ( n37851 , n30725 , n37827 );
and ( n37852 , n37850 , n37851 );
xor ( n37853 , n37850 , n37851 );
xor ( n37854 , n36652 , n36991 );
nor ( n37855 , n29596 , n37827 );
and ( n37856 , n37854 , n37855 );
xor ( n37857 , n37854 , n37855 );
xor ( n37858 , n36656 , n36989 );
nor ( n37859 , n28487 , n37827 );
and ( n37860 , n37858 , n37859 );
xor ( n37861 , n37858 , n37859 );
xor ( n37862 , n36660 , n36987 );
nor ( n37863 , n27397 , n37827 );
and ( n37864 , n37862 , n37863 );
xor ( n37865 , n37862 , n37863 );
xor ( n37866 , n36664 , n36985 );
nor ( n37867 , n26326 , n37827 );
and ( n37868 , n37866 , n37867 );
xor ( n37869 , n37866 , n37867 );
xor ( n37870 , n36668 , n36983 );
nor ( n37871 , n25272 , n37827 );
and ( n37872 , n37870 , n37871 );
xor ( n37873 , n37870 , n37871 );
xor ( n37874 , n36672 , n36981 );
nor ( n37875 , n24242 , n37827 );
and ( n37876 , n37874 , n37875 );
xor ( n37877 , n37874 , n37875 );
xor ( n37878 , n36676 , n36979 );
nor ( n37879 , n23225 , n37827 );
and ( n37880 , n37878 , n37879 );
xor ( n37881 , n37878 , n37879 );
xor ( n37882 , n36680 , n36977 );
nor ( n37883 , n22231 , n37827 );
and ( n37884 , n37882 , n37883 );
xor ( n37885 , n37882 , n37883 );
xor ( n37886 , n36684 , n36975 );
nor ( n37887 , n21258 , n37827 );
and ( n37888 , n37886 , n37887 );
xor ( n37889 , n37886 , n37887 );
xor ( n37890 , n36688 , n36973 );
nor ( n37891 , n20303 , n37827 );
and ( n37892 , n37890 , n37891 );
xor ( n37893 , n37890 , n37891 );
xor ( n37894 , n36692 , n36971 );
nor ( n37895 , n19365 , n37827 );
and ( n37896 , n37894 , n37895 );
xor ( n37897 , n37894 , n37895 );
xor ( n37898 , n36696 , n36969 );
nor ( n37899 , n18448 , n37827 );
and ( n37900 , n37898 , n37899 );
xor ( n37901 , n37898 , n37899 );
xor ( n37902 , n36700 , n36967 );
nor ( n37903 , n17548 , n37827 );
and ( n37904 , n37902 , n37903 );
xor ( n37905 , n37902 , n37903 );
xor ( n37906 , n36704 , n36965 );
nor ( n37907 , n16669 , n37827 );
and ( n37908 , n37906 , n37907 );
xor ( n37909 , n37906 , n37907 );
xor ( n37910 , n36708 , n36963 );
nor ( n37911 , n15809 , n37827 );
and ( n37912 , n37910 , n37911 );
xor ( n37913 , n37910 , n37911 );
xor ( n37914 , n36712 , n36961 );
nor ( n37915 , n14968 , n37827 );
and ( n37916 , n37914 , n37915 );
xor ( n37917 , n37914 , n37915 );
xor ( n37918 , n36716 , n36959 );
nor ( n37919 , n14147 , n37827 );
and ( n37920 , n37918 , n37919 );
xor ( n37921 , n37918 , n37919 );
xor ( n37922 , n36720 , n36957 );
nor ( n37923 , n13349 , n37827 );
and ( n37924 , n37922 , n37923 );
xor ( n37925 , n37922 , n37923 );
xor ( n37926 , n36724 , n36955 );
nor ( n37927 , n12564 , n37827 );
and ( n37928 , n37926 , n37927 );
xor ( n37929 , n37926 , n37927 );
xor ( n37930 , n36728 , n36953 );
nor ( n37931 , n11799 , n37827 );
and ( n37932 , n37930 , n37931 );
xor ( n37933 , n37930 , n37931 );
xor ( n37934 , n36732 , n36951 );
nor ( n37935 , n11050 , n37827 );
and ( n37936 , n37934 , n37935 );
xor ( n37937 , n37934 , n37935 );
xor ( n37938 , n36736 , n36949 );
nor ( n37939 , n10321 , n37827 );
and ( n37940 , n37938 , n37939 );
xor ( n37941 , n37938 , n37939 );
xor ( n37942 , n36740 , n36947 );
nor ( n37943 , n9429 , n37827 );
and ( n37944 , n37942 , n37943 );
xor ( n37945 , n37942 , n37943 );
xor ( n37946 , n36744 , n36945 );
nor ( n37947 , n8949 , n37827 );
and ( n37948 , n37946 , n37947 );
xor ( n37949 , n37946 , n37947 );
xor ( n37950 , n36748 , n36943 );
nor ( n37951 , n9437 , n37827 );
and ( n37952 , n37950 , n37951 );
xor ( n37953 , n37950 , n37951 );
xor ( n37954 , n36752 , n36941 );
nor ( n37955 , n9446 , n37827 );
and ( n37956 , n37954 , n37955 );
xor ( n37957 , n37954 , n37955 );
xor ( n37958 , n36756 , n36939 );
nor ( n37959 , n9455 , n37827 );
and ( n37960 , n37958 , n37959 );
xor ( n37961 , n37958 , n37959 );
xor ( n37962 , n36760 , n36937 );
nor ( n37963 , n9464 , n37827 );
and ( n37964 , n37962 , n37963 );
xor ( n37965 , n37962 , n37963 );
xor ( n37966 , n36764 , n36935 );
nor ( n37967 , n9473 , n37827 );
and ( n37968 , n37966 , n37967 );
xor ( n37969 , n37966 , n37967 );
xor ( n37970 , n36768 , n36933 );
nor ( n37971 , n9482 , n37827 );
and ( n37972 , n37970 , n37971 );
xor ( n37973 , n37970 , n37971 );
xor ( n37974 , n36772 , n36931 );
nor ( n37975 , n9491 , n37827 );
and ( n37976 , n37974 , n37975 );
xor ( n37977 , n37974 , n37975 );
xor ( n37978 , n36776 , n36929 );
nor ( n37979 , n9500 , n37827 );
and ( n37980 , n37978 , n37979 );
xor ( n37981 , n37978 , n37979 );
xor ( n37982 , n36780 , n36927 );
nor ( n37983 , n9509 , n37827 );
and ( n37984 , n37982 , n37983 );
xor ( n37985 , n37982 , n37983 );
xor ( n37986 , n36784 , n36925 );
nor ( n37987 , n9518 , n37827 );
and ( n37988 , n37986 , n37987 );
xor ( n37989 , n37986 , n37987 );
xor ( n37990 , n36788 , n36923 );
nor ( n37991 , n9527 , n37827 );
and ( n37992 , n37990 , n37991 );
xor ( n37993 , n37990 , n37991 );
xor ( n37994 , n36792 , n36921 );
nor ( n37995 , n9536 , n37827 );
and ( n37996 , n37994 , n37995 );
xor ( n37997 , n37994 , n37995 );
xor ( n37998 , n36796 , n36919 );
nor ( n37999 , n9545 , n37827 );
and ( n38000 , n37998 , n37999 );
xor ( n38001 , n37998 , n37999 );
xor ( n38002 , n36800 , n36917 );
nor ( n38003 , n9554 , n37827 );
and ( n38004 , n38002 , n38003 );
xor ( n38005 , n38002 , n38003 );
xor ( n38006 , n36804 , n36915 );
nor ( n38007 , n9563 , n37827 );
and ( n38008 , n38006 , n38007 );
xor ( n38009 , n38006 , n38007 );
xor ( n38010 , n36808 , n36913 );
nor ( n38011 , n9572 , n37827 );
and ( n38012 , n38010 , n38011 );
xor ( n38013 , n38010 , n38011 );
xor ( n38014 , n36812 , n36911 );
nor ( n38015 , n9581 , n37827 );
and ( n38016 , n38014 , n38015 );
xor ( n38017 , n38014 , n38015 );
xor ( n38018 , n36816 , n36909 );
nor ( n38019 , n9590 , n37827 );
and ( n38020 , n38018 , n38019 );
xor ( n38021 , n38018 , n38019 );
xor ( n38022 , n36820 , n36907 );
nor ( n38023 , n9599 , n37827 );
and ( n38024 , n38022 , n38023 );
xor ( n38025 , n38022 , n38023 );
xor ( n38026 , n36824 , n36905 );
nor ( n38027 , n9608 , n37827 );
and ( n38028 , n38026 , n38027 );
xor ( n38029 , n38026 , n38027 );
xor ( n38030 , n36828 , n36903 );
nor ( n38031 , n9617 , n37827 );
and ( n38032 , n38030 , n38031 );
xor ( n38033 , n38030 , n38031 );
xor ( n38034 , n36832 , n36901 );
nor ( n38035 , n9626 , n37827 );
and ( n38036 , n38034 , n38035 );
xor ( n38037 , n38034 , n38035 );
xor ( n38038 , n36836 , n36899 );
nor ( n38039 , n9635 , n37827 );
and ( n38040 , n38038 , n38039 );
xor ( n38041 , n38038 , n38039 );
xor ( n38042 , n36840 , n36897 );
nor ( n38043 , n9644 , n37827 );
and ( n38044 , n38042 , n38043 );
xor ( n38045 , n38042 , n38043 );
xor ( n38046 , n36844 , n36895 );
nor ( n38047 , n9653 , n37827 );
and ( n38048 , n38046 , n38047 );
xor ( n38049 , n38046 , n38047 );
xor ( n38050 , n36848 , n36893 );
nor ( n38051 , n9662 , n37827 );
and ( n38052 , n38050 , n38051 );
xor ( n38053 , n38050 , n38051 );
xor ( n38054 , n36852 , n36891 );
nor ( n38055 , n9671 , n37827 );
and ( n38056 , n38054 , n38055 );
xor ( n38057 , n38054 , n38055 );
xor ( n38058 , n36856 , n36889 );
nor ( n38059 , n9680 , n37827 );
and ( n38060 , n38058 , n38059 );
xor ( n38061 , n38058 , n38059 );
xor ( n38062 , n36860 , n36887 );
nor ( n38063 , n9689 , n37827 );
and ( n38064 , n38062 , n38063 );
xor ( n38065 , n38062 , n38063 );
xor ( n38066 , n36864 , n36885 );
nor ( n38067 , n9698 , n37827 );
and ( n38068 , n38066 , n38067 );
xor ( n38069 , n38066 , n38067 );
xor ( n38070 , n36868 , n36883 );
nor ( n38071 , n9707 , n37827 );
and ( n38072 , n38070 , n38071 );
xor ( n38073 , n38070 , n38071 );
xor ( n38074 , n36872 , n36881 );
nor ( n38075 , n9716 , n37827 );
and ( n38076 , n38074 , n38075 );
xor ( n38077 , n38074 , n38075 );
xor ( n38078 , n36876 , n36879 );
nor ( n38079 , n9725 , n37827 );
and ( n38080 , n38078 , n38079 );
xor ( n38081 , n38078 , n38079 );
xor ( n38082 , n36877 , n36878 );
nor ( n38083 , n9734 , n37827 );
and ( n38084 , n38082 , n38083 );
xor ( n38085 , n38082 , n38083 );
nor ( n38086 , n9752 , n36622 );
nor ( n38087 , n9743 , n37827 );
and ( n38088 , n38086 , n38087 );
and ( n38089 , n38085 , n38088 );
or ( n38090 , n38084 , n38089 );
and ( n38091 , n38081 , n38090 );
or ( n38092 , n38080 , n38091 );
and ( n38093 , n38077 , n38092 );
or ( n38094 , n38076 , n38093 );
and ( n38095 , n38073 , n38094 );
or ( n38096 , n38072 , n38095 );
and ( n38097 , n38069 , n38096 );
or ( n38098 , n38068 , n38097 );
and ( n38099 , n38065 , n38098 );
or ( n38100 , n38064 , n38099 );
and ( n38101 , n38061 , n38100 );
or ( n38102 , n38060 , n38101 );
and ( n38103 , n38057 , n38102 );
or ( n38104 , n38056 , n38103 );
and ( n38105 , n38053 , n38104 );
or ( n38106 , n38052 , n38105 );
and ( n38107 , n38049 , n38106 );
or ( n38108 , n38048 , n38107 );
and ( n38109 , n38045 , n38108 );
or ( n38110 , n38044 , n38109 );
and ( n38111 , n38041 , n38110 );
or ( n38112 , n38040 , n38111 );
and ( n38113 , n38037 , n38112 );
or ( n38114 , n38036 , n38113 );
and ( n38115 , n38033 , n38114 );
or ( n38116 , n38032 , n38115 );
and ( n38117 , n38029 , n38116 );
or ( n38118 , n38028 , n38117 );
and ( n38119 , n38025 , n38118 );
or ( n38120 , n38024 , n38119 );
and ( n38121 , n38021 , n38120 );
or ( n38122 , n38020 , n38121 );
and ( n38123 , n38017 , n38122 );
or ( n38124 , n38016 , n38123 );
and ( n38125 , n38013 , n38124 );
or ( n38126 , n38012 , n38125 );
and ( n38127 , n38009 , n38126 );
or ( n38128 , n38008 , n38127 );
and ( n38129 , n38005 , n38128 );
or ( n38130 , n38004 , n38129 );
and ( n38131 , n38001 , n38130 );
or ( n38132 , n38000 , n38131 );
and ( n38133 , n37997 , n38132 );
or ( n38134 , n37996 , n38133 );
and ( n38135 , n37993 , n38134 );
or ( n38136 , n37992 , n38135 );
and ( n38137 , n37989 , n38136 );
or ( n38138 , n37988 , n38137 );
and ( n38139 , n37985 , n38138 );
or ( n38140 , n37984 , n38139 );
and ( n38141 , n37981 , n38140 );
or ( n38142 , n37980 , n38141 );
and ( n38143 , n37977 , n38142 );
or ( n38144 , n37976 , n38143 );
and ( n38145 , n37973 , n38144 );
or ( n38146 , n37972 , n38145 );
and ( n38147 , n37969 , n38146 );
or ( n38148 , n37968 , n38147 );
and ( n38149 , n37965 , n38148 );
or ( n38150 , n37964 , n38149 );
and ( n38151 , n37961 , n38150 );
or ( n38152 , n37960 , n38151 );
and ( n38153 , n37957 , n38152 );
or ( n38154 , n37956 , n38153 );
and ( n38155 , n37953 , n38154 );
or ( n38156 , n37952 , n38155 );
and ( n38157 , n37949 , n38156 );
or ( n38158 , n37948 , n38157 );
and ( n38159 , n37945 , n38158 );
or ( n38160 , n37944 , n38159 );
and ( n38161 , n37941 , n38160 );
or ( n38162 , n37940 , n38161 );
and ( n38163 , n37937 , n38162 );
or ( n38164 , n37936 , n38163 );
and ( n38165 , n37933 , n38164 );
or ( n38166 , n37932 , n38165 );
and ( n38167 , n37929 , n38166 );
or ( n38168 , n37928 , n38167 );
and ( n38169 , n37925 , n38168 );
or ( n38170 , n37924 , n38169 );
and ( n38171 , n37921 , n38170 );
or ( n38172 , n37920 , n38171 );
and ( n38173 , n37917 , n38172 );
or ( n38174 , n37916 , n38173 );
and ( n38175 , n37913 , n38174 );
or ( n38176 , n37912 , n38175 );
and ( n38177 , n37909 , n38176 );
or ( n38178 , n37908 , n38177 );
and ( n38179 , n37905 , n38178 );
or ( n38180 , n37904 , n38179 );
and ( n38181 , n37901 , n38180 );
or ( n38182 , n37900 , n38181 );
and ( n38183 , n37897 , n38182 );
or ( n38184 , n37896 , n38183 );
and ( n38185 , n37893 , n38184 );
or ( n38186 , n37892 , n38185 );
and ( n38187 , n37889 , n38186 );
or ( n38188 , n37888 , n38187 );
and ( n38189 , n37885 , n38188 );
or ( n38190 , n37884 , n38189 );
and ( n38191 , n37881 , n38190 );
or ( n38192 , n37880 , n38191 );
and ( n38193 , n37877 , n38192 );
or ( n38194 , n37876 , n38193 );
and ( n38195 , n37873 , n38194 );
or ( n38196 , n37872 , n38195 );
and ( n38197 , n37869 , n38196 );
or ( n38198 , n37868 , n38197 );
and ( n38199 , n37865 , n38198 );
or ( n38200 , n37864 , n38199 );
and ( n38201 , n37861 , n38200 );
or ( n38202 , n37860 , n38201 );
and ( n38203 , n37857 , n38202 );
or ( n38204 , n37856 , n38203 );
and ( n38205 , n37853 , n38204 );
or ( n38206 , n37852 , n38205 );
and ( n38207 , n37849 , n38206 );
or ( n38208 , n37848 , n38207 );
and ( n38209 , n37845 , n38208 );
or ( n38210 , n37844 , n38209 );
and ( n38211 , n37841 , n38210 );
or ( n38212 , n37840 , n38211 );
and ( n38213 , n37837 , n38212 );
or ( n38214 , n37836 , n38213 );
and ( n38215 , n37833 , n38214 );
or ( n38216 , n37832 , n38215 );
xor ( n38217 , n37829 , n38216 );
and ( n38218 , n33403 , n683 );
nor ( n38219 , n684 , n38218 );
nor ( n38220 , n733 , n32231 );
xor ( n38221 , n38219 , n38220 );
and ( n38222 , n37008 , n37009 );
and ( n38223 , n37010 , n37012 );
or ( n38224 , n38222 , n38223 );
xor ( n38225 , n38221 , n38224 );
nor ( n38226 , n796 , n31083 );
xor ( n38227 , n38225 , n38226 );
and ( n38228 , n37013 , n37014 );
and ( n38229 , n37015 , n37018 );
or ( n38230 , n38228 , n38229 );
xor ( n38231 , n38227 , n38230 );
nor ( n38232 , n868 , n29948 );
xor ( n38233 , n38231 , n38232 );
and ( n38234 , n37019 , n37020 );
and ( n38235 , n37021 , n37024 );
or ( n38236 , n38234 , n38235 );
xor ( n38237 , n38233 , n38236 );
nor ( n38238 , n958 , n28833 );
xor ( n38239 , n38237 , n38238 );
and ( n38240 , n37025 , n37026 );
and ( n38241 , n37027 , n37030 );
or ( n38242 , n38240 , n38241 );
xor ( n38243 , n38239 , n38242 );
nor ( n38244 , n1062 , n27737 );
xor ( n38245 , n38243 , n38244 );
and ( n38246 , n37031 , n37032 );
and ( n38247 , n37033 , n37036 );
or ( n38248 , n38246 , n38247 );
xor ( n38249 , n38245 , n38248 );
nor ( n38250 , n1176 , n26660 );
xor ( n38251 , n38249 , n38250 );
and ( n38252 , n37037 , n37038 );
and ( n38253 , n37039 , n37042 );
or ( n38254 , n38252 , n38253 );
xor ( n38255 , n38251 , n38254 );
nor ( n38256 , n1303 , n25600 );
xor ( n38257 , n38255 , n38256 );
and ( n38258 , n37043 , n37044 );
and ( n38259 , n37045 , n37048 );
or ( n38260 , n38258 , n38259 );
xor ( n38261 , n38257 , n38260 );
nor ( n38262 , n1445 , n24564 );
xor ( n38263 , n38261 , n38262 );
and ( n38264 , n37049 , n37050 );
and ( n38265 , n37051 , n37054 );
or ( n38266 , n38264 , n38265 );
xor ( n38267 , n38263 , n38266 );
nor ( n38268 , n1598 , n23541 );
xor ( n38269 , n38267 , n38268 );
and ( n38270 , n37055 , n37056 );
and ( n38271 , n37057 , n37060 );
or ( n38272 , n38270 , n38271 );
xor ( n38273 , n38269 , n38272 );
nor ( n38274 , n1766 , n22541 );
xor ( n38275 , n38273 , n38274 );
and ( n38276 , n37061 , n37062 );
and ( n38277 , n37063 , n37066 );
or ( n38278 , n38276 , n38277 );
xor ( n38279 , n38275 , n38278 );
nor ( n38280 , n1945 , n21562 );
xor ( n38281 , n38279 , n38280 );
and ( n38282 , n37067 , n37068 );
and ( n38283 , n37069 , n37072 );
or ( n38284 , n38282 , n38283 );
xor ( n38285 , n38281 , n38284 );
nor ( n38286 , n2137 , n20601 );
xor ( n38287 , n38285 , n38286 );
and ( n38288 , n37073 , n37074 );
and ( n38289 , n37075 , n37078 );
or ( n38290 , n38288 , n38289 );
xor ( n38291 , n38287 , n38290 );
nor ( n38292 , n2343 , n19657 );
xor ( n38293 , n38291 , n38292 );
and ( n38294 , n37079 , n37080 );
and ( n38295 , n37081 , n37084 );
or ( n38296 , n38294 , n38295 );
xor ( n38297 , n38293 , n38296 );
nor ( n38298 , n2566 , n18734 );
xor ( n38299 , n38297 , n38298 );
and ( n38300 , n37085 , n37086 );
and ( n38301 , n37087 , n37090 );
or ( n38302 , n38300 , n38301 );
xor ( n38303 , n38299 , n38302 );
nor ( n38304 , n2797 , n17828 );
xor ( n38305 , n38303 , n38304 );
and ( n38306 , n37091 , n37092 );
and ( n38307 , n37093 , n37096 );
or ( n38308 , n38306 , n38307 );
xor ( n38309 , n38305 , n38308 );
nor ( n38310 , n3043 , n16943 );
xor ( n38311 , n38309 , n38310 );
and ( n38312 , n37097 , n37098 );
and ( n38313 , n37099 , n37102 );
or ( n38314 , n38312 , n38313 );
xor ( n38315 , n38311 , n38314 );
nor ( n38316 , n3300 , n16077 );
xor ( n38317 , n38315 , n38316 );
and ( n38318 , n37103 , n37104 );
and ( n38319 , n37105 , n37108 );
or ( n38320 , n38318 , n38319 );
xor ( n38321 , n38317 , n38320 );
nor ( n38322 , n3570 , n15230 );
xor ( n38323 , n38321 , n38322 );
and ( n38324 , n37109 , n37110 );
and ( n38325 , n37111 , n37114 );
or ( n38326 , n38324 , n38325 );
xor ( n38327 , n38323 , n38326 );
nor ( n38328 , n3853 , n14403 );
xor ( n38329 , n38327 , n38328 );
and ( n38330 , n37115 , n37116 );
and ( n38331 , n37117 , n37120 );
or ( n38332 , n38330 , n38331 );
xor ( n38333 , n38329 , n38332 );
nor ( n38334 , n4151 , n13599 );
xor ( n38335 , n38333 , n38334 );
and ( n38336 , n37121 , n37122 );
and ( n38337 , n37123 , n37126 );
or ( n38338 , n38336 , n38337 );
xor ( n38339 , n38335 , n38338 );
nor ( n38340 , n4458 , n12808 );
xor ( n38341 , n38339 , n38340 );
and ( n38342 , n37127 , n37128 );
and ( n38343 , n37129 , n37132 );
or ( n38344 , n38342 , n38343 );
xor ( n38345 , n38341 , n38344 );
nor ( n38346 , n4786 , n12037 );
xor ( n38347 , n38345 , n38346 );
and ( n38348 , n37133 , n37134 );
and ( n38349 , n37135 , n37138 );
or ( n38350 , n38348 , n38349 );
xor ( n38351 , n38347 , n38350 );
nor ( n38352 , n5126 , n11282 );
xor ( n38353 , n38351 , n38352 );
and ( n38354 , n37139 , n37140 );
and ( n38355 , n37141 , n37144 );
or ( n38356 , n38354 , n38355 );
xor ( n38357 , n38353 , n38356 );
nor ( n38358 , n5477 , n10547 );
xor ( n38359 , n38357 , n38358 );
and ( n38360 , n37145 , n37146 );
and ( n38361 , n37147 , n37150 );
or ( n38362 , n38360 , n38361 );
xor ( n38363 , n38359 , n38362 );
nor ( n38364 , n5838 , n9829 );
xor ( n38365 , n38363 , n38364 );
and ( n38366 , n37151 , n37152 );
and ( n38367 , n37153 , n37156 );
or ( n38368 , n38366 , n38367 );
xor ( n38369 , n38365 , n38368 );
nor ( n38370 , n6212 , n8955 );
xor ( n38371 , n38369 , n38370 );
and ( n38372 , n37157 , n37158 );
and ( n38373 , n37159 , n37162 );
or ( n38374 , n38372 , n38373 );
xor ( n38375 , n38371 , n38374 );
nor ( n38376 , n6596 , n603 );
xor ( n38377 , n38375 , n38376 );
and ( n38378 , n37163 , n37164 );
and ( n38379 , n37165 , n37168 );
or ( n38380 , n38378 , n38379 );
xor ( n38381 , n38377 , n38380 );
nor ( n38382 , n6997 , n652 );
xor ( n38383 , n38381 , n38382 );
and ( n38384 , n37169 , n37170 );
and ( n38385 , n37171 , n37174 );
or ( n38386 , n38384 , n38385 );
xor ( n38387 , n38383 , n38386 );
nor ( n38388 , n7413 , n624 );
xor ( n38389 , n38387 , n38388 );
and ( n38390 , n37175 , n37176 );
and ( n38391 , n37177 , n37180 );
or ( n38392 , n38390 , n38391 );
xor ( n38393 , n38389 , n38392 );
nor ( n38394 , n7841 , n648 );
xor ( n38395 , n38393 , n38394 );
and ( n38396 , n37181 , n37182 );
and ( n38397 , n37183 , n37186 );
or ( n38398 , n38396 , n38397 );
xor ( n38399 , n38395 , n38398 );
nor ( n38400 , n8281 , n686 );
xor ( n38401 , n38399 , n38400 );
and ( n38402 , n37187 , n37188 );
and ( n38403 , n37189 , n37192 );
or ( n38404 , n38402 , n38403 );
xor ( n38405 , n38401 , n38404 );
nor ( n38406 , n8737 , n735 );
xor ( n38407 , n38405 , n38406 );
and ( n38408 , n37193 , n37194 );
and ( n38409 , n37195 , n37198 );
or ( n38410 , n38408 , n38409 );
xor ( n38411 , n38407 , n38410 );
nor ( n38412 , n9420 , n798 );
xor ( n38413 , n38411 , n38412 );
and ( n38414 , n37199 , n37200 );
and ( n38415 , n37201 , n37204 );
or ( n38416 , n38414 , n38415 );
xor ( n38417 , n38413 , n38416 );
nor ( n38418 , n10312 , n870 );
xor ( n38419 , n38417 , n38418 );
and ( n38420 , n37205 , n37206 );
and ( n38421 , n37207 , n37210 );
or ( n38422 , n38420 , n38421 );
xor ( n38423 , n38419 , n38422 );
nor ( n38424 , n11041 , n960 );
xor ( n38425 , n38423 , n38424 );
and ( n38426 , n37211 , n37212 );
and ( n38427 , n37213 , n37216 );
or ( n38428 , n38426 , n38427 );
xor ( n38429 , n38425 , n38428 );
nor ( n38430 , n11790 , n1064 );
xor ( n38431 , n38429 , n38430 );
and ( n38432 , n37217 , n37218 );
and ( n38433 , n37219 , n37222 );
or ( n38434 , n38432 , n38433 );
xor ( n38435 , n38431 , n38434 );
nor ( n38436 , n12555 , n1178 );
xor ( n38437 , n38435 , n38436 );
and ( n38438 , n37223 , n37224 );
and ( n38439 , n37225 , n37228 );
or ( n38440 , n38438 , n38439 );
xor ( n38441 , n38437 , n38440 );
nor ( n38442 , n13340 , n1305 );
xor ( n38443 , n38441 , n38442 );
and ( n38444 , n37229 , n37230 );
and ( n38445 , n37231 , n37234 );
or ( n38446 , n38444 , n38445 );
xor ( n38447 , n38443 , n38446 );
nor ( n38448 , n14138 , n1447 );
xor ( n38449 , n38447 , n38448 );
and ( n38450 , n37235 , n37236 );
and ( n38451 , n37237 , n37240 );
or ( n38452 , n38450 , n38451 );
xor ( n38453 , n38449 , n38452 );
nor ( n38454 , n14959 , n1600 );
xor ( n38455 , n38453 , n38454 );
and ( n38456 , n37241 , n37242 );
and ( n38457 , n37243 , n37246 );
or ( n38458 , n38456 , n38457 );
xor ( n38459 , n38455 , n38458 );
nor ( n38460 , n15800 , n1768 );
xor ( n38461 , n38459 , n38460 );
and ( n38462 , n37247 , n37248 );
and ( n38463 , n37249 , n37252 );
or ( n38464 , n38462 , n38463 );
xor ( n38465 , n38461 , n38464 );
nor ( n38466 , n16660 , n1947 );
xor ( n38467 , n38465 , n38466 );
and ( n38468 , n37253 , n37254 );
and ( n38469 , n37255 , n37258 );
or ( n38470 , n38468 , n38469 );
xor ( n38471 , n38467 , n38470 );
nor ( n38472 , n17539 , n2139 );
xor ( n38473 , n38471 , n38472 );
and ( n38474 , n37259 , n37260 );
and ( n38475 , n37261 , n37264 );
or ( n38476 , n38474 , n38475 );
xor ( n38477 , n38473 , n38476 );
nor ( n38478 , n18439 , n2345 );
xor ( n38479 , n38477 , n38478 );
and ( n38480 , n37265 , n37266 );
and ( n38481 , n37267 , n37270 );
or ( n38482 , n38480 , n38481 );
xor ( n38483 , n38479 , n38482 );
nor ( n38484 , n19356 , n2568 );
xor ( n38485 , n38483 , n38484 );
and ( n38486 , n37271 , n37272 );
and ( n38487 , n37273 , n37276 );
or ( n38488 , n38486 , n38487 );
xor ( n38489 , n38485 , n38488 );
nor ( n38490 , n20294 , n2799 );
xor ( n38491 , n38489 , n38490 );
and ( n38492 , n37277 , n37278 );
and ( n38493 , n37279 , n37282 );
or ( n38494 , n38492 , n38493 );
xor ( n38495 , n38491 , n38494 );
nor ( n38496 , n21249 , n3045 );
xor ( n38497 , n38495 , n38496 );
and ( n38498 , n37283 , n37284 );
and ( n38499 , n37285 , n37288 );
or ( n38500 , n38498 , n38499 );
xor ( n38501 , n38497 , n38500 );
nor ( n38502 , n22222 , n3302 );
xor ( n38503 , n38501 , n38502 );
and ( n38504 , n37289 , n37290 );
and ( n38505 , n37291 , n37294 );
or ( n38506 , n38504 , n38505 );
xor ( n38507 , n38503 , n38506 );
nor ( n38508 , n23216 , n3572 );
xor ( n38509 , n38507 , n38508 );
and ( n38510 , n37295 , n37296 );
and ( n38511 , n37297 , n37300 );
or ( n38512 , n38510 , n38511 );
xor ( n38513 , n38509 , n38512 );
nor ( n38514 , n24233 , n3855 );
xor ( n38515 , n38513 , n38514 );
and ( n38516 , n37301 , n37302 );
and ( n38517 , n37303 , n37306 );
or ( n38518 , n38516 , n38517 );
xor ( n38519 , n38515 , n38518 );
nor ( n38520 , n25263 , n4153 );
xor ( n38521 , n38519 , n38520 );
and ( n38522 , n37307 , n37308 );
and ( n38523 , n37309 , n37312 );
or ( n38524 , n38522 , n38523 );
xor ( n38525 , n38521 , n38524 );
nor ( n38526 , n26317 , n4460 );
xor ( n38527 , n38525 , n38526 );
and ( n38528 , n37313 , n37314 );
and ( n38529 , n37315 , n37318 );
or ( n38530 , n38528 , n38529 );
xor ( n38531 , n38527 , n38530 );
nor ( n38532 , n27388 , n4788 );
xor ( n38533 , n38531 , n38532 );
and ( n38534 , n37319 , n37320 );
and ( n38535 , n37321 , n37324 );
or ( n38536 , n38534 , n38535 );
xor ( n38537 , n38533 , n38536 );
nor ( n38538 , n28478 , n5128 );
xor ( n38539 , n38537 , n38538 );
and ( n38540 , n37325 , n37326 );
and ( n38541 , n37327 , n37330 );
or ( n38542 , n38540 , n38541 );
xor ( n38543 , n38539 , n38542 );
nor ( n38544 , n29587 , n5479 );
xor ( n38545 , n38543 , n38544 );
and ( n38546 , n37331 , n37332 );
and ( n38547 , n37333 , n37336 );
or ( n38548 , n38546 , n38547 );
xor ( n38549 , n38545 , n38548 );
nor ( n38550 , n30716 , n5840 );
xor ( n38551 , n38549 , n38550 );
and ( n38552 , n37337 , n37338 );
and ( n38553 , n37339 , n37342 );
or ( n38554 , n38552 , n38553 );
xor ( n38555 , n38551 , n38554 );
nor ( n38556 , n31858 , n6214 );
xor ( n38557 , n38555 , n38556 );
and ( n38558 , n37343 , n37344 );
and ( n38559 , n37345 , n37348 );
or ( n38560 , n38558 , n38559 );
xor ( n38561 , n38557 , n38560 );
nor ( n38562 , n33024 , n6598 );
xor ( n38563 , n38561 , n38562 );
and ( n38564 , n37349 , n37350 );
and ( n38565 , n37351 , n37354 );
or ( n38566 , n38564 , n38565 );
xor ( n38567 , n38563 , n38566 );
nor ( n38568 , n34215 , n6999 );
xor ( n38569 , n38567 , n38568 );
and ( n38570 , n37355 , n37356 );
and ( n38571 , n37357 , n37360 );
or ( n38572 , n38570 , n38571 );
xor ( n38573 , n38569 , n38572 );
nor ( n38574 , n35410 , n7415 );
xor ( n38575 , n38573 , n38574 );
and ( n38576 , n37361 , n37362 );
and ( n38577 , n37363 , n37366 );
or ( n38578 , n38576 , n38577 );
xor ( n38579 , n38575 , n38578 );
nor ( n38580 , n36611 , n7843 );
xor ( n38581 , n38579 , n38580 );
and ( n38582 , n37367 , n37368 );
and ( n38583 , n37369 , n37372 );
or ( n38584 , n38582 , n38583 );
xor ( n38585 , n38581 , n38584 );
nor ( n38586 , n37816 , n8283 );
xor ( n38587 , n38585 , n38586 );
and ( n38588 , n37373 , n37374 );
and ( n38589 , n37375 , n37378 );
or ( n38590 , n38588 , n38589 );
xor ( n38591 , n38587 , n38590 );
and ( n38592 , n37391 , n37395 );
and ( n38593 , n37395 , n37802 );
and ( n38594 , n37391 , n37802 );
or ( n38595 , n38592 , n38593 , n38594 );
and ( n38596 , n33774 , n663 );
not ( n38597 , n663 );
nor ( n38598 , n38596 , n38597 );
xor ( n38599 , n38595 , n38598 );
and ( n38600 , n37404 , n37408 );
and ( n38601 , n37408 , n37476 );
and ( n38602 , n37404 , n37476 );
or ( n38603 , n38600 , n38601 , n38602 );
and ( n38604 , n37400 , n37477 );
and ( n38605 , n37477 , n37801 );
and ( n38606 , n37400 , n37801 );
or ( n38607 , n38604 , n38605 , n38606 );
xor ( n38608 , n38603 , n38607 );
and ( n38609 , n37482 , n37602 );
and ( n38610 , n37602 , n37800 );
and ( n38611 , n37482 , n37800 );
or ( n38612 , n38609 , n38610 , n38611 );
and ( n38613 , n37413 , n37417 );
and ( n38614 , n37417 , n37475 );
and ( n38615 , n37413 , n37475 );
or ( n38616 , n38613 , n38614 , n38615 );
and ( n38617 , n37486 , n37490 );
and ( n38618 , n37490 , n37601 );
and ( n38619 , n37486 , n37601 );
or ( n38620 , n38617 , n38618 , n38619 );
xor ( n38621 , n38616 , n38620 );
and ( n38622 , n37444 , n37448 );
and ( n38623 , n37448 , n37454 );
and ( n38624 , n37444 , n37454 );
or ( n38625 , n38622 , n38623 , n38624 );
and ( n38626 , n37422 , n37426 );
and ( n38627 , n37426 , n37474 );
and ( n38628 , n37422 , n37474 );
or ( n38629 , n38626 , n38627 , n38628 );
xor ( n38630 , n38625 , n38629 );
and ( n38631 , n37431 , n37435 );
and ( n38632 , n37435 , n37473 );
and ( n38633 , n37431 , n37473 );
or ( n38634 , n38631 , n38632 , n38633 );
and ( n38635 , n37499 , n37524 );
and ( n38636 , n37524 , n37562 );
and ( n38637 , n37499 , n37562 );
or ( n38638 , n38635 , n38636 , n38637 );
xor ( n38639 , n38634 , n38638 );
and ( n38640 , n37440 , n37455 );
and ( n38641 , n37455 , n37472 );
and ( n38642 , n37440 , n37472 );
or ( n38643 , n38640 , n38641 , n38642 );
and ( n38644 , n37503 , n37507 );
and ( n38645 , n37507 , n37523 );
and ( n38646 , n37503 , n37523 );
or ( n38647 , n38644 , n38645 , n38646 );
xor ( n38648 , n38643 , n38647 );
and ( n38649 , n37460 , n37465 );
and ( n38650 , n37465 , n37471 );
and ( n38651 , n37460 , n37471 );
or ( n38652 , n38649 , n38650 , n38651 );
and ( n38653 , n37450 , n37451 );
and ( n38654 , n37451 , n37453 );
and ( n38655 , n37450 , n37453 );
or ( n38656 , n38653 , n38654 , n38655 );
and ( n38657 , n37461 , n37462 );
and ( n38658 , n37462 , n37464 );
and ( n38659 , n37461 , n37464 );
or ( n38660 , n38657 , n38658 , n38659 );
xor ( n38661 , n38656 , n38660 );
and ( n38662 , n30695 , n840 );
and ( n38663 , n31836 , n771 );
xor ( n38664 , n38662 , n38663 );
and ( n38665 , n32649 , n719 );
xor ( n38666 , n38664 , n38665 );
xor ( n38667 , n38661 , n38666 );
xor ( n38668 , n38652 , n38667 );
and ( n38669 , n37467 , n37468 );
and ( n38670 , n37468 , n37470 );
and ( n38671 , n37467 , n37470 );
or ( n38672 , n38669 , n38670 , n38671 );
and ( n38673 , n27361 , n1134 );
and ( n38674 , n28456 , n1034 );
xor ( n38675 , n38673 , n38674 );
and ( n38676 , n29559 , n940 );
xor ( n38677 , n38675 , n38676 );
xor ( n38678 , n38672 , n38677 );
and ( n38679 , n24214 , n1551 );
and ( n38680 , n25243 , n1424 );
xor ( n38681 , n38679 , n38680 );
and ( n38682 , n26296 , n1254 );
xor ( n38683 , n38681 , n38682 );
xor ( n38684 , n38678 , n38683 );
xor ( n38685 , n38668 , n38684 );
xor ( n38686 , n38648 , n38685 );
xor ( n38687 , n38639 , n38686 );
xor ( n38688 , n38630 , n38687 );
xor ( n38689 , n38621 , n38688 );
xor ( n38690 , n38612 , n38689 );
and ( n38691 , n37607 , n37685 );
and ( n38692 , n37685 , n37799 );
and ( n38693 , n37607 , n37799 );
or ( n38694 , n38691 , n38692 , n38693 );
and ( n38695 , n37495 , n37563 );
and ( n38696 , n37563 , n37600 );
and ( n38697 , n37495 , n37600 );
or ( n38698 , n38695 , n38696 , n38697 );
and ( n38699 , n37611 , n37615 );
and ( n38700 , n37615 , n37684 );
and ( n38701 , n37611 , n37684 );
or ( n38702 , n38699 , n38700 , n38701 );
xor ( n38703 , n38698 , n38702 );
and ( n38704 , n37568 , n37572 );
and ( n38705 , n37572 , n37599 );
and ( n38706 , n37568 , n37599 );
or ( n38707 , n38704 , n38705 , n38706 );
and ( n38708 , n37529 , n37545 );
and ( n38709 , n37545 , n37561 );
and ( n38710 , n37529 , n37561 );
or ( n38711 , n38708 , n38709 , n38710 );
and ( n38712 , n37512 , n37516 );
and ( n38713 , n37516 , n37522 );
and ( n38714 , n37512 , n37522 );
or ( n38715 , n38712 , n38713 , n38714 );
and ( n38716 , n37533 , n37538 );
and ( n38717 , n37538 , n37544 );
and ( n38718 , n37533 , n37544 );
or ( n38719 , n38716 , n38717 , n38718 );
xor ( n38720 , n38715 , n38719 );
and ( n38721 , n37518 , n37519 );
and ( n38722 , n37519 , n37521 );
and ( n38723 , n37518 , n37521 );
or ( n38724 , n38721 , n38722 , n38723 );
and ( n38725 , n37534 , n37535 );
and ( n38726 , n37535 , n37537 );
and ( n38727 , n37534 , n37537 );
or ( n38728 , n38725 , n38726 , n38727 );
xor ( n38729 , n38724 , n38728 );
and ( n38730 , n21216 , n2100 );
and ( n38731 , n22186 , n1882 );
xor ( n38732 , n38730 , n38731 );
and ( n38733 , n22892 , n1738 );
xor ( n38734 , n38732 , n38733 );
xor ( n38735 , n38729 , n38734 );
xor ( n38736 , n38720 , n38735 );
xor ( n38737 , n38711 , n38736 );
and ( n38738 , n37550 , n37554 );
and ( n38739 , n37554 , n37560 );
and ( n38740 , n37550 , n37560 );
or ( n38741 , n38738 , n38739 , n38740 );
and ( n38742 , n37540 , n37541 );
and ( n38743 , n37541 , n37543 );
and ( n38744 , n37540 , n37543 );
or ( n38745 , n38742 , n38743 , n38744 );
and ( n38746 , n18144 , n2739 );
and ( n38747 , n19324 , n2544 );
xor ( n38748 , n38746 , n38747 );
and ( n38749 , n20233 , n2298 );
xor ( n38750 , n38748 , n38749 );
xor ( n38751 , n38745 , n38750 );
and ( n38752 , n15758 , n3495 );
and ( n38753 , n16637 , n3271 );
xor ( n38754 , n38752 , n38753 );
and ( n38755 , n17512 , n2981 );
xor ( n38756 , n38754 , n38755 );
xor ( n38757 , n38751 , n38756 );
xor ( n38758 , n38741 , n38757 );
and ( n38759 , n37556 , n37557 );
and ( n38760 , n37557 , n37559 );
and ( n38761 , n37556 , n37559 );
or ( n38762 , n38759 , n38760 , n38761 );
and ( n38763 , n37587 , n37588 );
and ( n38764 , n37588 , n37590 );
and ( n38765 , n37587 , n37590 );
or ( n38766 , n38763 , n38764 , n38765 );
xor ( n38767 , n38762 , n38766 );
and ( n38768 , n13322 , n4403 );
and ( n38769 , n14118 , n4102 );
xor ( n38770 , n38768 , n38769 );
and ( n38771 , n14938 , n3749 );
xor ( n38772 , n38770 , n38771 );
xor ( n38773 , n38767 , n38772 );
xor ( n38774 , n38758 , n38773 );
xor ( n38775 , n38737 , n38774 );
xor ( n38776 , n38707 , n38775 );
and ( n38777 , n37577 , n37581 );
and ( n38778 , n37581 , n37598 );
and ( n38779 , n37577 , n37598 );
or ( n38780 , n38777 , n38778 , n38779 );
and ( n38781 , n37624 , n37639 );
and ( n38782 , n37639 , n37656 );
and ( n38783 , n37624 , n37656 );
or ( n38784 , n38781 , n38782 , n38783 );
xor ( n38785 , n38780 , n38784 );
and ( n38786 , n37586 , n37591 );
and ( n38787 , n37591 , n37597 );
and ( n38788 , n37586 , n37597 );
or ( n38789 , n38786 , n38787 , n38788 );
and ( n38790 , n37628 , n37632 );
and ( n38791 , n37632 , n37638 );
and ( n38792 , n37628 , n37638 );
or ( n38793 , n38790 , n38791 , n38792 );
xor ( n38794 , n38789 , n38793 );
and ( n38795 , n37593 , n37594 );
and ( n38796 , n37594 , n37596 );
and ( n38797 , n37593 , n37596 );
or ( n38798 , n38795 , n38796 , n38797 );
and ( n38799 , n11015 , n5408 );
and ( n38800 , n11769 , n5103 );
xor ( n38801 , n38799 , n38800 );
and ( n38802 , n12320 , n4730 );
xor ( n38803 , n38801 , n38802 );
xor ( n38804 , n38798 , n38803 );
and ( n38805 , n8718 , n6504 );
and ( n38806 , n9400 , n6132 );
xor ( n38807 , n38805 , n38806 );
and ( n38808 , n10291 , n5765 );
xor ( n38809 , n38807 , n38808 );
xor ( n38810 , n38804 , n38809 );
xor ( n38811 , n38794 , n38810 );
xor ( n38812 , n38785 , n38811 );
xor ( n38813 , n38776 , n38812 );
xor ( n38814 , n38703 , n38813 );
xor ( n38815 , n38694 , n38814 );
and ( n38816 , n37690 , n37737 );
and ( n38817 , n37737 , n37798 );
and ( n38818 , n37690 , n37798 );
or ( n38819 , n38816 , n38817 , n38818 );
and ( n38820 , n37620 , n37657 );
and ( n38821 , n37657 , n37683 );
and ( n38822 , n37620 , n37683 );
or ( n38823 , n38820 , n38821 , n38822 );
and ( n38824 , n37694 , n37698 );
and ( n38825 , n37698 , n37736 );
and ( n38826 , n37694 , n37736 );
or ( n38827 , n38824 , n38825 , n38826 );
xor ( n38828 , n38823 , n38827 );
and ( n38829 , n37662 , n37666 );
and ( n38830 , n37666 , n37682 );
and ( n38831 , n37662 , n37682 );
or ( n38832 , n38829 , n38830 , n38831 );
and ( n38833 , n37644 , n37649 );
and ( n38834 , n37649 , n37655 );
and ( n38835 , n37644 , n37655 );
or ( n38836 , n38833 , n38834 , n38835 );
and ( n38837 , n37634 , n37635 );
and ( n38838 , n37635 , n37637 );
and ( n38839 , n37634 , n37637 );
or ( n38840 , n38837 , n38838 , n38839 );
and ( n38841 , n37645 , n37646 );
and ( n38842 , n37646 , n37648 );
and ( n38843 , n37645 , n37648 );
or ( n38844 , n38841 , n38842 , n38843 );
xor ( n38845 , n38840 , n38844 );
and ( n38846 , n8079 , n6971 );
buf ( n38847 , n38846 );
xor ( n38848 , n38845 , n38847 );
xor ( n38849 , n38836 , n38848 );
and ( n38850 , n37651 , n37652 );
and ( n38851 , n37652 , n37654 );
and ( n38852 , n37651 , n37654 );
or ( n38853 , n38850 , n38851 , n38852 );
and ( n38854 , n6187 , n9348 );
and ( n38855 , n6569 , n8669 );
xor ( n38856 , n38854 , n38855 );
and ( n38857 , n6816 , n8243 );
xor ( n38858 , n38856 , n38857 );
xor ( n38859 , n38853 , n38858 );
and ( n38860 , n4959 , n11718 );
and ( n38861 , n5459 , n10977 );
xor ( n38862 , n38860 , n38861 );
and ( n38863 , n5819 , n10239 );
xor ( n38864 , n38862 , n38863 );
xor ( n38865 , n38859 , n38864 );
xor ( n38866 , n38849 , n38865 );
xor ( n38867 , n38832 , n38866 );
and ( n38868 , n37671 , n37675 );
and ( n38869 , n37675 , n37681 );
and ( n38870 , n37671 , n37681 );
or ( n38871 , n38868 , n38869 , n38870 );
and ( n38872 , n37707 , n37712 );
and ( n38873 , n37712 , n37718 );
and ( n38874 , n37707 , n37718 );
or ( n38875 , n38872 , n38873 , n38874 );
xor ( n38876 , n38871 , n38875 );
and ( n38877 , n37677 , n37678 );
and ( n38878 , n37678 , n37680 );
and ( n38879 , n37677 , n37680 );
or ( n38880 , n38877 , n38878 , n38879 );
and ( n38881 , n37708 , n37709 );
and ( n38882 , n37709 , n37711 );
and ( n38883 , n37708 , n37711 );
or ( n38884 , n38881 , n38882 , n38883 );
xor ( n38885 , n38880 , n38884 );
and ( n38886 , n4132 , n14044 );
and ( n38887 , n4438 , n13256 );
xor ( n38888 , n38886 , n38887 );
and ( n38889 , n4766 , n12531 );
xor ( n38890 , n38888 , n38889 );
xor ( n38891 , n38885 , n38890 );
xor ( n38892 , n38876 , n38891 );
xor ( n38893 , n38867 , n38892 );
xor ( n38894 , n38828 , n38893 );
xor ( n38895 , n38819 , n38894 );
and ( n38896 , n37742 , n37768 );
and ( n38897 , n37768 , n37797 );
and ( n38898 , n37742 , n37797 );
or ( n38899 , n38896 , n38897 , n38898 );
and ( n38900 , n37703 , n37719 );
and ( n38901 , n37719 , n37735 );
and ( n38902 , n37703 , n37735 );
or ( n38903 , n38900 , n38901 , n38902 );
and ( n38904 , n37746 , n37750 );
and ( n38905 , n37750 , n37767 );
and ( n38906 , n37746 , n37767 );
or ( n38907 , n38904 , n38905 , n38906 );
xor ( n38908 , n38903 , n38907 );
and ( n38909 , n37724 , n37728 );
and ( n38910 , n37728 , n37734 );
and ( n38911 , n37724 , n37734 );
or ( n38912 , n38909 , n38910 , n38911 );
and ( n38913 , n37714 , n37715 );
and ( n38914 , n37715 , n37717 );
and ( n38915 , n37714 , n37717 );
or ( n38916 , n38913 , n38914 , n38915 );
and ( n38917 , n3182 , n16550 );
and ( n38918 , n3545 , n15691 );
xor ( n38919 , n38917 , n38918 );
and ( n38920 , n3801 , n14838 );
xor ( n38921 , n38919 , n38920 );
xor ( n38922 , n38916 , n38921 );
and ( n38923 , n2462 , n19222 );
and ( n38924 , n2779 , n18407 );
xor ( n38925 , n38923 , n38924 );
and ( n38926 , n3024 , n17422 );
xor ( n38927 , n38925 , n38926 );
xor ( n38928 , n38922 , n38927 );
xor ( n38929 , n38912 , n38928 );
and ( n38930 , n37730 , n37731 );
and ( n38931 , n37731 , n37733 );
and ( n38932 , n37730 , n37733 );
or ( n38933 , n38930 , n38931 , n38932 );
and ( n38934 , n37756 , n37757 );
and ( n38935 , n37757 , n37759 );
and ( n38936 , n37756 , n37759 );
or ( n38937 , n38934 , n38935 , n38936 );
xor ( n38938 , n38933 , n38937 );
and ( n38939 , n1933 , n22065 );
and ( n38940 , n2120 , n20976 );
xor ( n38941 , n38939 , n38940 );
and ( n38942 , n2324 , n20156 );
xor ( n38943 , n38941 , n38942 );
xor ( n38944 , n38938 , n38943 );
xor ( n38945 , n38929 , n38944 );
xor ( n38946 , n38908 , n38945 );
xor ( n38947 , n38899 , n38946 );
and ( n38948 , n37773 , n37780 );
and ( n38949 , n37780 , n37796 );
and ( n38950 , n37773 , n37796 );
or ( n38951 , n38948 , n38949 , n38950 );
and ( n38952 , n37755 , n37760 );
and ( n38953 , n37760 , n37766 );
and ( n38954 , n37755 , n37766 );
or ( n38955 , n38952 , n38953 , n38954 );
and ( n38956 , n37785 , n37789 );
and ( n38957 , n37789 , n37795 );
and ( n38958 , n37785 , n37795 );
or ( n38959 , n38956 , n38957 , n38958 );
xor ( n38960 , n38955 , n38959 );
and ( n38961 , n37762 , n37763 );
and ( n38962 , n37763 , n37765 );
and ( n38963 , n37762 , n37765 );
or ( n38964 , n38961 , n38962 , n38963 );
and ( n38965 , n1383 , n25163 );
and ( n38966 , n1580 , n24137 );
xor ( n38967 , n38965 , n38966 );
and ( n38968 , n1694 , n23075 );
xor ( n38969 , n38967 , n38968 );
xor ( n38970 , n38964 , n38969 );
and ( n38971 , n1047 , n28406 );
and ( n38972 , n1164 , n27296 );
xor ( n38973 , n38971 , n38972 );
and ( n38974 , n1287 , n26216 );
xor ( n38975 , n38973 , n38974 );
xor ( n38976 , n38970 , n38975 );
xor ( n38977 , n38960 , n38976 );
xor ( n38978 , n38951 , n38977 );
and ( n38979 , n37776 , n37777 );
and ( n38980 , n37777 , n37779 );
and ( n38981 , n37776 , n37779 );
or ( n38982 , n38979 , n38980 , n38981 );
and ( n38983 , n37791 , n37792 );
and ( n38984 , n37792 , n37794 );
and ( n38985 , n37791 , n37794 );
or ( n38986 , n38983 , n38984 , n38985 );
xor ( n38987 , n38982 , n38986 );
and ( n38988 , n783 , n31761 );
and ( n38989 , n856 , n30629 );
xor ( n38990 , n38988 , n38989 );
and ( n38991 , n925 , n29508 );
xor ( n38992 , n38990 , n38991 );
xor ( n38993 , n38987 , n38992 );
not ( n38994 , n671 );
and ( n38995 , n34193 , n671 );
nor ( n38996 , n38994 , n38995 );
and ( n38997 , n715 , n32999 );
xor ( n38998 , n38996 , n38997 );
xor ( n38999 , n38993 , n38998 );
xor ( n39000 , n38978 , n38999 );
xor ( n39001 , n38947 , n39000 );
xor ( n39002 , n38895 , n39001 );
xor ( n39003 , n38815 , n39002 );
xor ( n39004 , n38690 , n39003 );
xor ( n39005 , n38608 , n39004 );
xor ( n39006 , n38599 , n39005 );
and ( n39007 , n37383 , n37386 );
and ( n39008 , n37386 , n37803 );
and ( n39009 , n37383 , n37803 );
or ( n39010 , n39007 , n39008 , n39009 );
xor ( n39011 , n39006 , n39010 );
and ( n39012 , n37804 , n37808 );
and ( n39013 , n37809 , n37812 );
or ( n39014 , n39012 , n39013 );
xor ( n39015 , n39011 , n39014 );
buf ( n39016 , n39015 );
buf ( n39017 , n39016 );
not ( n39018 , n39017 );
nor ( n39019 , n39018 , n8739 );
xor ( n39020 , n38591 , n39019 );
and ( n39021 , n37379 , n37817 );
and ( n39022 , n37818 , n37821 );
or ( n39023 , n39021 , n39022 );
xor ( n39024 , n39020 , n39023 );
buf ( n39025 , n39024 );
buf ( n39026 , n39025 );
not ( n39027 , n39026 );
buf ( n39028 , n566 );
not ( n39029 , n39028 );
nor ( n39030 , n39027 , n39029 );
xor ( n39031 , n38217 , n39030 );
xor ( n39032 , n37833 , n38214 );
nor ( n39033 , n37825 , n39029 );
and ( n39034 , n39032 , n39033 );
xor ( n39035 , n39032 , n39033 );
xor ( n39036 , n37837 , n38212 );
nor ( n39037 , n36620 , n39029 );
and ( n39038 , n39036 , n39037 );
xor ( n39039 , n39036 , n39037 );
xor ( n39040 , n37841 , n38210 );
nor ( n39041 , n35419 , n39029 );
and ( n39042 , n39040 , n39041 );
xor ( n39043 , n39040 , n39041 );
xor ( n39044 , n37845 , n38208 );
nor ( n39045 , n34224 , n39029 );
and ( n39046 , n39044 , n39045 );
xor ( n39047 , n39044 , n39045 );
xor ( n39048 , n37849 , n38206 );
nor ( n39049 , n33033 , n39029 );
and ( n39050 , n39048 , n39049 );
xor ( n39051 , n39048 , n39049 );
xor ( n39052 , n37853 , n38204 );
nor ( n39053 , n31867 , n39029 );
and ( n39054 , n39052 , n39053 );
xor ( n39055 , n39052 , n39053 );
xor ( n39056 , n37857 , n38202 );
nor ( n39057 , n30725 , n39029 );
and ( n39058 , n39056 , n39057 );
xor ( n39059 , n39056 , n39057 );
xor ( n39060 , n37861 , n38200 );
nor ( n39061 , n29596 , n39029 );
and ( n39062 , n39060 , n39061 );
xor ( n39063 , n39060 , n39061 );
xor ( n39064 , n37865 , n38198 );
nor ( n39065 , n28487 , n39029 );
and ( n39066 , n39064 , n39065 );
xor ( n39067 , n39064 , n39065 );
xor ( n39068 , n37869 , n38196 );
nor ( n39069 , n27397 , n39029 );
and ( n39070 , n39068 , n39069 );
xor ( n39071 , n39068 , n39069 );
xor ( n39072 , n37873 , n38194 );
nor ( n39073 , n26326 , n39029 );
and ( n39074 , n39072 , n39073 );
xor ( n39075 , n39072 , n39073 );
xor ( n39076 , n37877 , n38192 );
nor ( n39077 , n25272 , n39029 );
and ( n39078 , n39076 , n39077 );
xor ( n39079 , n39076 , n39077 );
xor ( n39080 , n37881 , n38190 );
nor ( n39081 , n24242 , n39029 );
and ( n39082 , n39080 , n39081 );
xor ( n39083 , n39080 , n39081 );
xor ( n39084 , n37885 , n38188 );
nor ( n39085 , n23225 , n39029 );
and ( n39086 , n39084 , n39085 );
xor ( n39087 , n39084 , n39085 );
xor ( n39088 , n37889 , n38186 );
nor ( n39089 , n22231 , n39029 );
and ( n39090 , n39088 , n39089 );
xor ( n39091 , n39088 , n39089 );
xor ( n39092 , n37893 , n38184 );
nor ( n39093 , n21258 , n39029 );
and ( n39094 , n39092 , n39093 );
xor ( n39095 , n39092 , n39093 );
xor ( n39096 , n37897 , n38182 );
nor ( n39097 , n20303 , n39029 );
and ( n39098 , n39096 , n39097 );
xor ( n39099 , n39096 , n39097 );
xor ( n39100 , n37901 , n38180 );
nor ( n39101 , n19365 , n39029 );
and ( n39102 , n39100 , n39101 );
xor ( n39103 , n39100 , n39101 );
xor ( n39104 , n37905 , n38178 );
nor ( n39105 , n18448 , n39029 );
and ( n39106 , n39104 , n39105 );
xor ( n39107 , n39104 , n39105 );
xor ( n39108 , n37909 , n38176 );
nor ( n39109 , n17548 , n39029 );
and ( n39110 , n39108 , n39109 );
xor ( n39111 , n39108 , n39109 );
xor ( n39112 , n37913 , n38174 );
nor ( n39113 , n16669 , n39029 );
and ( n39114 , n39112 , n39113 );
xor ( n39115 , n39112 , n39113 );
xor ( n39116 , n37917 , n38172 );
nor ( n39117 , n15809 , n39029 );
and ( n39118 , n39116 , n39117 );
xor ( n39119 , n39116 , n39117 );
xor ( n39120 , n37921 , n38170 );
nor ( n39121 , n14968 , n39029 );
and ( n39122 , n39120 , n39121 );
xor ( n39123 , n39120 , n39121 );
xor ( n39124 , n37925 , n38168 );
nor ( n39125 , n14147 , n39029 );
and ( n39126 , n39124 , n39125 );
xor ( n39127 , n39124 , n39125 );
xor ( n39128 , n37929 , n38166 );
nor ( n39129 , n13349 , n39029 );
and ( n39130 , n39128 , n39129 );
xor ( n39131 , n39128 , n39129 );
xor ( n39132 , n37933 , n38164 );
nor ( n39133 , n12564 , n39029 );
and ( n39134 , n39132 , n39133 );
xor ( n39135 , n39132 , n39133 );
xor ( n39136 , n37937 , n38162 );
nor ( n39137 , n11799 , n39029 );
and ( n39138 , n39136 , n39137 );
xor ( n39139 , n39136 , n39137 );
xor ( n39140 , n37941 , n38160 );
nor ( n39141 , n11050 , n39029 );
and ( n39142 , n39140 , n39141 );
xor ( n39143 , n39140 , n39141 );
xor ( n39144 , n37945 , n38158 );
nor ( n39145 , n10321 , n39029 );
and ( n39146 , n39144 , n39145 );
xor ( n39147 , n39144 , n39145 );
xor ( n39148 , n37949 , n38156 );
nor ( n39149 , n9429 , n39029 );
and ( n39150 , n39148 , n39149 );
xor ( n39151 , n39148 , n39149 );
xor ( n39152 , n37953 , n38154 );
nor ( n39153 , n8949 , n39029 );
and ( n39154 , n39152 , n39153 );
xor ( n39155 , n39152 , n39153 );
xor ( n39156 , n37957 , n38152 );
nor ( n39157 , n9437 , n39029 );
and ( n39158 , n39156 , n39157 );
xor ( n39159 , n39156 , n39157 );
xor ( n39160 , n37961 , n38150 );
nor ( n39161 , n9446 , n39029 );
and ( n39162 , n39160 , n39161 );
xor ( n39163 , n39160 , n39161 );
xor ( n39164 , n37965 , n38148 );
nor ( n39165 , n9455 , n39029 );
and ( n39166 , n39164 , n39165 );
xor ( n39167 , n39164 , n39165 );
xor ( n39168 , n37969 , n38146 );
nor ( n39169 , n9464 , n39029 );
and ( n39170 , n39168 , n39169 );
xor ( n39171 , n39168 , n39169 );
xor ( n39172 , n37973 , n38144 );
nor ( n39173 , n9473 , n39029 );
and ( n39174 , n39172 , n39173 );
xor ( n39175 , n39172 , n39173 );
xor ( n39176 , n37977 , n38142 );
nor ( n39177 , n9482 , n39029 );
and ( n39178 , n39176 , n39177 );
xor ( n39179 , n39176 , n39177 );
xor ( n39180 , n37981 , n38140 );
nor ( n39181 , n9491 , n39029 );
and ( n39182 , n39180 , n39181 );
xor ( n39183 , n39180 , n39181 );
xor ( n39184 , n37985 , n38138 );
nor ( n39185 , n9500 , n39029 );
and ( n39186 , n39184 , n39185 );
xor ( n39187 , n39184 , n39185 );
xor ( n39188 , n37989 , n38136 );
nor ( n39189 , n9509 , n39029 );
and ( n39190 , n39188 , n39189 );
xor ( n39191 , n39188 , n39189 );
xor ( n39192 , n37993 , n38134 );
nor ( n39193 , n9518 , n39029 );
and ( n39194 , n39192 , n39193 );
xor ( n39195 , n39192 , n39193 );
xor ( n39196 , n37997 , n38132 );
nor ( n39197 , n9527 , n39029 );
and ( n39198 , n39196 , n39197 );
xor ( n39199 , n39196 , n39197 );
xor ( n39200 , n38001 , n38130 );
nor ( n39201 , n9536 , n39029 );
and ( n39202 , n39200 , n39201 );
xor ( n39203 , n39200 , n39201 );
xor ( n39204 , n38005 , n38128 );
nor ( n39205 , n9545 , n39029 );
and ( n39206 , n39204 , n39205 );
xor ( n39207 , n39204 , n39205 );
xor ( n39208 , n38009 , n38126 );
nor ( n39209 , n9554 , n39029 );
and ( n39210 , n39208 , n39209 );
xor ( n39211 , n39208 , n39209 );
xor ( n39212 , n38013 , n38124 );
nor ( n39213 , n9563 , n39029 );
and ( n39214 , n39212 , n39213 );
xor ( n39215 , n39212 , n39213 );
xor ( n39216 , n38017 , n38122 );
nor ( n39217 , n9572 , n39029 );
and ( n39218 , n39216 , n39217 );
xor ( n39219 , n39216 , n39217 );
xor ( n39220 , n38021 , n38120 );
nor ( n39221 , n9581 , n39029 );
and ( n39222 , n39220 , n39221 );
xor ( n39223 , n39220 , n39221 );
xor ( n39224 , n38025 , n38118 );
nor ( n39225 , n9590 , n39029 );
and ( n39226 , n39224 , n39225 );
xor ( n39227 , n39224 , n39225 );
xor ( n39228 , n38029 , n38116 );
nor ( n39229 , n9599 , n39029 );
and ( n39230 , n39228 , n39229 );
xor ( n39231 , n39228 , n39229 );
xor ( n39232 , n38033 , n38114 );
nor ( n39233 , n9608 , n39029 );
and ( n39234 , n39232 , n39233 );
xor ( n39235 , n39232 , n39233 );
xor ( n39236 , n38037 , n38112 );
nor ( n39237 , n9617 , n39029 );
and ( n39238 , n39236 , n39237 );
xor ( n39239 , n39236 , n39237 );
xor ( n39240 , n38041 , n38110 );
nor ( n39241 , n9626 , n39029 );
and ( n39242 , n39240 , n39241 );
xor ( n39243 , n39240 , n39241 );
xor ( n39244 , n38045 , n38108 );
nor ( n39245 , n9635 , n39029 );
and ( n39246 , n39244 , n39245 );
xor ( n39247 , n39244 , n39245 );
xor ( n39248 , n38049 , n38106 );
nor ( n39249 , n9644 , n39029 );
and ( n39250 , n39248 , n39249 );
xor ( n39251 , n39248 , n39249 );
xor ( n39252 , n38053 , n38104 );
nor ( n39253 , n9653 , n39029 );
and ( n39254 , n39252 , n39253 );
xor ( n39255 , n39252 , n39253 );
xor ( n39256 , n38057 , n38102 );
nor ( n39257 , n9662 , n39029 );
and ( n39258 , n39256 , n39257 );
xor ( n39259 , n39256 , n39257 );
xor ( n39260 , n38061 , n38100 );
nor ( n39261 , n9671 , n39029 );
and ( n39262 , n39260 , n39261 );
xor ( n39263 , n39260 , n39261 );
xor ( n39264 , n38065 , n38098 );
nor ( n39265 , n9680 , n39029 );
and ( n39266 , n39264 , n39265 );
xor ( n39267 , n39264 , n39265 );
xor ( n39268 , n38069 , n38096 );
nor ( n39269 , n9689 , n39029 );
and ( n39270 , n39268 , n39269 );
xor ( n39271 , n39268 , n39269 );
xor ( n39272 , n38073 , n38094 );
nor ( n39273 , n9698 , n39029 );
and ( n39274 , n39272 , n39273 );
xor ( n39275 , n39272 , n39273 );
xor ( n39276 , n38077 , n38092 );
nor ( n39277 , n9707 , n39029 );
and ( n39278 , n39276 , n39277 );
xor ( n39279 , n39276 , n39277 );
xor ( n39280 , n38081 , n38090 );
nor ( n39281 , n9716 , n39029 );
and ( n39282 , n39280 , n39281 );
xor ( n39283 , n39280 , n39281 );
xor ( n39284 , n38085 , n38088 );
nor ( n39285 , n9725 , n39029 );
and ( n39286 , n39284 , n39285 );
xor ( n39287 , n39284 , n39285 );
xor ( n39288 , n38086 , n38087 );
nor ( n39289 , n9734 , n39029 );
and ( n39290 , n39288 , n39289 );
xor ( n39291 , n39288 , n39289 );
nor ( n39292 , n9752 , n37827 );
nor ( n39293 , n9743 , n39029 );
and ( n39294 , n39292 , n39293 );
and ( n39295 , n39291 , n39294 );
or ( n39296 , n39290 , n39295 );
and ( n39297 , n39287 , n39296 );
or ( n39298 , n39286 , n39297 );
and ( n39299 , n39283 , n39298 );
or ( n39300 , n39282 , n39299 );
and ( n39301 , n39279 , n39300 );
or ( n39302 , n39278 , n39301 );
and ( n39303 , n39275 , n39302 );
or ( n39304 , n39274 , n39303 );
and ( n39305 , n39271 , n39304 );
or ( n39306 , n39270 , n39305 );
and ( n39307 , n39267 , n39306 );
or ( n39308 , n39266 , n39307 );
and ( n39309 , n39263 , n39308 );
or ( n39310 , n39262 , n39309 );
and ( n39311 , n39259 , n39310 );
or ( n39312 , n39258 , n39311 );
and ( n39313 , n39255 , n39312 );
or ( n39314 , n39254 , n39313 );
and ( n39315 , n39251 , n39314 );
or ( n39316 , n39250 , n39315 );
and ( n39317 , n39247 , n39316 );
or ( n39318 , n39246 , n39317 );
and ( n39319 , n39243 , n39318 );
or ( n39320 , n39242 , n39319 );
and ( n39321 , n39239 , n39320 );
or ( n39322 , n39238 , n39321 );
and ( n39323 , n39235 , n39322 );
or ( n39324 , n39234 , n39323 );
and ( n39325 , n39231 , n39324 );
or ( n39326 , n39230 , n39325 );
and ( n39327 , n39227 , n39326 );
or ( n39328 , n39226 , n39327 );
and ( n39329 , n39223 , n39328 );
or ( n39330 , n39222 , n39329 );
and ( n39331 , n39219 , n39330 );
or ( n39332 , n39218 , n39331 );
and ( n39333 , n39215 , n39332 );
or ( n39334 , n39214 , n39333 );
and ( n39335 , n39211 , n39334 );
or ( n39336 , n39210 , n39335 );
and ( n39337 , n39207 , n39336 );
or ( n39338 , n39206 , n39337 );
and ( n39339 , n39203 , n39338 );
or ( n39340 , n39202 , n39339 );
and ( n39341 , n39199 , n39340 );
or ( n39342 , n39198 , n39341 );
and ( n39343 , n39195 , n39342 );
or ( n39344 , n39194 , n39343 );
and ( n39345 , n39191 , n39344 );
or ( n39346 , n39190 , n39345 );
and ( n39347 , n39187 , n39346 );
or ( n39348 , n39186 , n39347 );
and ( n39349 , n39183 , n39348 );
or ( n39350 , n39182 , n39349 );
and ( n39351 , n39179 , n39350 );
or ( n39352 , n39178 , n39351 );
and ( n39353 , n39175 , n39352 );
or ( n39354 , n39174 , n39353 );
and ( n39355 , n39171 , n39354 );
or ( n39356 , n39170 , n39355 );
and ( n39357 , n39167 , n39356 );
or ( n39358 , n39166 , n39357 );
and ( n39359 , n39163 , n39358 );
or ( n39360 , n39162 , n39359 );
and ( n39361 , n39159 , n39360 );
or ( n39362 , n39158 , n39361 );
and ( n39363 , n39155 , n39362 );
or ( n39364 , n39154 , n39363 );
and ( n39365 , n39151 , n39364 );
or ( n39366 , n39150 , n39365 );
and ( n39367 , n39147 , n39366 );
or ( n39368 , n39146 , n39367 );
and ( n39369 , n39143 , n39368 );
or ( n39370 , n39142 , n39369 );
and ( n39371 , n39139 , n39370 );
or ( n39372 , n39138 , n39371 );
and ( n39373 , n39135 , n39372 );
or ( n39374 , n39134 , n39373 );
and ( n39375 , n39131 , n39374 );
or ( n39376 , n39130 , n39375 );
and ( n39377 , n39127 , n39376 );
or ( n39378 , n39126 , n39377 );
and ( n39379 , n39123 , n39378 );
or ( n39380 , n39122 , n39379 );
and ( n39381 , n39119 , n39380 );
or ( n39382 , n39118 , n39381 );
and ( n39383 , n39115 , n39382 );
or ( n39384 , n39114 , n39383 );
and ( n39385 , n39111 , n39384 );
or ( n39386 , n39110 , n39385 );
and ( n39387 , n39107 , n39386 );
or ( n39388 , n39106 , n39387 );
and ( n39389 , n39103 , n39388 );
or ( n39390 , n39102 , n39389 );
and ( n39391 , n39099 , n39390 );
or ( n39392 , n39098 , n39391 );
and ( n39393 , n39095 , n39392 );
or ( n39394 , n39094 , n39393 );
and ( n39395 , n39091 , n39394 );
or ( n39396 , n39090 , n39395 );
and ( n39397 , n39087 , n39396 );
or ( n39398 , n39086 , n39397 );
and ( n39399 , n39083 , n39398 );
or ( n39400 , n39082 , n39399 );
and ( n39401 , n39079 , n39400 );
or ( n39402 , n39078 , n39401 );
and ( n39403 , n39075 , n39402 );
or ( n39404 , n39074 , n39403 );
and ( n39405 , n39071 , n39404 );
or ( n39406 , n39070 , n39405 );
and ( n39407 , n39067 , n39406 );
or ( n39408 , n39066 , n39407 );
and ( n39409 , n39063 , n39408 );
or ( n39410 , n39062 , n39409 );
and ( n39411 , n39059 , n39410 );
or ( n39412 , n39058 , n39411 );
and ( n39413 , n39055 , n39412 );
or ( n39414 , n39054 , n39413 );
and ( n39415 , n39051 , n39414 );
or ( n39416 , n39050 , n39415 );
and ( n39417 , n39047 , n39416 );
or ( n39418 , n39046 , n39417 );
and ( n39419 , n39043 , n39418 );
or ( n39420 , n39042 , n39419 );
and ( n39421 , n39039 , n39420 );
or ( n39422 , n39038 , n39421 );
and ( n39423 , n39035 , n39422 );
or ( n39424 , n39034 , n39423 );
xor ( n39425 , n39031 , n39424 );
and ( n39426 , n33403 , n732 );
nor ( n39427 , n733 , n39426 );
nor ( n39428 , n796 , n32231 );
xor ( n39429 , n39427 , n39428 );
and ( n39430 , n38219 , n38220 );
and ( n39431 , n38221 , n38224 );
or ( n39432 , n39430 , n39431 );
xor ( n39433 , n39429 , n39432 );
nor ( n39434 , n868 , n31083 );
xor ( n39435 , n39433 , n39434 );
and ( n39436 , n38225 , n38226 );
and ( n39437 , n38227 , n38230 );
or ( n39438 , n39436 , n39437 );
xor ( n39439 , n39435 , n39438 );
nor ( n39440 , n958 , n29948 );
xor ( n39441 , n39439 , n39440 );
and ( n39442 , n38231 , n38232 );
and ( n39443 , n38233 , n38236 );
or ( n39444 , n39442 , n39443 );
xor ( n39445 , n39441 , n39444 );
nor ( n39446 , n1062 , n28833 );
xor ( n39447 , n39445 , n39446 );
and ( n39448 , n38237 , n38238 );
and ( n39449 , n38239 , n38242 );
or ( n39450 , n39448 , n39449 );
xor ( n39451 , n39447 , n39450 );
nor ( n39452 , n1176 , n27737 );
xor ( n39453 , n39451 , n39452 );
and ( n39454 , n38243 , n38244 );
and ( n39455 , n38245 , n38248 );
or ( n39456 , n39454 , n39455 );
xor ( n39457 , n39453 , n39456 );
nor ( n39458 , n1303 , n26660 );
xor ( n39459 , n39457 , n39458 );
and ( n39460 , n38249 , n38250 );
and ( n39461 , n38251 , n38254 );
or ( n39462 , n39460 , n39461 );
xor ( n39463 , n39459 , n39462 );
nor ( n39464 , n1445 , n25600 );
xor ( n39465 , n39463 , n39464 );
and ( n39466 , n38255 , n38256 );
and ( n39467 , n38257 , n38260 );
or ( n39468 , n39466 , n39467 );
xor ( n39469 , n39465 , n39468 );
nor ( n39470 , n1598 , n24564 );
xor ( n39471 , n39469 , n39470 );
and ( n39472 , n38261 , n38262 );
and ( n39473 , n38263 , n38266 );
or ( n39474 , n39472 , n39473 );
xor ( n39475 , n39471 , n39474 );
nor ( n39476 , n1766 , n23541 );
xor ( n39477 , n39475 , n39476 );
and ( n39478 , n38267 , n38268 );
and ( n39479 , n38269 , n38272 );
or ( n39480 , n39478 , n39479 );
xor ( n39481 , n39477 , n39480 );
nor ( n39482 , n1945 , n22541 );
xor ( n39483 , n39481 , n39482 );
and ( n39484 , n38273 , n38274 );
and ( n39485 , n38275 , n38278 );
or ( n39486 , n39484 , n39485 );
xor ( n39487 , n39483 , n39486 );
nor ( n39488 , n2137 , n21562 );
xor ( n39489 , n39487 , n39488 );
and ( n39490 , n38279 , n38280 );
and ( n39491 , n38281 , n38284 );
or ( n39492 , n39490 , n39491 );
xor ( n39493 , n39489 , n39492 );
nor ( n39494 , n2343 , n20601 );
xor ( n39495 , n39493 , n39494 );
and ( n39496 , n38285 , n38286 );
and ( n39497 , n38287 , n38290 );
or ( n39498 , n39496 , n39497 );
xor ( n39499 , n39495 , n39498 );
nor ( n39500 , n2566 , n19657 );
xor ( n39501 , n39499 , n39500 );
and ( n39502 , n38291 , n38292 );
and ( n39503 , n38293 , n38296 );
or ( n39504 , n39502 , n39503 );
xor ( n39505 , n39501 , n39504 );
nor ( n39506 , n2797 , n18734 );
xor ( n39507 , n39505 , n39506 );
and ( n39508 , n38297 , n38298 );
and ( n39509 , n38299 , n38302 );
or ( n39510 , n39508 , n39509 );
xor ( n39511 , n39507 , n39510 );
nor ( n39512 , n3043 , n17828 );
xor ( n39513 , n39511 , n39512 );
and ( n39514 , n38303 , n38304 );
and ( n39515 , n38305 , n38308 );
or ( n39516 , n39514 , n39515 );
xor ( n39517 , n39513 , n39516 );
nor ( n39518 , n3300 , n16943 );
xor ( n39519 , n39517 , n39518 );
and ( n39520 , n38309 , n38310 );
and ( n39521 , n38311 , n38314 );
or ( n39522 , n39520 , n39521 );
xor ( n39523 , n39519 , n39522 );
nor ( n39524 , n3570 , n16077 );
xor ( n39525 , n39523 , n39524 );
and ( n39526 , n38315 , n38316 );
and ( n39527 , n38317 , n38320 );
or ( n39528 , n39526 , n39527 );
xor ( n39529 , n39525 , n39528 );
nor ( n39530 , n3853 , n15230 );
xor ( n39531 , n39529 , n39530 );
and ( n39532 , n38321 , n38322 );
and ( n39533 , n38323 , n38326 );
or ( n39534 , n39532 , n39533 );
xor ( n39535 , n39531 , n39534 );
nor ( n39536 , n4151 , n14403 );
xor ( n39537 , n39535 , n39536 );
and ( n39538 , n38327 , n38328 );
and ( n39539 , n38329 , n38332 );
or ( n39540 , n39538 , n39539 );
xor ( n39541 , n39537 , n39540 );
nor ( n39542 , n4458 , n13599 );
xor ( n39543 , n39541 , n39542 );
and ( n39544 , n38333 , n38334 );
and ( n39545 , n38335 , n38338 );
or ( n39546 , n39544 , n39545 );
xor ( n39547 , n39543 , n39546 );
nor ( n39548 , n4786 , n12808 );
xor ( n39549 , n39547 , n39548 );
and ( n39550 , n38339 , n38340 );
and ( n39551 , n38341 , n38344 );
or ( n39552 , n39550 , n39551 );
xor ( n39553 , n39549 , n39552 );
nor ( n39554 , n5126 , n12037 );
xor ( n39555 , n39553 , n39554 );
and ( n39556 , n38345 , n38346 );
and ( n39557 , n38347 , n38350 );
or ( n39558 , n39556 , n39557 );
xor ( n39559 , n39555 , n39558 );
nor ( n39560 , n5477 , n11282 );
xor ( n39561 , n39559 , n39560 );
and ( n39562 , n38351 , n38352 );
and ( n39563 , n38353 , n38356 );
or ( n39564 , n39562 , n39563 );
xor ( n39565 , n39561 , n39564 );
nor ( n39566 , n5838 , n10547 );
xor ( n39567 , n39565 , n39566 );
and ( n39568 , n38357 , n38358 );
and ( n39569 , n38359 , n38362 );
or ( n39570 , n39568 , n39569 );
xor ( n39571 , n39567 , n39570 );
nor ( n39572 , n6212 , n9829 );
xor ( n39573 , n39571 , n39572 );
and ( n39574 , n38363 , n38364 );
and ( n39575 , n38365 , n38368 );
or ( n39576 , n39574 , n39575 );
xor ( n39577 , n39573 , n39576 );
nor ( n39578 , n6596 , n8955 );
xor ( n39579 , n39577 , n39578 );
and ( n39580 , n38369 , n38370 );
and ( n39581 , n38371 , n38374 );
or ( n39582 , n39580 , n39581 );
xor ( n39583 , n39579 , n39582 );
nor ( n39584 , n6997 , n603 );
xor ( n39585 , n39583 , n39584 );
and ( n39586 , n38375 , n38376 );
and ( n39587 , n38377 , n38380 );
or ( n39588 , n39586 , n39587 );
xor ( n39589 , n39585 , n39588 );
nor ( n39590 , n7413 , n652 );
xor ( n39591 , n39589 , n39590 );
and ( n39592 , n38381 , n38382 );
and ( n39593 , n38383 , n38386 );
or ( n39594 , n39592 , n39593 );
xor ( n39595 , n39591 , n39594 );
nor ( n39596 , n7841 , n624 );
xor ( n39597 , n39595 , n39596 );
and ( n39598 , n38387 , n38388 );
and ( n39599 , n38389 , n38392 );
or ( n39600 , n39598 , n39599 );
xor ( n39601 , n39597 , n39600 );
nor ( n39602 , n8281 , n648 );
xor ( n39603 , n39601 , n39602 );
and ( n39604 , n38393 , n38394 );
and ( n39605 , n38395 , n38398 );
or ( n39606 , n39604 , n39605 );
xor ( n39607 , n39603 , n39606 );
nor ( n39608 , n8737 , n686 );
xor ( n39609 , n39607 , n39608 );
and ( n39610 , n38399 , n38400 );
and ( n39611 , n38401 , n38404 );
or ( n39612 , n39610 , n39611 );
xor ( n39613 , n39609 , n39612 );
nor ( n39614 , n9420 , n735 );
xor ( n39615 , n39613 , n39614 );
and ( n39616 , n38405 , n38406 );
and ( n39617 , n38407 , n38410 );
or ( n39618 , n39616 , n39617 );
xor ( n39619 , n39615 , n39618 );
nor ( n39620 , n10312 , n798 );
xor ( n39621 , n39619 , n39620 );
and ( n39622 , n38411 , n38412 );
and ( n39623 , n38413 , n38416 );
or ( n39624 , n39622 , n39623 );
xor ( n39625 , n39621 , n39624 );
nor ( n39626 , n11041 , n870 );
xor ( n39627 , n39625 , n39626 );
and ( n39628 , n38417 , n38418 );
and ( n39629 , n38419 , n38422 );
or ( n39630 , n39628 , n39629 );
xor ( n39631 , n39627 , n39630 );
nor ( n39632 , n11790 , n960 );
xor ( n39633 , n39631 , n39632 );
and ( n39634 , n38423 , n38424 );
and ( n39635 , n38425 , n38428 );
or ( n39636 , n39634 , n39635 );
xor ( n39637 , n39633 , n39636 );
nor ( n39638 , n12555 , n1064 );
xor ( n39639 , n39637 , n39638 );
and ( n39640 , n38429 , n38430 );
and ( n39641 , n38431 , n38434 );
or ( n39642 , n39640 , n39641 );
xor ( n39643 , n39639 , n39642 );
nor ( n39644 , n13340 , n1178 );
xor ( n39645 , n39643 , n39644 );
and ( n39646 , n38435 , n38436 );
and ( n39647 , n38437 , n38440 );
or ( n39648 , n39646 , n39647 );
xor ( n39649 , n39645 , n39648 );
nor ( n39650 , n14138 , n1305 );
xor ( n39651 , n39649 , n39650 );
and ( n39652 , n38441 , n38442 );
and ( n39653 , n38443 , n38446 );
or ( n39654 , n39652 , n39653 );
xor ( n39655 , n39651 , n39654 );
nor ( n39656 , n14959 , n1447 );
xor ( n39657 , n39655 , n39656 );
and ( n39658 , n38447 , n38448 );
and ( n39659 , n38449 , n38452 );
or ( n39660 , n39658 , n39659 );
xor ( n39661 , n39657 , n39660 );
nor ( n39662 , n15800 , n1600 );
xor ( n39663 , n39661 , n39662 );
and ( n39664 , n38453 , n38454 );
and ( n39665 , n38455 , n38458 );
or ( n39666 , n39664 , n39665 );
xor ( n39667 , n39663 , n39666 );
nor ( n39668 , n16660 , n1768 );
xor ( n39669 , n39667 , n39668 );
and ( n39670 , n38459 , n38460 );
and ( n39671 , n38461 , n38464 );
or ( n39672 , n39670 , n39671 );
xor ( n39673 , n39669 , n39672 );
nor ( n39674 , n17539 , n1947 );
xor ( n39675 , n39673 , n39674 );
and ( n39676 , n38465 , n38466 );
and ( n39677 , n38467 , n38470 );
or ( n39678 , n39676 , n39677 );
xor ( n39679 , n39675 , n39678 );
nor ( n39680 , n18439 , n2139 );
xor ( n39681 , n39679 , n39680 );
and ( n39682 , n38471 , n38472 );
and ( n39683 , n38473 , n38476 );
or ( n39684 , n39682 , n39683 );
xor ( n39685 , n39681 , n39684 );
nor ( n39686 , n19356 , n2345 );
xor ( n39687 , n39685 , n39686 );
and ( n39688 , n38477 , n38478 );
and ( n39689 , n38479 , n38482 );
or ( n39690 , n39688 , n39689 );
xor ( n39691 , n39687 , n39690 );
nor ( n39692 , n20294 , n2568 );
xor ( n39693 , n39691 , n39692 );
and ( n39694 , n38483 , n38484 );
and ( n39695 , n38485 , n38488 );
or ( n39696 , n39694 , n39695 );
xor ( n39697 , n39693 , n39696 );
nor ( n39698 , n21249 , n2799 );
xor ( n39699 , n39697 , n39698 );
and ( n39700 , n38489 , n38490 );
and ( n39701 , n38491 , n38494 );
or ( n39702 , n39700 , n39701 );
xor ( n39703 , n39699 , n39702 );
nor ( n39704 , n22222 , n3045 );
xor ( n39705 , n39703 , n39704 );
and ( n39706 , n38495 , n38496 );
and ( n39707 , n38497 , n38500 );
or ( n39708 , n39706 , n39707 );
xor ( n39709 , n39705 , n39708 );
nor ( n39710 , n23216 , n3302 );
xor ( n39711 , n39709 , n39710 );
and ( n39712 , n38501 , n38502 );
and ( n39713 , n38503 , n38506 );
or ( n39714 , n39712 , n39713 );
xor ( n39715 , n39711 , n39714 );
nor ( n39716 , n24233 , n3572 );
xor ( n39717 , n39715 , n39716 );
and ( n39718 , n38507 , n38508 );
and ( n39719 , n38509 , n38512 );
or ( n39720 , n39718 , n39719 );
xor ( n39721 , n39717 , n39720 );
nor ( n39722 , n25263 , n3855 );
xor ( n39723 , n39721 , n39722 );
and ( n39724 , n38513 , n38514 );
and ( n39725 , n38515 , n38518 );
or ( n39726 , n39724 , n39725 );
xor ( n39727 , n39723 , n39726 );
nor ( n39728 , n26317 , n4153 );
xor ( n39729 , n39727 , n39728 );
and ( n39730 , n38519 , n38520 );
and ( n39731 , n38521 , n38524 );
or ( n39732 , n39730 , n39731 );
xor ( n39733 , n39729 , n39732 );
nor ( n39734 , n27388 , n4460 );
xor ( n39735 , n39733 , n39734 );
and ( n39736 , n38525 , n38526 );
and ( n39737 , n38527 , n38530 );
or ( n39738 , n39736 , n39737 );
xor ( n39739 , n39735 , n39738 );
nor ( n39740 , n28478 , n4788 );
xor ( n39741 , n39739 , n39740 );
and ( n39742 , n38531 , n38532 );
and ( n39743 , n38533 , n38536 );
or ( n39744 , n39742 , n39743 );
xor ( n39745 , n39741 , n39744 );
nor ( n39746 , n29587 , n5128 );
xor ( n39747 , n39745 , n39746 );
and ( n39748 , n38537 , n38538 );
and ( n39749 , n38539 , n38542 );
or ( n39750 , n39748 , n39749 );
xor ( n39751 , n39747 , n39750 );
nor ( n39752 , n30716 , n5479 );
xor ( n39753 , n39751 , n39752 );
and ( n39754 , n38543 , n38544 );
and ( n39755 , n38545 , n38548 );
or ( n39756 , n39754 , n39755 );
xor ( n39757 , n39753 , n39756 );
nor ( n39758 , n31858 , n5840 );
xor ( n39759 , n39757 , n39758 );
and ( n39760 , n38549 , n38550 );
and ( n39761 , n38551 , n38554 );
or ( n39762 , n39760 , n39761 );
xor ( n39763 , n39759 , n39762 );
nor ( n39764 , n33024 , n6214 );
xor ( n39765 , n39763 , n39764 );
and ( n39766 , n38555 , n38556 );
and ( n39767 , n38557 , n38560 );
or ( n39768 , n39766 , n39767 );
xor ( n39769 , n39765 , n39768 );
nor ( n39770 , n34215 , n6598 );
xor ( n39771 , n39769 , n39770 );
and ( n39772 , n38561 , n38562 );
and ( n39773 , n38563 , n38566 );
or ( n39774 , n39772 , n39773 );
xor ( n39775 , n39771 , n39774 );
nor ( n39776 , n35410 , n6999 );
xor ( n39777 , n39775 , n39776 );
and ( n39778 , n38567 , n38568 );
and ( n39779 , n38569 , n38572 );
or ( n39780 , n39778 , n39779 );
xor ( n39781 , n39777 , n39780 );
nor ( n39782 , n36611 , n7415 );
xor ( n39783 , n39781 , n39782 );
and ( n39784 , n38573 , n38574 );
and ( n39785 , n38575 , n38578 );
or ( n39786 , n39784 , n39785 );
xor ( n39787 , n39783 , n39786 );
nor ( n39788 , n37816 , n7843 );
xor ( n39789 , n39787 , n39788 );
and ( n39790 , n38579 , n38580 );
and ( n39791 , n38581 , n38584 );
or ( n39792 , n39790 , n39791 );
xor ( n39793 , n39789 , n39792 );
nor ( n39794 , n39018 , n8283 );
xor ( n39795 , n39793 , n39794 );
and ( n39796 , n38585 , n38586 );
and ( n39797 , n38587 , n38590 );
or ( n39798 , n39796 , n39797 );
xor ( n39799 , n39795 , n39798 );
and ( n39800 , n38603 , n38607 );
and ( n39801 , n38607 , n39004 );
and ( n39802 , n38603 , n39004 );
or ( n39803 , n39800 , n39801 , n39802 );
and ( n39804 , n33774 , n719 );
not ( n39805 , n719 );
nor ( n39806 , n39804 , n39805 );
xor ( n39807 , n39803 , n39806 );
and ( n39808 , n38616 , n38620 );
and ( n39809 , n38620 , n38688 );
and ( n39810 , n38616 , n38688 );
or ( n39811 , n39808 , n39809 , n39810 );
and ( n39812 , n38612 , n38689 );
and ( n39813 , n38689 , n39003 );
and ( n39814 , n38612 , n39003 );
or ( n39815 , n39812 , n39813 , n39814 );
xor ( n39816 , n39811 , n39815 );
and ( n39817 , n38694 , n38814 );
and ( n39818 , n38814 , n39002 );
and ( n39819 , n38694 , n39002 );
or ( n39820 , n39817 , n39818 , n39819 );
and ( n39821 , n38625 , n38629 );
and ( n39822 , n38629 , n38687 );
and ( n39823 , n38625 , n38687 );
or ( n39824 , n39821 , n39822 , n39823 );
and ( n39825 , n38698 , n38702 );
and ( n39826 , n38702 , n38813 );
and ( n39827 , n38698 , n38813 );
or ( n39828 , n39825 , n39826 , n39827 );
xor ( n39829 , n39824 , n39828 );
and ( n39830 , n38656 , n38660 );
and ( n39831 , n38660 , n38666 );
and ( n39832 , n38656 , n38666 );
or ( n39833 , n39830 , n39831 , n39832 );
and ( n39834 , n38634 , n38638 );
and ( n39835 , n38638 , n38686 );
and ( n39836 , n38634 , n38686 );
or ( n39837 , n39834 , n39835 , n39836 );
xor ( n39838 , n39833 , n39837 );
and ( n39839 , n38711 , n38736 );
and ( n39840 , n38736 , n38774 );
and ( n39841 , n38711 , n38774 );
or ( n39842 , n39839 , n39840 , n39841 );
and ( n39843 , n38643 , n38647 );
and ( n39844 , n38647 , n38685 );
and ( n39845 , n38643 , n38685 );
or ( n39846 , n39843 , n39844 , n39845 );
xor ( n39847 , n39842 , n39846 );
and ( n39848 , n38652 , n38667 );
and ( n39849 , n38667 , n38684 );
and ( n39850 , n38652 , n38684 );
or ( n39851 , n39848 , n39849 , n39850 );
and ( n39852 , n38715 , n38719 );
and ( n39853 , n38719 , n38735 );
and ( n39854 , n38715 , n38735 );
or ( n39855 , n39852 , n39853 , n39854 );
xor ( n39856 , n39851 , n39855 );
and ( n39857 , n38672 , n38677 );
and ( n39858 , n38677 , n38683 );
and ( n39859 , n38672 , n38683 );
or ( n39860 , n39857 , n39858 , n39859 );
and ( n39861 , n38662 , n38663 );
and ( n39862 , n38663 , n38665 );
and ( n39863 , n38662 , n38665 );
or ( n39864 , n39861 , n39862 , n39863 );
and ( n39865 , n38673 , n38674 );
and ( n39866 , n38674 , n38676 );
and ( n39867 , n38673 , n38676 );
or ( n39868 , n39865 , n39866 , n39867 );
xor ( n39869 , n39864 , n39868 );
and ( n39870 , n30695 , n940 );
and ( n39871 , n31836 , n840 );
xor ( n39872 , n39870 , n39871 );
and ( n39873 , n32649 , n771 );
xor ( n39874 , n39872 , n39873 );
xor ( n39875 , n39869 , n39874 );
xor ( n39876 , n39860 , n39875 );
and ( n39877 , n38679 , n38680 );
and ( n39878 , n38680 , n38682 );
and ( n39879 , n38679 , n38682 );
or ( n39880 , n39877 , n39878 , n39879 );
and ( n39881 , n27361 , n1254 );
and ( n39882 , n28456 , n1134 );
xor ( n39883 , n39881 , n39882 );
and ( n39884 , n29559 , n1034 );
xor ( n39885 , n39883 , n39884 );
xor ( n39886 , n39880 , n39885 );
and ( n39887 , n24214 , n1738 );
and ( n39888 , n25243 , n1551 );
xor ( n39889 , n39887 , n39888 );
and ( n39890 , n26296 , n1424 );
xor ( n39891 , n39889 , n39890 );
xor ( n39892 , n39886 , n39891 );
xor ( n39893 , n39876 , n39892 );
xor ( n39894 , n39856 , n39893 );
xor ( n39895 , n39847 , n39894 );
xor ( n39896 , n39838 , n39895 );
xor ( n39897 , n39829 , n39896 );
xor ( n39898 , n39820 , n39897 );
and ( n39899 , n38819 , n38894 );
and ( n39900 , n38894 , n39001 );
and ( n39901 , n38819 , n39001 );
or ( n39902 , n39899 , n39900 , n39901 );
and ( n39903 , n38707 , n38775 );
and ( n39904 , n38775 , n38812 );
and ( n39905 , n38707 , n38812 );
or ( n39906 , n39903 , n39904 , n39905 );
and ( n39907 , n38823 , n38827 );
and ( n39908 , n38827 , n38893 );
and ( n39909 , n38823 , n38893 );
or ( n39910 , n39907 , n39908 , n39909 );
xor ( n39911 , n39906 , n39910 );
and ( n39912 , n38780 , n38784 );
and ( n39913 , n38784 , n38811 );
and ( n39914 , n38780 , n38811 );
or ( n39915 , n39912 , n39913 , n39914 );
and ( n39916 , n38741 , n38757 );
and ( n39917 , n38757 , n38773 );
and ( n39918 , n38741 , n38773 );
or ( n39919 , n39916 , n39917 , n39918 );
and ( n39920 , n38724 , n38728 );
and ( n39921 , n38728 , n38734 );
and ( n39922 , n38724 , n38734 );
or ( n39923 , n39920 , n39921 , n39922 );
and ( n39924 , n38745 , n38750 );
and ( n39925 , n38750 , n38756 );
and ( n39926 , n38745 , n38756 );
or ( n39927 , n39924 , n39925 , n39926 );
xor ( n39928 , n39923 , n39927 );
and ( n39929 , n38730 , n38731 );
and ( n39930 , n38731 , n38733 );
and ( n39931 , n38730 , n38733 );
or ( n39932 , n39929 , n39930 , n39931 );
and ( n39933 , n38746 , n38747 );
and ( n39934 , n38747 , n38749 );
and ( n39935 , n38746 , n38749 );
or ( n39936 , n39933 , n39934 , n39935 );
xor ( n39937 , n39932 , n39936 );
and ( n39938 , n21216 , n2298 );
and ( n39939 , n22186 , n2100 );
xor ( n39940 , n39938 , n39939 );
and ( n39941 , n22892 , n1882 );
xor ( n39942 , n39940 , n39941 );
xor ( n39943 , n39937 , n39942 );
xor ( n39944 , n39928 , n39943 );
xor ( n39945 , n39919 , n39944 );
and ( n39946 , n38762 , n38766 );
and ( n39947 , n38766 , n38772 );
and ( n39948 , n38762 , n38772 );
or ( n39949 , n39946 , n39947 , n39948 );
and ( n39950 , n38752 , n38753 );
and ( n39951 , n38753 , n38755 );
and ( n39952 , n38752 , n38755 );
or ( n39953 , n39950 , n39951 , n39952 );
and ( n39954 , n18144 , n2981 );
and ( n39955 , n19324 , n2739 );
xor ( n39956 , n39954 , n39955 );
and ( n39957 , n20233 , n2544 );
xor ( n39958 , n39956 , n39957 );
xor ( n39959 , n39953 , n39958 );
and ( n39960 , n15758 , n3749 );
and ( n39961 , n16637 , n3495 );
xor ( n39962 , n39960 , n39961 );
and ( n39963 , n17512 , n3271 );
xor ( n39964 , n39962 , n39963 );
xor ( n39965 , n39959 , n39964 );
xor ( n39966 , n39949 , n39965 );
and ( n39967 , n38768 , n38769 );
and ( n39968 , n38769 , n38771 );
and ( n39969 , n38768 , n38771 );
or ( n39970 , n39967 , n39968 , n39969 );
and ( n39971 , n38799 , n38800 );
and ( n39972 , n38800 , n38802 );
and ( n39973 , n38799 , n38802 );
or ( n39974 , n39971 , n39972 , n39973 );
xor ( n39975 , n39970 , n39974 );
and ( n39976 , n13322 , n4730 );
and ( n39977 , n14118 , n4403 );
xor ( n39978 , n39976 , n39977 );
and ( n39979 , n14938 , n4102 );
xor ( n39980 , n39978 , n39979 );
xor ( n39981 , n39975 , n39980 );
xor ( n39982 , n39966 , n39981 );
xor ( n39983 , n39945 , n39982 );
xor ( n39984 , n39915 , n39983 );
and ( n39985 , n38789 , n38793 );
and ( n39986 , n38793 , n38810 );
and ( n39987 , n38789 , n38810 );
or ( n39988 , n39985 , n39986 , n39987 );
and ( n39989 , n38836 , n38848 );
and ( n39990 , n38848 , n38865 );
and ( n39991 , n38836 , n38865 );
or ( n39992 , n39989 , n39990 , n39991 );
xor ( n39993 , n39988 , n39992 );
and ( n39994 , n38798 , n38803 );
and ( n39995 , n38803 , n38809 );
and ( n39996 , n38798 , n38809 );
or ( n39997 , n39994 , n39995 , n39996 );
and ( n39998 , n38840 , n38844 );
and ( n39999 , n38844 , n38847 );
and ( n40000 , n38840 , n38847 );
or ( n40001 , n39998 , n39999 , n40000 );
xor ( n40002 , n39997 , n40001 );
and ( n40003 , n38805 , n38806 );
and ( n40004 , n38806 , n38808 );
and ( n40005 , n38805 , n38808 );
or ( n40006 , n40003 , n40004 , n40005 );
and ( n40007 , n11015 , n5765 );
and ( n40008 , n11769 , n5408 );
xor ( n40009 , n40007 , n40008 );
and ( n40010 , n12320 , n5103 );
xor ( n40011 , n40009 , n40010 );
xor ( n40012 , n40006 , n40011 );
and ( n40013 , n8718 , n6971 );
and ( n40014 , n9400 , n6504 );
xor ( n40015 , n40013 , n40014 );
and ( n40016 , n10291 , n6132 );
xor ( n40017 , n40015 , n40016 );
xor ( n40018 , n40012 , n40017 );
xor ( n40019 , n40002 , n40018 );
xor ( n40020 , n39993 , n40019 );
xor ( n40021 , n39984 , n40020 );
xor ( n40022 , n39911 , n40021 );
xor ( n40023 , n39902 , n40022 );
and ( n40024 , n38899 , n38946 );
and ( n40025 , n38946 , n39000 );
and ( n40026 , n38899 , n39000 );
or ( n40027 , n40024 , n40025 , n40026 );
and ( n40028 , n38832 , n38866 );
and ( n40029 , n38866 , n38892 );
and ( n40030 , n38832 , n38892 );
or ( n40031 , n40028 , n40029 , n40030 );
and ( n40032 , n38903 , n38907 );
and ( n40033 , n38907 , n38945 );
and ( n40034 , n38903 , n38945 );
or ( n40035 , n40032 , n40033 , n40034 );
xor ( n40036 , n40031 , n40035 );
and ( n40037 , n38871 , n38875 );
and ( n40038 , n38875 , n38891 );
and ( n40039 , n38871 , n38891 );
or ( n40040 , n40037 , n40038 , n40039 );
and ( n40041 , n38853 , n38858 );
and ( n40042 , n38858 , n38864 );
and ( n40043 , n38853 , n38864 );
or ( n40044 , n40041 , n40042 , n40043 );
and ( n40045 , n7385 , n7662 );
and ( n40046 , n7808 , n7310 );
and ( n40047 , n40045 , n40046 );
and ( n40048 , n40046 , n38846 );
and ( n40049 , n40045 , n38846 );
or ( n40050 , n40047 , n40048 , n40049 );
and ( n40051 , n38854 , n38855 );
and ( n40052 , n38855 , n38857 );
and ( n40053 , n38854 , n38857 );
or ( n40054 , n40051 , n40052 , n40053 );
xor ( n40055 , n40050 , n40054 );
and ( n40056 , n7385 , n8243 );
buf ( n40057 , n7808 );
xor ( n40058 , n40056 , n40057 );
and ( n40059 , n8079 , n7310 );
xor ( n40060 , n40058 , n40059 );
xor ( n40061 , n40055 , n40060 );
xor ( n40062 , n40044 , n40061 );
and ( n40063 , n38860 , n38861 );
and ( n40064 , n38861 , n38863 );
and ( n40065 , n38860 , n38863 );
or ( n40066 , n40063 , n40064 , n40065 );
and ( n40067 , n6187 , n10239 );
and ( n40068 , n6569 , n9348 );
xor ( n40069 , n40067 , n40068 );
and ( n40070 , n6816 , n8669 );
xor ( n40071 , n40069 , n40070 );
xor ( n40072 , n40066 , n40071 );
and ( n40073 , n4959 , n12531 );
and ( n40074 , n5459 , n11718 );
xor ( n40075 , n40073 , n40074 );
and ( n40076 , n5819 , n10977 );
xor ( n40077 , n40075 , n40076 );
xor ( n40078 , n40072 , n40077 );
xor ( n40079 , n40062 , n40078 );
xor ( n40080 , n40040 , n40079 );
and ( n40081 , n38880 , n38884 );
and ( n40082 , n38884 , n38890 );
and ( n40083 , n38880 , n38890 );
or ( n40084 , n40081 , n40082 , n40083 );
and ( n40085 , n38916 , n38921 );
and ( n40086 , n38921 , n38927 );
and ( n40087 , n38916 , n38927 );
or ( n40088 , n40085 , n40086 , n40087 );
xor ( n40089 , n40084 , n40088 );
and ( n40090 , n38886 , n38887 );
and ( n40091 , n38887 , n38889 );
and ( n40092 , n38886 , n38889 );
or ( n40093 , n40090 , n40091 , n40092 );
and ( n40094 , n38917 , n38918 );
and ( n40095 , n38918 , n38920 );
and ( n40096 , n38917 , n38920 );
or ( n40097 , n40094 , n40095 , n40096 );
xor ( n40098 , n40093 , n40097 );
and ( n40099 , n4132 , n14838 );
and ( n40100 , n4438 , n14044 );
xor ( n40101 , n40099 , n40100 );
and ( n40102 , n4766 , n13256 );
xor ( n40103 , n40101 , n40102 );
xor ( n40104 , n40098 , n40103 );
xor ( n40105 , n40089 , n40104 );
xor ( n40106 , n40080 , n40105 );
xor ( n40107 , n40036 , n40106 );
xor ( n40108 , n40027 , n40107 );
and ( n40109 , n38951 , n38977 );
and ( n40110 , n38977 , n38999 );
and ( n40111 , n38951 , n38999 );
or ( n40112 , n40109 , n40110 , n40111 );
and ( n40113 , n38912 , n38928 );
and ( n40114 , n38928 , n38944 );
and ( n40115 , n38912 , n38944 );
or ( n40116 , n40113 , n40114 , n40115 );
and ( n40117 , n38955 , n38959 );
and ( n40118 , n38959 , n38976 );
and ( n40119 , n38955 , n38976 );
or ( n40120 , n40117 , n40118 , n40119 );
xor ( n40121 , n40116 , n40120 );
and ( n40122 , n38933 , n38937 );
and ( n40123 , n38937 , n38943 );
and ( n40124 , n38933 , n38943 );
or ( n40125 , n40122 , n40123 , n40124 );
and ( n40126 , n38923 , n38924 );
and ( n40127 , n38924 , n38926 );
and ( n40128 , n38923 , n38926 );
or ( n40129 , n40126 , n40127 , n40128 );
and ( n40130 , n3182 , n17422 );
and ( n40131 , n3545 , n16550 );
xor ( n40132 , n40130 , n40131 );
and ( n40133 , n3801 , n15691 );
xor ( n40134 , n40132 , n40133 );
xor ( n40135 , n40129 , n40134 );
and ( n40136 , n2462 , n20156 );
and ( n40137 , n2779 , n19222 );
xor ( n40138 , n40136 , n40137 );
and ( n40139 , n3024 , n18407 );
xor ( n40140 , n40138 , n40139 );
xor ( n40141 , n40135 , n40140 );
xor ( n40142 , n40125 , n40141 );
and ( n40143 , n38939 , n38940 );
and ( n40144 , n38940 , n38942 );
and ( n40145 , n38939 , n38942 );
or ( n40146 , n40143 , n40144 , n40145 );
and ( n40147 , n38965 , n38966 );
and ( n40148 , n38966 , n38968 );
and ( n40149 , n38965 , n38968 );
or ( n40150 , n40147 , n40148 , n40149 );
xor ( n40151 , n40146 , n40150 );
and ( n40152 , n1933 , n23075 );
and ( n40153 , n2120 , n22065 );
xor ( n40154 , n40152 , n40153 );
and ( n40155 , n2324 , n20976 );
xor ( n40156 , n40154 , n40155 );
xor ( n40157 , n40151 , n40156 );
xor ( n40158 , n40142 , n40157 );
xor ( n40159 , n40121 , n40158 );
xor ( n40160 , n40112 , n40159 );
and ( n40161 , n38993 , n38998 );
and ( n40162 , n38982 , n38986 );
and ( n40163 , n38986 , n38992 );
and ( n40164 , n38982 , n38992 );
or ( n40165 , n40162 , n40163 , n40164 );
and ( n40166 , n38964 , n38969 );
and ( n40167 , n38969 , n38975 );
and ( n40168 , n38964 , n38975 );
or ( n40169 , n40166 , n40167 , n40168 );
xor ( n40170 , n40165 , n40169 );
and ( n40171 , n38971 , n38972 );
and ( n40172 , n38972 , n38974 );
and ( n40173 , n38971 , n38974 );
or ( n40174 , n40171 , n40172 , n40173 );
and ( n40175 , n1383 , n26216 );
and ( n40176 , n1580 , n25163 );
xor ( n40177 , n40175 , n40176 );
and ( n40178 , n1694 , n24137 );
xor ( n40179 , n40177 , n40178 );
xor ( n40180 , n40174 , n40179 );
and ( n40181 , n1047 , n29508 );
and ( n40182 , n1164 , n28406 );
xor ( n40183 , n40181 , n40182 );
and ( n40184 , n1287 , n27296 );
xor ( n40185 , n40183 , n40184 );
xor ( n40186 , n40180 , n40185 );
xor ( n40187 , n40170 , n40186 );
xor ( n40188 , n40161 , n40187 );
not ( n40189 , n715 );
and ( n40190 , n34193 , n715 );
nor ( n40191 , n40189 , n40190 );
and ( n40192 , n38988 , n38989 );
and ( n40193 , n38989 , n38991 );
and ( n40194 , n38988 , n38991 );
or ( n40195 , n40192 , n40193 , n40194 );
and ( n40196 , n38996 , n38997 );
xor ( n40197 , n40195 , n40196 );
and ( n40198 , n783 , n32999 );
and ( n40199 , n856 , n31761 );
xor ( n40200 , n40198 , n40199 );
and ( n40201 , n925 , n30629 );
xor ( n40202 , n40200 , n40201 );
xor ( n40203 , n40197 , n40202 );
xor ( n40204 , n40191 , n40203 );
xor ( n40205 , n40188 , n40204 );
xor ( n40206 , n40160 , n40205 );
xor ( n40207 , n40108 , n40206 );
xor ( n40208 , n40023 , n40207 );
xor ( n40209 , n39898 , n40208 );
xor ( n40210 , n39816 , n40209 );
xor ( n40211 , n39807 , n40210 );
and ( n40212 , n38595 , n38598 );
and ( n40213 , n38598 , n39005 );
and ( n40214 , n38595 , n39005 );
or ( n40215 , n40212 , n40213 , n40214 );
xor ( n40216 , n40211 , n40215 );
and ( n40217 , n39006 , n39010 );
and ( n40218 , n39011 , n39014 );
or ( n40219 , n40217 , n40218 );
xor ( n40220 , n40216 , n40219 );
buf ( n40221 , n40220 );
buf ( n40222 , n40221 );
not ( n40223 , n40222 );
nor ( n40224 , n40223 , n8739 );
xor ( n40225 , n39799 , n40224 );
and ( n40226 , n38591 , n39019 );
and ( n40227 , n39020 , n39023 );
or ( n40228 , n40226 , n40227 );
xor ( n40229 , n40225 , n40228 );
buf ( n40230 , n40229 );
buf ( n40231 , n40230 );
not ( n40232 , n40231 );
buf ( n40233 , n567 );
not ( n40234 , n40233 );
nor ( n40235 , n40232 , n40234 );
xor ( n40236 , n39425 , n40235 );
xor ( n40237 , n39035 , n39422 );
nor ( n40238 , n39027 , n40234 );
and ( n40239 , n40237 , n40238 );
xor ( n40240 , n40237 , n40238 );
xor ( n40241 , n39039 , n39420 );
nor ( n40242 , n37825 , n40234 );
and ( n40243 , n40241 , n40242 );
xor ( n40244 , n40241 , n40242 );
xor ( n40245 , n39043 , n39418 );
nor ( n40246 , n36620 , n40234 );
and ( n40247 , n40245 , n40246 );
xor ( n40248 , n40245 , n40246 );
xor ( n40249 , n39047 , n39416 );
nor ( n40250 , n35419 , n40234 );
and ( n40251 , n40249 , n40250 );
xor ( n40252 , n40249 , n40250 );
xor ( n40253 , n39051 , n39414 );
nor ( n40254 , n34224 , n40234 );
and ( n40255 , n40253 , n40254 );
xor ( n40256 , n40253 , n40254 );
xor ( n40257 , n39055 , n39412 );
nor ( n40258 , n33033 , n40234 );
and ( n40259 , n40257 , n40258 );
xor ( n40260 , n40257 , n40258 );
xor ( n40261 , n39059 , n39410 );
nor ( n40262 , n31867 , n40234 );
and ( n40263 , n40261 , n40262 );
xor ( n40264 , n40261 , n40262 );
xor ( n40265 , n39063 , n39408 );
nor ( n40266 , n30725 , n40234 );
and ( n40267 , n40265 , n40266 );
xor ( n40268 , n40265 , n40266 );
xor ( n40269 , n39067 , n39406 );
nor ( n40270 , n29596 , n40234 );
and ( n40271 , n40269 , n40270 );
xor ( n40272 , n40269 , n40270 );
xor ( n40273 , n39071 , n39404 );
nor ( n40274 , n28487 , n40234 );
and ( n40275 , n40273 , n40274 );
xor ( n40276 , n40273 , n40274 );
xor ( n40277 , n39075 , n39402 );
nor ( n40278 , n27397 , n40234 );
and ( n40279 , n40277 , n40278 );
xor ( n40280 , n40277 , n40278 );
xor ( n40281 , n39079 , n39400 );
nor ( n40282 , n26326 , n40234 );
and ( n40283 , n40281 , n40282 );
xor ( n40284 , n40281 , n40282 );
xor ( n40285 , n39083 , n39398 );
nor ( n40286 , n25272 , n40234 );
and ( n40287 , n40285 , n40286 );
xor ( n40288 , n40285 , n40286 );
xor ( n40289 , n39087 , n39396 );
nor ( n40290 , n24242 , n40234 );
and ( n40291 , n40289 , n40290 );
xor ( n40292 , n40289 , n40290 );
xor ( n40293 , n39091 , n39394 );
nor ( n40294 , n23225 , n40234 );
and ( n40295 , n40293 , n40294 );
xor ( n40296 , n40293 , n40294 );
xor ( n40297 , n39095 , n39392 );
nor ( n40298 , n22231 , n40234 );
and ( n40299 , n40297 , n40298 );
xor ( n40300 , n40297 , n40298 );
xor ( n40301 , n39099 , n39390 );
nor ( n40302 , n21258 , n40234 );
and ( n40303 , n40301 , n40302 );
xor ( n40304 , n40301 , n40302 );
xor ( n40305 , n39103 , n39388 );
nor ( n40306 , n20303 , n40234 );
and ( n40307 , n40305 , n40306 );
xor ( n40308 , n40305 , n40306 );
xor ( n40309 , n39107 , n39386 );
nor ( n40310 , n19365 , n40234 );
and ( n40311 , n40309 , n40310 );
xor ( n40312 , n40309 , n40310 );
xor ( n40313 , n39111 , n39384 );
nor ( n40314 , n18448 , n40234 );
and ( n40315 , n40313 , n40314 );
xor ( n40316 , n40313 , n40314 );
xor ( n40317 , n39115 , n39382 );
nor ( n40318 , n17548 , n40234 );
and ( n40319 , n40317 , n40318 );
xor ( n40320 , n40317 , n40318 );
xor ( n40321 , n39119 , n39380 );
nor ( n40322 , n16669 , n40234 );
and ( n40323 , n40321 , n40322 );
xor ( n40324 , n40321 , n40322 );
xor ( n40325 , n39123 , n39378 );
nor ( n40326 , n15809 , n40234 );
and ( n40327 , n40325 , n40326 );
xor ( n40328 , n40325 , n40326 );
xor ( n40329 , n39127 , n39376 );
nor ( n40330 , n14968 , n40234 );
and ( n40331 , n40329 , n40330 );
xor ( n40332 , n40329 , n40330 );
xor ( n40333 , n39131 , n39374 );
nor ( n40334 , n14147 , n40234 );
and ( n40335 , n40333 , n40334 );
xor ( n40336 , n40333 , n40334 );
xor ( n40337 , n39135 , n39372 );
nor ( n40338 , n13349 , n40234 );
and ( n40339 , n40337 , n40338 );
xor ( n40340 , n40337 , n40338 );
xor ( n40341 , n39139 , n39370 );
nor ( n40342 , n12564 , n40234 );
and ( n40343 , n40341 , n40342 );
xor ( n40344 , n40341 , n40342 );
xor ( n40345 , n39143 , n39368 );
nor ( n40346 , n11799 , n40234 );
and ( n40347 , n40345 , n40346 );
xor ( n40348 , n40345 , n40346 );
xor ( n40349 , n39147 , n39366 );
nor ( n40350 , n11050 , n40234 );
and ( n40351 , n40349 , n40350 );
xor ( n40352 , n40349 , n40350 );
xor ( n40353 , n39151 , n39364 );
nor ( n40354 , n10321 , n40234 );
and ( n40355 , n40353 , n40354 );
xor ( n40356 , n40353 , n40354 );
xor ( n40357 , n39155 , n39362 );
nor ( n40358 , n9429 , n40234 );
and ( n40359 , n40357 , n40358 );
xor ( n40360 , n40357 , n40358 );
xor ( n40361 , n39159 , n39360 );
nor ( n40362 , n8949 , n40234 );
and ( n40363 , n40361 , n40362 );
xor ( n40364 , n40361 , n40362 );
xor ( n40365 , n39163 , n39358 );
nor ( n40366 , n9437 , n40234 );
and ( n40367 , n40365 , n40366 );
xor ( n40368 , n40365 , n40366 );
xor ( n40369 , n39167 , n39356 );
nor ( n40370 , n9446 , n40234 );
and ( n40371 , n40369 , n40370 );
xor ( n40372 , n40369 , n40370 );
xor ( n40373 , n39171 , n39354 );
nor ( n40374 , n9455 , n40234 );
and ( n40375 , n40373 , n40374 );
xor ( n40376 , n40373 , n40374 );
xor ( n40377 , n39175 , n39352 );
nor ( n40378 , n9464 , n40234 );
and ( n40379 , n40377 , n40378 );
xor ( n40380 , n40377 , n40378 );
xor ( n40381 , n39179 , n39350 );
nor ( n40382 , n9473 , n40234 );
and ( n40383 , n40381 , n40382 );
xor ( n40384 , n40381 , n40382 );
xor ( n40385 , n39183 , n39348 );
nor ( n40386 , n9482 , n40234 );
and ( n40387 , n40385 , n40386 );
xor ( n40388 , n40385 , n40386 );
xor ( n40389 , n39187 , n39346 );
nor ( n40390 , n9491 , n40234 );
and ( n40391 , n40389 , n40390 );
xor ( n40392 , n40389 , n40390 );
xor ( n40393 , n39191 , n39344 );
nor ( n40394 , n9500 , n40234 );
and ( n40395 , n40393 , n40394 );
xor ( n40396 , n40393 , n40394 );
xor ( n40397 , n39195 , n39342 );
nor ( n40398 , n9509 , n40234 );
and ( n40399 , n40397 , n40398 );
xor ( n40400 , n40397 , n40398 );
xor ( n40401 , n39199 , n39340 );
nor ( n40402 , n9518 , n40234 );
and ( n40403 , n40401 , n40402 );
xor ( n40404 , n40401 , n40402 );
xor ( n40405 , n39203 , n39338 );
nor ( n40406 , n9527 , n40234 );
and ( n40407 , n40405 , n40406 );
xor ( n40408 , n40405 , n40406 );
xor ( n40409 , n39207 , n39336 );
nor ( n40410 , n9536 , n40234 );
and ( n40411 , n40409 , n40410 );
xor ( n40412 , n40409 , n40410 );
xor ( n40413 , n39211 , n39334 );
nor ( n40414 , n9545 , n40234 );
and ( n40415 , n40413 , n40414 );
xor ( n40416 , n40413 , n40414 );
xor ( n40417 , n39215 , n39332 );
nor ( n40418 , n9554 , n40234 );
and ( n40419 , n40417 , n40418 );
xor ( n40420 , n40417 , n40418 );
xor ( n40421 , n39219 , n39330 );
nor ( n40422 , n9563 , n40234 );
and ( n40423 , n40421 , n40422 );
xor ( n40424 , n40421 , n40422 );
xor ( n40425 , n39223 , n39328 );
nor ( n40426 , n9572 , n40234 );
and ( n40427 , n40425 , n40426 );
xor ( n40428 , n40425 , n40426 );
xor ( n40429 , n39227 , n39326 );
nor ( n40430 , n9581 , n40234 );
and ( n40431 , n40429 , n40430 );
xor ( n40432 , n40429 , n40430 );
xor ( n40433 , n39231 , n39324 );
nor ( n40434 , n9590 , n40234 );
and ( n40435 , n40433 , n40434 );
xor ( n40436 , n40433 , n40434 );
xor ( n40437 , n39235 , n39322 );
nor ( n40438 , n9599 , n40234 );
and ( n40439 , n40437 , n40438 );
xor ( n40440 , n40437 , n40438 );
xor ( n40441 , n39239 , n39320 );
nor ( n40442 , n9608 , n40234 );
and ( n40443 , n40441 , n40442 );
xor ( n40444 , n40441 , n40442 );
xor ( n40445 , n39243 , n39318 );
nor ( n40446 , n9617 , n40234 );
and ( n40447 , n40445 , n40446 );
xor ( n40448 , n40445 , n40446 );
xor ( n40449 , n39247 , n39316 );
nor ( n40450 , n9626 , n40234 );
and ( n40451 , n40449 , n40450 );
xor ( n40452 , n40449 , n40450 );
xor ( n40453 , n39251 , n39314 );
nor ( n40454 , n9635 , n40234 );
and ( n40455 , n40453 , n40454 );
xor ( n40456 , n40453 , n40454 );
xor ( n40457 , n39255 , n39312 );
nor ( n40458 , n9644 , n40234 );
and ( n40459 , n40457 , n40458 );
xor ( n40460 , n40457 , n40458 );
xor ( n40461 , n39259 , n39310 );
nor ( n40462 , n9653 , n40234 );
and ( n40463 , n40461 , n40462 );
xor ( n40464 , n40461 , n40462 );
xor ( n40465 , n39263 , n39308 );
nor ( n40466 , n9662 , n40234 );
and ( n40467 , n40465 , n40466 );
xor ( n40468 , n40465 , n40466 );
xor ( n40469 , n39267 , n39306 );
nor ( n40470 , n9671 , n40234 );
and ( n40471 , n40469 , n40470 );
xor ( n40472 , n40469 , n40470 );
xor ( n40473 , n39271 , n39304 );
nor ( n40474 , n9680 , n40234 );
and ( n40475 , n40473 , n40474 );
xor ( n40476 , n40473 , n40474 );
xor ( n40477 , n39275 , n39302 );
nor ( n40478 , n9689 , n40234 );
and ( n40479 , n40477 , n40478 );
xor ( n40480 , n40477 , n40478 );
xor ( n40481 , n39279 , n39300 );
nor ( n40482 , n9698 , n40234 );
and ( n40483 , n40481 , n40482 );
xor ( n40484 , n40481 , n40482 );
xor ( n40485 , n39283 , n39298 );
nor ( n40486 , n9707 , n40234 );
and ( n40487 , n40485 , n40486 );
xor ( n40488 , n40485 , n40486 );
xor ( n40489 , n39287 , n39296 );
nor ( n40490 , n9716 , n40234 );
and ( n40491 , n40489 , n40490 );
xor ( n40492 , n40489 , n40490 );
xor ( n40493 , n39291 , n39294 );
nor ( n40494 , n9725 , n40234 );
and ( n40495 , n40493 , n40494 );
xor ( n40496 , n40493 , n40494 );
xor ( n40497 , n39292 , n39293 );
nor ( n40498 , n9734 , n40234 );
and ( n40499 , n40497 , n40498 );
xor ( n40500 , n40497 , n40498 );
nor ( n40501 , n9752 , n39029 );
nor ( n40502 , n9743 , n40234 );
and ( n40503 , n40501 , n40502 );
and ( n40504 , n40500 , n40503 );
or ( n40505 , n40499 , n40504 );
and ( n40506 , n40496 , n40505 );
or ( n40507 , n40495 , n40506 );
and ( n40508 , n40492 , n40507 );
or ( n40509 , n40491 , n40508 );
and ( n40510 , n40488 , n40509 );
or ( n40511 , n40487 , n40510 );
and ( n40512 , n40484 , n40511 );
or ( n40513 , n40483 , n40512 );
and ( n40514 , n40480 , n40513 );
or ( n40515 , n40479 , n40514 );
and ( n40516 , n40476 , n40515 );
or ( n40517 , n40475 , n40516 );
and ( n40518 , n40472 , n40517 );
or ( n40519 , n40471 , n40518 );
and ( n40520 , n40468 , n40519 );
or ( n40521 , n40467 , n40520 );
and ( n40522 , n40464 , n40521 );
or ( n40523 , n40463 , n40522 );
and ( n40524 , n40460 , n40523 );
or ( n40525 , n40459 , n40524 );
and ( n40526 , n40456 , n40525 );
or ( n40527 , n40455 , n40526 );
and ( n40528 , n40452 , n40527 );
or ( n40529 , n40451 , n40528 );
and ( n40530 , n40448 , n40529 );
or ( n40531 , n40447 , n40530 );
and ( n40532 , n40444 , n40531 );
or ( n40533 , n40443 , n40532 );
and ( n40534 , n40440 , n40533 );
or ( n40535 , n40439 , n40534 );
and ( n40536 , n40436 , n40535 );
or ( n40537 , n40435 , n40536 );
and ( n40538 , n40432 , n40537 );
or ( n40539 , n40431 , n40538 );
and ( n40540 , n40428 , n40539 );
or ( n40541 , n40427 , n40540 );
and ( n40542 , n40424 , n40541 );
or ( n40543 , n40423 , n40542 );
and ( n40544 , n40420 , n40543 );
or ( n40545 , n40419 , n40544 );
and ( n40546 , n40416 , n40545 );
or ( n40547 , n40415 , n40546 );
and ( n40548 , n40412 , n40547 );
or ( n40549 , n40411 , n40548 );
and ( n40550 , n40408 , n40549 );
or ( n40551 , n40407 , n40550 );
and ( n40552 , n40404 , n40551 );
or ( n40553 , n40403 , n40552 );
and ( n40554 , n40400 , n40553 );
or ( n40555 , n40399 , n40554 );
and ( n40556 , n40396 , n40555 );
or ( n40557 , n40395 , n40556 );
and ( n40558 , n40392 , n40557 );
or ( n40559 , n40391 , n40558 );
and ( n40560 , n40388 , n40559 );
or ( n40561 , n40387 , n40560 );
and ( n40562 , n40384 , n40561 );
or ( n40563 , n40383 , n40562 );
and ( n40564 , n40380 , n40563 );
or ( n40565 , n40379 , n40564 );
and ( n40566 , n40376 , n40565 );
or ( n40567 , n40375 , n40566 );
and ( n40568 , n40372 , n40567 );
or ( n40569 , n40371 , n40568 );
and ( n40570 , n40368 , n40569 );
or ( n40571 , n40367 , n40570 );
and ( n40572 , n40364 , n40571 );
or ( n40573 , n40363 , n40572 );
and ( n40574 , n40360 , n40573 );
or ( n40575 , n40359 , n40574 );
and ( n40576 , n40356 , n40575 );
or ( n40577 , n40355 , n40576 );
and ( n40578 , n40352 , n40577 );
or ( n40579 , n40351 , n40578 );
and ( n40580 , n40348 , n40579 );
or ( n40581 , n40347 , n40580 );
and ( n40582 , n40344 , n40581 );
or ( n40583 , n40343 , n40582 );
and ( n40584 , n40340 , n40583 );
or ( n40585 , n40339 , n40584 );
and ( n40586 , n40336 , n40585 );
or ( n40587 , n40335 , n40586 );
and ( n40588 , n40332 , n40587 );
or ( n40589 , n40331 , n40588 );
and ( n40590 , n40328 , n40589 );
or ( n40591 , n40327 , n40590 );
and ( n40592 , n40324 , n40591 );
or ( n40593 , n40323 , n40592 );
and ( n40594 , n40320 , n40593 );
or ( n40595 , n40319 , n40594 );
and ( n40596 , n40316 , n40595 );
or ( n40597 , n40315 , n40596 );
and ( n40598 , n40312 , n40597 );
or ( n40599 , n40311 , n40598 );
and ( n40600 , n40308 , n40599 );
or ( n40601 , n40307 , n40600 );
and ( n40602 , n40304 , n40601 );
or ( n40603 , n40303 , n40602 );
and ( n40604 , n40300 , n40603 );
or ( n40605 , n40299 , n40604 );
and ( n40606 , n40296 , n40605 );
or ( n40607 , n40295 , n40606 );
and ( n40608 , n40292 , n40607 );
or ( n40609 , n40291 , n40608 );
and ( n40610 , n40288 , n40609 );
or ( n40611 , n40287 , n40610 );
and ( n40612 , n40284 , n40611 );
or ( n40613 , n40283 , n40612 );
and ( n40614 , n40280 , n40613 );
or ( n40615 , n40279 , n40614 );
and ( n40616 , n40276 , n40615 );
or ( n40617 , n40275 , n40616 );
and ( n40618 , n40272 , n40617 );
or ( n40619 , n40271 , n40618 );
and ( n40620 , n40268 , n40619 );
or ( n40621 , n40267 , n40620 );
and ( n40622 , n40264 , n40621 );
or ( n40623 , n40263 , n40622 );
and ( n40624 , n40260 , n40623 );
or ( n40625 , n40259 , n40624 );
and ( n40626 , n40256 , n40625 );
or ( n40627 , n40255 , n40626 );
and ( n40628 , n40252 , n40627 );
or ( n40629 , n40251 , n40628 );
and ( n40630 , n40248 , n40629 );
or ( n40631 , n40247 , n40630 );
and ( n40632 , n40244 , n40631 );
or ( n40633 , n40243 , n40632 );
and ( n40634 , n40240 , n40633 );
or ( n40635 , n40239 , n40634 );
xor ( n40636 , n40236 , n40635 );
and ( n40637 , n33403 , n795 );
nor ( n40638 , n796 , n40637 );
nor ( n40639 , n868 , n32231 );
xor ( n40640 , n40638 , n40639 );
and ( n40641 , n39427 , n39428 );
and ( n40642 , n39429 , n39432 );
or ( n40643 , n40641 , n40642 );
xor ( n40644 , n40640 , n40643 );
nor ( n40645 , n958 , n31083 );
xor ( n40646 , n40644 , n40645 );
and ( n40647 , n39433 , n39434 );
and ( n40648 , n39435 , n39438 );
or ( n40649 , n40647 , n40648 );
xor ( n40650 , n40646 , n40649 );
nor ( n40651 , n1062 , n29948 );
xor ( n40652 , n40650 , n40651 );
and ( n40653 , n39439 , n39440 );
and ( n40654 , n39441 , n39444 );
or ( n40655 , n40653 , n40654 );
xor ( n40656 , n40652 , n40655 );
nor ( n40657 , n1176 , n28833 );
xor ( n40658 , n40656 , n40657 );
and ( n40659 , n39445 , n39446 );
and ( n40660 , n39447 , n39450 );
or ( n40661 , n40659 , n40660 );
xor ( n40662 , n40658 , n40661 );
nor ( n40663 , n1303 , n27737 );
xor ( n40664 , n40662 , n40663 );
and ( n40665 , n39451 , n39452 );
and ( n40666 , n39453 , n39456 );
or ( n40667 , n40665 , n40666 );
xor ( n40668 , n40664 , n40667 );
nor ( n40669 , n1445 , n26660 );
xor ( n40670 , n40668 , n40669 );
and ( n40671 , n39457 , n39458 );
and ( n40672 , n39459 , n39462 );
or ( n40673 , n40671 , n40672 );
xor ( n40674 , n40670 , n40673 );
nor ( n40675 , n1598 , n25600 );
xor ( n40676 , n40674 , n40675 );
and ( n40677 , n39463 , n39464 );
and ( n40678 , n39465 , n39468 );
or ( n40679 , n40677 , n40678 );
xor ( n40680 , n40676 , n40679 );
nor ( n40681 , n1766 , n24564 );
xor ( n40682 , n40680 , n40681 );
and ( n40683 , n39469 , n39470 );
and ( n40684 , n39471 , n39474 );
or ( n40685 , n40683 , n40684 );
xor ( n40686 , n40682 , n40685 );
nor ( n40687 , n1945 , n23541 );
xor ( n40688 , n40686 , n40687 );
and ( n40689 , n39475 , n39476 );
and ( n40690 , n39477 , n39480 );
or ( n40691 , n40689 , n40690 );
xor ( n40692 , n40688 , n40691 );
nor ( n40693 , n2137 , n22541 );
xor ( n40694 , n40692 , n40693 );
and ( n40695 , n39481 , n39482 );
and ( n40696 , n39483 , n39486 );
or ( n40697 , n40695 , n40696 );
xor ( n40698 , n40694 , n40697 );
nor ( n40699 , n2343 , n21562 );
xor ( n40700 , n40698 , n40699 );
and ( n40701 , n39487 , n39488 );
and ( n40702 , n39489 , n39492 );
or ( n40703 , n40701 , n40702 );
xor ( n40704 , n40700 , n40703 );
nor ( n40705 , n2566 , n20601 );
xor ( n40706 , n40704 , n40705 );
and ( n40707 , n39493 , n39494 );
and ( n40708 , n39495 , n39498 );
or ( n40709 , n40707 , n40708 );
xor ( n40710 , n40706 , n40709 );
nor ( n40711 , n2797 , n19657 );
xor ( n40712 , n40710 , n40711 );
and ( n40713 , n39499 , n39500 );
and ( n40714 , n39501 , n39504 );
or ( n40715 , n40713 , n40714 );
xor ( n40716 , n40712 , n40715 );
nor ( n40717 , n3043 , n18734 );
xor ( n40718 , n40716 , n40717 );
and ( n40719 , n39505 , n39506 );
and ( n40720 , n39507 , n39510 );
or ( n40721 , n40719 , n40720 );
xor ( n40722 , n40718 , n40721 );
nor ( n40723 , n3300 , n17828 );
xor ( n40724 , n40722 , n40723 );
and ( n40725 , n39511 , n39512 );
and ( n40726 , n39513 , n39516 );
or ( n40727 , n40725 , n40726 );
xor ( n40728 , n40724 , n40727 );
nor ( n40729 , n3570 , n16943 );
xor ( n40730 , n40728 , n40729 );
and ( n40731 , n39517 , n39518 );
and ( n40732 , n39519 , n39522 );
or ( n40733 , n40731 , n40732 );
xor ( n40734 , n40730 , n40733 );
nor ( n40735 , n3853 , n16077 );
xor ( n40736 , n40734 , n40735 );
and ( n40737 , n39523 , n39524 );
and ( n40738 , n39525 , n39528 );
or ( n40739 , n40737 , n40738 );
xor ( n40740 , n40736 , n40739 );
nor ( n40741 , n4151 , n15230 );
xor ( n40742 , n40740 , n40741 );
and ( n40743 , n39529 , n39530 );
and ( n40744 , n39531 , n39534 );
or ( n40745 , n40743 , n40744 );
xor ( n40746 , n40742 , n40745 );
nor ( n40747 , n4458 , n14403 );
xor ( n40748 , n40746 , n40747 );
and ( n40749 , n39535 , n39536 );
and ( n40750 , n39537 , n39540 );
or ( n40751 , n40749 , n40750 );
xor ( n40752 , n40748 , n40751 );
nor ( n40753 , n4786 , n13599 );
xor ( n40754 , n40752 , n40753 );
and ( n40755 , n39541 , n39542 );
and ( n40756 , n39543 , n39546 );
or ( n40757 , n40755 , n40756 );
xor ( n40758 , n40754 , n40757 );
nor ( n40759 , n5126 , n12808 );
xor ( n40760 , n40758 , n40759 );
and ( n40761 , n39547 , n39548 );
and ( n40762 , n39549 , n39552 );
or ( n40763 , n40761 , n40762 );
xor ( n40764 , n40760 , n40763 );
nor ( n40765 , n5477 , n12037 );
xor ( n40766 , n40764 , n40765 );
and ( n40767 , n39553 , n39554 );
and ( n40768 , n39555 , n39558 );
or ( n40769 , n40767 , n40768 );
xor ( n40770 , n40766 , n40769 );
nor ( n40771 , n5838 , n11282 );
xor ( n40772 , n40770 , n40771 );
and ( n40773 , n39559 , n39560 );
and ( n40774 , n39561 , n39564 );
or ( n40775 , n40773 , n40774 );
xor ( n40776 , n40772 , n40775 );
nor ( n40777 , n6212 , n10547 );
xor ( n40778 , n40776 , n40777 );
and ( n40779 , n39565 , n39566 );
and ( n40780 , n39567 , n39570 );
or ( n40781 , n40779 , n40780 );
xor ( n40782 , n40778 , n40781 );
nor ( n40783 , n6596 , n9829 );
xor ( n40784 , n40782 , n40783 );
and ( n40785 , n39571 , n39572 );
and ( n40786 , n39573 , n39576 );
or ( n40787 , n40785 , n40786 );
xor ( n40788 , n40784 , n40787 );
nor ( n40789 , n6997 , n8955 );
xor ( n40790 , n40788 , n40789 );
and ( n40791 , n39577 , n39578 );
and ( n40792 , n39579 , n39582 );
or ( n40793 , n40791 , n40792 );
xor ( n40794 , n40790 , n40793 );
nor ( n40795 , n7413 , n603 );
xor ( n40796 , n40794 , n40795 );
and ( n40797 , n39583 , n39584 );
and ( n40798 , n39585 , n39588 );
or ( n40799 , n40797 , n40798 );
xor ( n40800 , n40796 , n40799 );
nor ( n40801 , n7841 , n652 );
xor ( n40802 , n40800 , n40801 );
and ( n40803 , n39589 , n39590 );
and ( n40804 , n39591 , n39594 );
or ( n40805 , n40803 , n40804 );
xor ( n40806 , n40802 , n40805 );
nor ( n40807 , n8281 , n624 );
xor ( n40808 , n40806 , n40807 );
and ( n40809 , n39595 , n39596 );
and ( n40810 , n39597 , n39600 );
or ( n40811 , n40809 , n40810 );
xor ( n40812 , n40808 , n40811 );
nor ( n40813 , n8737 , n648 );
xor ( n40814 , n40812 , n40813 );
and ( n40815 , n39601 , n39602 );
and ( n40816 , n39603 , n39606 );
or ( n40817 , n40815 , n40816 );
xor ( n40818 , n40814 , n40817 );
nor ( n40819 , n9420 , n686 );
xor ( n40820 , n40818 , n40819 );
and ( n40821 , n39607 , n39608 );
and ( n40822 , n39609 , n39612 );
or ( n40823 , n40821 , n40822 );
xor ( n40824 , n40820 , n40823 );
nor ( n40825 , n10312 , n735 );
xor ( n40826 , n40824 , n40825 );
and ( n40827 , n39613 , n39614 );
and ( n40828 , n39615 , n39618 );
or ( n40829 , n40827 , n40828 );
xor ( n40830 , n40826 , n40829 );
nor ( n40831 , n11041 , n798 );
xor ( n40832 , n40830 , n40831 );
and ( n40833 , n39619 , n39620 );
and ( n40834 , n39621 , n39624 );
or ( n40835 , n40833 , n40834 );
xor ( n40836 , n40832 , n40835 );
nor ( n40837 , n11790 , n870 );
xor ( n40838 , n40836 , n40837 );
and ( n40839 , n39625 , n39626 );
and ( n40840 , n39627 , n39630 );
or ( n40841 , n40839 , n40840 );
xor ( n40842 , n40838 , n40841 );
nor ( n40843 , n12555 , n960 );
xor ( n40844 , n40842 , n40843 );
and ( n40845 , n39631 , n39632 );
and ( n40846 , n39633 , n39636 );
or ( n40847 , n40845 , n40846 );
xor ( n40848 , n40844 , n40847 );
nor ( n40849 , n13340 , n1064 );
xor ( n40850 , n40848 , n40849 );
and ( n40851 , n39637 , n39638 );
and ( n40852 , n39639 , n39642 );
or ( n40853 , n40851 , n40852 );
xor ( n40854 , n40850 , n40853 );
nor ( n40855 , n14138 , n1178 );
xor ( n40856 , n40854 , n40855 );
and ( n40857 , n39643 , n39644 );
and ( n40858 , n39645 , n39648 );
or ( n40859 , n40857 , n40858 );
xor ( n40860 , n40856 , n40859 );
nor ( n40861 , n14959 , n1305 );
xor ( n40862 , n40860 , n40861 );
and ( n40863 , n39649 , n39650 );
and ( n40864 , n39651 , n39654 );
or ( n40865 , n40863 , n40864 );
xor ( n40866 , n40862 , n40865 );
nor ( n40867 , n15800 , n1447 );
xor ( n40868 , n40866 , n40867 );
and ( n40869 , n39655 , n39656 );
and ( n40870 , n39657 , n39660 );
or ( n40871 , n40869 , n40870 );
xor ( n40872 , n40868 , n40871 );
nor ( n40873 , n16660 , n1600 );
xor ( n40874 , n40872 , n40873 );
and ( n40875 , n39661 , n39662 );
and ( n40876 , n39663 , n39666 );
or ( n40877 , n40875 , n40876 );
xor ( n40878 , n40874 , n40877 );
nor ( n40879 , n17539 , n1768 );
xor ( n40880 , n40878 , n40879 );
and ( n40881 , n39667 , n39668 );
and ( n40882 , n39669 , n39672 );
or ( n40883 , n40881 , n40882 );
xor ( n40884 , n40880 , n40883 );
nor ( n40885 , n18439 , n1947 );
xor ( n40886 , n40884 , n40885 );
and ( n40887 , n39673 , n39674 );
and ( n40888 , n39675 , n39678 );
or ( n40889 , n40887 , n40888 );
xor ( n40890 , n40886 , n40889 );
nor ( n40891 , n19356 , n2139 );
xor ( n40892 , n40890 , n40891 );
and ( n40893 , n39679 , n39680 );
and ( n40894 , n39681 , n39684 );
or ( n40895 , n40893 , n40894 );
xor ( n40896 , n40892 , n40895 );
nor ( n40897 , n20294 , n2345 );
xor ( n40898 , n40896 , n40897 );
and ( n40899 , n39685 , n39686 );
and ( n40900 , n39687 , n39690 );
or ( n40901 , n40899 , n40900 );
xor ( n40902 , n40898 , n40901 );
nor ( n40903 , n21249 , n2568 );
xor ( n40904 , n40902 , n40903 );
and ( n40905 , n39691 , n39692 );
and ( n40906 , n39693 , n39696 );
or ( n40907 , n40905 , n40906 );
xor ( n40908 , n40904 , n40907 );
nor ( n40909 , n22222 , n2799 );
xor ( n40910 , n40908 , n40909 );
and ( n40911 , n39697 , n39698 );
and ( n40912 , n39699 , n39702 );
or ( n40913 , n40911 , n40912 );
xor ( n40914 , n40910 , n40913 );
nor ( n40915 , n23216 , n3045 );
xor ( n40916 , n40914 , n40915 );
and ( n40917 , n39703 , n39704 );
and ( n40918 , n39705 , n39708 );
or ( n40919 , n40917 , n40918 );
xor ( n40920 , n40916 , n40919 );
nor ( n40921 , n24233 , n3302 );
xor ( n40922 , n40920 , n40921 );
and ( n40923 , n39709 , n39710 );
and ( n40924 , n39711 , n39714 );
or ( n40925 , n40923 , n40924 );
xor ( n40926 , n40922 , n40925 );
nor ( n40927 , n25263 , n3572 );
xor ( n40928 , n40926 , n40927 );
and ( n40929 , n39715 , n39716 );
and ( n40930 , n39717 , n39720 );
or ( n40931 , n40929 , n40930 );
xor ( n40932 , n40928 , n40931 );
nor ( n40933 , n26317 , n3855 );
xor ( n40934 , n40932 , n40933 );
and ( n40935 , n39721 , n39722 );
and ( n40936 , n39723 , n39726 );
or ( n40937 , n40935 , n40936 );
xor ( n40938 , n40934 , n40937 );
nor ( n40939 , n27388 , n4153 );
xor ( n40940 , n40938 , n40939 );
and ( n40941 , n39727 , n39728 );
and ( n40942 , n39729 , n39732 );
or ( n40943 , n40941 , n40942 );
xor ( n40944 , n40940 , n40943 );
nor ( n40945 , n28478 , n4460 );
xor ( n40946 , n40944 , n40945 );
and ( n40947 , n39733 , n39734 );
and ( n40948 , n39735 , n39738 );
or ( n40949 , n40947 , n40948 );
xor ( n40950 , n40946 , n40949 );
nor ( n40951 , n29587 , n4788 );
xor ( n40952 , n40950 , n40951 );
and ( n40953 , n39739 , n39740 );
and ( n40954 , n39741 , n39744 );
or ( n40955 , n40953 , n40954 );
xor ( n40956 , n40952 , n40955 );
nor ( n40957 , n30716 , n5128 );
xor ( n40958 , n40956 , n40957 );
and ( n40959 , n39745 , n39746 );
and ( n40960 , n39747 , n39750 );
or ( n40961 , n40959 , n40960 );
xor ( n40962 , n40958 , n40961 );
nor ( n40963 , n31858 , n5479 );
xor ( n40964 , n40962 , n40963 );
and ( n40965 , n39751 , n39752 );
and ( n40966 , n39753 , n39756 );
or ( n40967 , n40965 , n40966 );
xor ( n40968 , n40964 , n40967 );
nor ( n40969 , n33024 , n5840 );
xor ( n40970 , n40968 , n40969 );
and ( n40971 , n39757 , n39758 );
and ( n40972 , n39759 , n39762 );
or ( n40973 , n40971 , n40972 );
xor ( n40974 , n40970 , n40973 );
nor ( n40975 , n34215 , n6214 );
xor ( n40976 , n40974 , n40975 );
and ( n40977 , n39763 , n39764 );
and ( n40978 , n39765 , n39768 );
or ( n40979 , n40977 , n40978 );
xor ( n40980 , n40976 , n40979 );
nor ( n40981 , n35410 , n6598 );
xor ( n40982 , n40980 , n40981 );
and ( n40983 , n39769 , n39770 );
and ( n40984 , n39771 , n39774 );
or ( n40985 , n40983 , n40984 );
xor ( n40986 , n40982 , n40985 );
nor ( n40987 , n36611 , n6999 );
xor ( n40988 , n40986 , n40987 );
and ( n40989 , n39775 , n39776 );
and ( n40990 , n39777 , n39780 );
or ( n40991 , n40989 , n40990 );
xor ( n40992 , n40988 , n40991 );
nor ( n40993 , n37816 , n7415 );
xor ( n40994 , n40992 , n40993 );
and ( n40995 , n39781 , n39782 );
and ( n40996 , n39783 , n39786 );
or ( n40997 , n40995 , n40996 );
xor ( n40998 , n40994 , n40997 );
nor ( n40999 , n39018 , n7843 );
xor ( n41000 , n40998 , n40999 );
and ( n41001 , n39787 , n39788 );
and ( n41002 , n39789 , n39792 );
or ( n41003 , n41001 , n41002 );
xor ( n41004 , n41000 , n41003 );
nor ( n41005 , n40223 , n8283 );
xor ( n41006 , n41004 , n41005 );
and ( n41007 , n39793 , n39794 );
and ( n41008 , n39795 , n39798 );
or ( n41009 , n41007 , n41008 );
xor ( n41010 , n41006 , n41009 );
and ( n41011 , n39811 , n39815 );
and ( n41012 , n39815 , n40209 );
and ( n41013 , n39811 , n40209 );
or ( n41014 , n41011 , n41012 , n41013 );
and ( n41015 , n33774 , n771 );
not ( n41016 , n771 );
nor ( n41017 , n41015 , n41016 );
xor ( n41018 , n41014 , n41017 );
and ( n41019 , n39824 , n39828 );
and ( n41020 , n39828 , n39896 );
and ( n41021 , n39824 , n39896 );
or ( n41022 , n41019 , n41020 , n41021 );
and ( n41023 , n39820 , n39897 );
and ( n41024 , n39897 , n40208 );
and ( n41025 , n39820 , n40208 );
or ( n41026 , n41023 , n41024 , n41025 );
xor ( n41027 , n41022 , n41026 );
and ( n41028 , n39902 , n40022 );
and ( n41029 , n40022 , n40207 );
and ( n41030 , n39902 , n40207 );
or ( n41031 , n41028 , n41029 , n41030 );
and ( n41032 , n39833 , n39837 );
and ( n41033 , n39837 , n39895 );
and ( n41034 , n39833 , n39895 );
or ( n41035 , n41032 , n41033 , n41034 );
and ( n41036 , n39906 , n39910 );
and ( n41037 , n39910 , n40021 );
and ( n41038 , n39906 , n40021 );
or ( n41039 , n41036 , n41037 , n41038 );
xor ( n41040 , n41035 , n41039 );
and ( n41041 , n39864 , n39868 );
and ( n41042 , n39868 , n39874 );
and ( n41043 , n39864 , n39874 );
or ( n41044 , n41041 , n41042 , n41043 );
and ( n41045 , n39842 , n39846 );
and ( n41046 , n39846 , n39894 );
and ( n41047 , n39842 , n39894 );
or ( n41048 , n41045 , n41046 , n41047 );
xor ( n41049 , n41044 , n41048 );
and ( n41050 , n39851 , n39855 );
and ( n41051 , n39855 , n39893 );
and ( n41052 , n39851 , n39893 );
or ( n41053 , n41050 , n41051 , n41052 );
and ( n41054 , n39919 , n39944 );
and ( n41055 , n39944 , n39982 );
and ( n41056 , n39919 , n39982 );
or ( n41057 , n41054 , n41055 , n41056 );
xor ( n41058 , n41053 , n41057 );
and ( n41059 , n39860 , n39875 );
and ( n41060 , n39875 , n39892 );
and ( n41061 , n39860 , n39892 );
or ( n41062 , n41059 , n41060 , n41061 );
and ( n41063 , n39923 , n39927 );
and ( n41064 , n39927 , n39943 );
and ( n41065 , n39923 , n39943 );
or ( n41066 , n41063 , n41064 , n41065 );
xor ( n41067 , n41062 , n41066 );
and ( n41068 , n39880 , n39885 );
and ( n41069 , n39885 , n39891 );
and ( n41070 , n39880 , n39891 );
or ( n41071 , n41068 , n41069 , n41070 );
and ( n41072 , n39870 , n39871 );
and ( n41073 , n39871 , n39873 );
and ( n41074 , n39870 , n39873 );
or ( n41075 , n41072 , n41073 , n41074 );
and ( n41076 , n39881 , n39882 );
and ( n41077 , n39882 , n39884 );
and ( n41078 , n39881 , n39884 );
or ( n41079 , n41076 , n41077 , n41078 );
xor ( n41080 , n41075 , n41079 );
and ( n41081 , n30695 , n1034 );
and ( n41082 , n31836 , n940 );
xor ( n41083 , n41081 , n41082 );
and ( n41084 , n32649 , n840 );
xor ( n41085 , n41083 , n41084 );
xor ( n41086 , n41080 , n41085 );
xor ( n41087 , n41071 , n41086 );
and ( n41088 , n39887 , n39888 );
and ( n41089 , n39888 , n39890 );
and ( n41090 , n39887 , n39890 );
or ( n41091 , n41088 , n41089 , n41090 );
and ( n41092 , n27361 , n1424 );
and ( n41093 , n28456 , n1254 );
xor ( n41094 , n41092 , n41093 );
and ( n41095 , n29559 , n1134 );
xor ( n41096 , n41094 , n41095 );
xor ( n41097 , n41091 , n41096 );
and ( n41098 , n24214 , n1882 );
and ( n41099 , n25243 , n1738 );
xor ( n41100 , n41098 , n41099 );
and ( n41101 , n26296 , n1551 );
xor ( n41102 , n41100 , n41101 );
xor ( n41103 , n41097 , n41102 );
xor ( n41104 , n41087 , n41103 );
xor ( n41105 , n41067 , n41104 );
xor ( n41106 , n41058 , n41105 );
xor ( n41107 , n41049 , n41106 );
xor ( n41108 , n41040 , n41107 );
xor ( n41109 , n41031 , n41108 );
and ( n41110 , n40027 , n40107 );
and ( n41111 , n40107 , n40206 );
and ( n41112 , n40027 , n40206 );
or ( n41113 , n41110 , n41111 , n41112 );
and ( n41114 , n39915 , n39983 );
and ( n41115 , n39983 , n40020 );
and ( n41116 , n39915 , n40020 );
or ( n41117 , n41114 , n41115 , n41116 );
and ( n41118 , n40031 , n40035 );
and ( n41119 , n40035 , n40106 );
and ( n41120 , n40031 , n40106 );
or ( n41121 , n41118 , n41119 , n41120 );
xor ( n41122 , n41117 , n41121 );
and ( n41123 , n39988 , n39992 );
and ( n41124 , n39992 , n40019 );
and ( n41125 , n39988 , n40019 );
or ( n41126 , n41123 , n41124 , n41125 );
and ( n41127 , n39949 , n39965 );
and ( n41128 , n39965 , n39981 );
and ( n41129 , n39949 , n39981 );
or ( n41130 , n41127 , n41128 , n41129 );
and ( n41131 , n39932 , n39936 );
and ( n41132 , n39936 , n39942 );
and ( n41133 , n39932 , n39942 );
or ( n41134 , n41131 , n41132 , n41133 );
and ( n41135 , n39953 , n39958 );
and ( n41136 , n39958 , n39964 );
and ( n41137 , n39953 , n39964 );
or ( n41138 , n41135 , n41136 , n41137 );
xor ( n41139 , n41134 , n41138 );
and ( n41140 , n39938 , n39939 );
and ( n41141 , n39939 , n39941 );
and ( n41142 , n39938 , n39941 );
or ( n41143 , n41140 , n41141 , n41142 );
and ( n41144 , n39954 , n39955 );
and ( n41145 , n39955 , n39957 );
and ( n41146 , n39954 , n39957 );
or ( n41147 , n41144 , n41145 , n41146 );
xor ( n41148 , n41143 , n41147 );
and ( n41149 , n21216 , n2544 );
and ( n41150 , n22186 , n2298 );
xor ( n41151 , n41149 , n41150 );
and ( n41152 , n22892 , n2100 );
xor ( n41153 , n41151 , n41152 );
xor ( n41154 , n41148 , n41153 );
xor ( n41155 , n41139 , n41154 );
xor ( n41156 , n41130 , n41155 );
and ( n41157 , n39970 , n39974 );
and ( n41158 , n39974 , n39980 );
and ( n41159 , n39970 , n39980 );
or ( n41160 , n41157 , n41158 , n41159 );
and ( n41161 , n39960 , n39961 );
and ( n41162 , n39961 , n39963 );
and ( n41163 , n39960 , n39963 );
or ( n41164 , n41161 , n41162 , n41163 );
and ( n41165 , n18144 , n3271 );
and ( n41166 , n19324 , n2981 );
xor ( n41167 , n41165 , n41166 );
and ( n41168 , n20233 , n2739 );
xor ( n41169 , n41167 , n41168 );
xor ( n41170 , n41164 , n41169 );
and ( n41171 , n15758 , n4102 );
and ( n41172 , n16637 , n3749 );
xor ( n41173 , n41171 , n41172 );
and ( n41174 , n17512 , n3495 );
xor ( n41175 , n41173 , n41174 );
xor ( n41176 , n41170 , n41175 );
xor ( n41177 , n41160 , n41176 );
and ( n41178 , n39976 , n39977 );
and ( n41179 , n39977 , n39979 );
and ( n41180 , n39976 , n39979 );
or ( n41181 , n41178 , n41179 , n41180 );
and ( n41182 , n40007 , n40008 );
and ( n41183 , n40008 , n40010 );
and ( n41184 , n40007 , n40010 );
or ( n41185 , n41182 , n41183 , n41184 );
xor ( n41186 , n41181 , n41185 );
and ( n41187 , n13322 , n5103 );
and ( n41188 , n14118 , n4730 );
xor ( n41189 , n41187 , n41188 );
and ( n41190 , n14938 , n4403 );
xor ( n41191 , n41189 , n41190 );
xor ( n41192 , n41186 , n41191 );
xor ( n41193 , n41177 , n41192 );
xor ( n41194 , n41156 , n41193 );
xor ( n41195 , n41126 , n41194 );
and ( n41196 , n39997 , n40001 );
and ( n41197 , n40001 , n40018 );
and ( n41198 , n39997 , n40018 );
or ( n41199 , n41196 , n41197 , n41198 );
and ( n41200 , n40044 , n40061 );
and ( n41201 , n40061 , n40078 );
and ( n41202 , n40044 , n40078 );
or ( n41203 , n41200 , n41201 , n41202 );
xor ( n41204 , n41199 , n41203 );
and ( n41205 , n40006 , n40011 );
and ( n41206 , n40011 , n40017 );
and ( n41207 , n40006 , n40017 );
or ( n41208 , n41205 , n41206 , n41207 );
and ( n41209 , n40050 , n40054 );
and ( n41210 , n40054 , n40060 );
and ( n41211 , n40050 , n40060 );
or ( n41212 , n41209 , n41210 , n41211 );
xor ( n41213 , n41208 , n41212 );
and ( n41214 , n40013 , n40014 );
and ( n41215 , n40014 , n40016 );
and ( n41216 , n40013 , n40016 );
or ( n41217 , n41214 , n41215 , n41216 );
and ( n41218 , n11015 , n6132 );
and ( n41219 , n11769 , n5765 );
xor ( n41220 , n41218 , n41219 );
and ( n41221 , n12320 , n5408 );
xor ( n41222 , n41220 , n41221 );
xor ( n41223 , n41217 , n41222 );
and ( n41224 , n8718 , n7310 );
and ( n41225 , n9400 , n6971 );
xor ( n41226 , n41224 , n41225 );
and ( n41227 , n10291 , n6504 );
xor ( n41228 , n41226 , n41227 );
xor ( n41229 , n41223 , n41228 );
xor ( n41230 , n41213 , n41229 );
xor ( n41231 , n41204 , n41230 );
xor ( n41232 , n41195 , n41231 );
xor ( n41233 , n41122 , n41232 );
xor ( n41234 , n41113 , n41233 );
and ( n41235 , n40112 , n40159 );
and ( n41236 , n40159 , n40205 );
and ( n41237 , n40112 , n40205 );
or ( n41238 , n41235 , n41236 , n41237 );
and ( n41239 , n40040 , n40079 );
and ( n41240 , n40079 , n40105 );
and ( n41241 , n40040 , n40105 );
or ( n41242 , n41239 , n41240 , n41241 );
and ( n41243 , n40116 , n40120 );
and ( n41244 , n40120 , n40158 );
and ( n41245 , n40116 , n40158 );
or ( n41246 , n41243 , n41244 , n41245 );
xor ( n41247 , n41242 , n41246 );
and ( n41248 , n40084 , n40088 );
and ( n41249 , n40088 , n40104 );
and ( n41250 , n40084 , n40104 );
or ( n41251 , n41248 , n41249 , n41250 );
and ( n41252 , n40066 , n40071 );
and ( n41253 , n40071 , n40077 );
and ( n41254 , n40066 , n40077 );
or ( n41255 , n41252 , n41253 , n41254 );
and ( n41256 , n40056 , n40057 );
and ( n41257 , n40057 , n40059 );
and ( n41258 , n40056 , n40059 );
or ( n41259 , n41256 , n41257 , n41258 );
and ( n41260 , n40067 , n40068 );
and ( n41261 , n40068 , n40070 );
and ( n41262 , n40067 , n40070 );
or ( n41263 , n41260 , n41261 , n41262 );
xor ( n41264 , n41259 , n41263 );
and ( n41265 , n7385 , n8669 );
and ( n41266 , n7808 , n8243 );
xor ( n41267 , n41265 , n41266 );
and ( n41268 , n8079 , n7662 );
xor ( n41269 , n41267 , n41268 );
xor ( n41270 , n41264 , n41269 );
xor ( n41271 , n41255 , n41270 );
and ( n41272 , n40073 , n40074 );
and ( n41273 , n40074 , n40076 );
and ( n41274 , n40073 , n40076 );
or ( n41275 , n41272 , n41273 , n41274 );
and ( n41276 , n6187 , n10977 );
and ( n41277 , n6569 , n10239 );
xor ( n41278 , n41276 , n41277 );
and ( n41279 , n6816 , n9348 );
xor ( n41280 , n41278 , n41279 );
xor ( n41281 , n41275 , n41280 );
and ( n41282 , n4959 , n13256 );
and ( n41283 , n5459 , n12531 );
xor ( n41284 , n41282 , n41283 );
and ( n41285 , n5819 , n11718 );
xor ( n41286 , n41284 , n41285 );
xor ( n41287 , n41281 , n41286 );
xor ( n41288 , n41271 , n41287 );
xor ( n41289 , n41251 , n41288 );
and ( n41290 , n40093 , n40097 );
and ( n41291 , n40097 , n40103 );
and ( n41292 , n40093 , n40103 );
or ( n41293 , n41290 , n41291 , n41292 );
and ( n41294 , n40129 , n40134 );
and ( n41295 , n40134 , n40140 );
and ( n41296 , n40129 , n40140 );
or ( n41297 , n41294 , n41295 , n41296 );
xor ( n41298 , n41293 , n41297 );
and ( n41299 , n40099 , n40100 );
and ( n41300 , n40100 , n40102 );
and ( n41301 , n40099 , n40102 );
or ( n41302 , n41299 , n41300 , n41301 );
and ( n41303 , n40130 , n40131 );
and ( n41304 , n40131 , n40133 );
and ( n41305 , n40130 , n40133 );
or ( n41306 , n41303 , n41304 , n41305 );
xor ( n41307 , n41302 , n41306 );
and ( n41308 , n4132 , n15691 );
and ( n41309 , n4438 , n14838 );
xor ( n41310 , n41308 , n41309 );
and ( n41311 , n4766 , n14044 );
xor ( n41312 , n41310 , n41311 );
xor ( n41313 , n41307 , n41312 );
xor ( n41314 , n41298 , n41313 );
xor ( n41315 , n41289 , n41314 );
xor ( n41316 , n41247 , n41315 );
xor ( n41317 , n41238 , n41316 );
and ( n41318 , n40161 , n40187 );
and ( n41319 , n40187 , n40204 );
and ( n41320 , n40161 , n40204 );
or ( n41321 , n41318 , n41319 , n41320 );
and ( n41322 , n40125 , n40141 );
and ( n41323 , n40141 , n40157 );
and ( n41324 , n40125 , n40157 );
or ( n41325 , n41322 , n41323 , n41324 );
and ( n41326 , n40165 , n40169 );
and ( n41327 , n40169 , n40186 );
and ( n41328 , n40165 , n40186 );
or ( n41329 , n41326 , n41327 , n41328 );
xor ( n41330 , n41325 , n41329 );
and ( n41331 , n40146 , n40150 );
and ( n41332 , n40150 , n40156 );
and ( n41333 , n40146 , n40156 );
or ( n41334 , n41331 , n41332 , n41333 );
and ( n41335 , n40136 , n40137 );
and ( n41336 , n40137 , n40139 );
and ( n41337 , n40136 , n40139 );
or ( n41338 , n41335 , n41336 , n41337 );
and ( n41339 , n3182 , n18407 );
and ( n41340 , n3545 , n17422 );
xor ( n41341 , n41339 , n41340 );
and ( n41342 , n3801 , n16550 );
xor ( n41343 , n41341 , n41342 );
xor ( n41344 , n41338 , n41343 );
and ( n41345 , n2462 , n20976 );
and ( n41346 , n2779 , n20156 );
xor ( n41347 , n41345 , n41346 );
and ( n41348 , n3024 , n19222 );
xor ( n41349 , n41347 , n41348 );
xor ( n41350 , n41344 , n41349 );
xor ( n41351 , n41334 , n41350 );
and ( n41352 , n40152 , n40153 );
and ( n41353 , n40153 , n40155 );
and ( n41354 , n40152 , n40155 );
or ( n41355 , n41352 , n41353 , n41354 );
and ( n41356 , n40175 , n40176 );
and ( n41357 , n40176 , n40178 );
and ( n41358 , n40175 , n40178 );
or ( n41359 , n41356 , n41357 , n41358 );
xor ( n41360 , n41355 , n41359 );
and ( n41361 , n1933 , n24137 );
and ( n41362 , n2120 , n23075 );
xor ( n41363 , n41361 , n41362 );
and ( n41364 , n2324 , n22065 );
xor ( n41365 , n41363 , n41364 );
xor ( n41366 , n41360 , n41365 );
xor ( n41367 , n41351 , n41366 );
xor ( n41368 , n41330 , n41367 );
xor ( n41369 , n41321 , n41368 );
and ( n41370 , n40191 , n40203 );
and ( n41371 , n40195 , n40196 );
and ( n41372 , n40196 , n40202 );
and ( n41373 , n40195 , n40202 );
or ( n41374 , n41371 , n41372 , n41373 );
and ( n41375 , n40174 , n40179 );
and ( n41376 , n40179 , n40185 );
and ( n41377 , n40174 , n40185 );
or ( n41378 , n41375 , n41376 , n41377 );
xor ( n41379 , n41374 , n41378 );
and ( n41380 , n40181 , n40182 );
and ( n41381 , n40182 , n40184 );
and ( n41382 , n40181 , n40184 );
or ( n41383 , n41380 , n41381 , n41382 );
and ( n41384 , n1383 , n27296 );
and ( n41385 , n1580 , n26216 );
xor ( n41386 , n41384 , n41385 );
and ( n41387 , n1694 , n25163 );
xor ( n41388 , n41386 , n41387 );
xor ( n41389 , n41383 , n41388 );
and ( n41390 , n1047 , n30629 );
and ( n41391 , n1164 , n29508 );
xor ( n41392 , n41390 , n41391 );
and ( n41393 , n1287 , n28406 );
xor ( n41394 , n41392 , n41393 );
xor ( n41395 , n41389 , n41394 );
xor ( n41396 , n41379 , n41395 );
xor ( n41397 , n41370 , n41396 );
and ( n41398 , n40198 , n40199 );
and ( n41399 , n40199 , n40201 );
and ( n41400 , n40198 , n40201 );
or ( n41401 , n41398 , n41399 , n41400 );
not ( n41402 , n783 );
and ( n41403 , n34193 , n783 );
nor ( n41404 , n41402 , n41403 );
and ( n41405 , n856 , n32999 );
xor ( n41406 , n41404 , n41405 );
and ( n41407 , n925 , n31761 );
xor ( n41408 , n41406 , n41407 );
xor ( n41409 , n41401 , n41408 );
xor ( n41410 , n41397 , n41409 );
xor ( n41411 , n41369 , n41410 );
xor ( n41412 , n41317 , n41411 );
xor ( n41413 , n41234 , n41412 );
xor ( n41414 , n41109 , n41413 );
xor ( n41415 , n41027 , n41414 );
xor ( n41416 , n41018 , n41415 );
and ( n41417 , n39803 , n39806 );
and ( n41418 , n39806 , n40210 );
and ( n41419 , n39803 , n40210 );
or ( n41420 , n41417 , n41418 , n41419 );
xor ( n41421 , n41416 , n41420 );
and ( n41422 , n40211 , n40215 );
and ( n41423 , n40216 , n40219 );
or ( n41424 , n41422 , n41423 );
xor ( n41425 , n41421 , n41424 );
buf ( n41426 , n41425 );
buf ( n41427 , n41426 );
not ( n41428 , n41427 );
nor ( n41429 , n41428 , n8739 );
xor ( n41430 , n41010 , n41429 );
and ( n41431 , n39799 , n40224 );
and ( n41432 , n40225 , n40228 );
or ( n41433 , n41431 , n41432 );
xor ( n41434 , n41430 , n41433 );
buf ( n41435 , n41434 );
buf ( n41436 , n41435 );
not ( n41437 , n41436 );
buf ( n41438 , n568 );
not ( n41439 , n41438 );
nor ( n41440 , n41437 , n41439 );
xor ( n41441 , n40636 , n41440 );
xor ( n41442 , n40240 , n40633 );
nor ( n41443 , n40232 , n41439 );
and ( n41444 , n41442 , n41443 );
xor ( n41445 , n41442 , n41443 );
xor ( n41446 , n40244 , n40631 );
nor ( n41447 , n39027 , n41439 );
and ( n41448 , n41446 , n41447 );
xor ( n41449 , n41446 , n41447 );
xor ( n41450 , n40248 , n40629 );
nor ( n41451 , n37825 , n41439 );
and ( n41452 , n41450 , n41451 );
xor ( n41453 , n41450 , n41451 );
xor ( n41454 , n40252 , n40627 );
nor ( n41455 , n36620 , n41439 );
and ( n41456 , n41454 , n41455 );
xor ( n41457 , n41454 , n41455 );
xor ( n41458 , n40256 , n40625 );
nor ( n41459 , n35419 , n41439 );
and ( n41460 , n41458 , n41459 );
xor ( n41461 , n41458 , n41459 );
xor ( n41462 , n40260 , n40623 );
nor ( n41463 , n34224 , n41439 );
and ( n41464 , n41462 , n41463 );
xor ( n41465 , n41462 , n41463 );
xor ( n41466 , n40264 , n40621 );
nor ( n41467 , n33033 , n41439 );
and ( n41468 , n41466 , n41467 );
xor ( n41469 , n41466 , n41467 );
xor ( n41470 , n40268 , n40619 );
nor ( n41471 , n31867 , n41439 );
and ( n41472 , n41470 , n41471 );
xor ( n41473 , n41470 , n41471 );
xor ( n41474 , n40272 , n40617 );
nor ( n41475 , n30725 , n41439 );
and ( n41476 , n41474 , n41475 );
xor ( n41477 , n41474 , n41475 );
xor ( n41478 , n40276 , n40615 );
nor ( n41479 , n29596 , n41439 );
and ( n41480 , n41478 , n41479 );
xor ( n41481 , n41478 , n41479 );
xor ( n41482 , n40280 , n40613 );
nor ( n41483 , n28487 , n41439 );
and ( n41484 , n41482 , n41483 );
xor ( n41485 , n41482 , n41483 );
xor ( n41486 , n40284 , n40611 );
nor ( n41487 , n27397 , n41439 );
and ( n41488 , n41486 , n41487 );
xor ( n41489 , n41486 , n41487 );
xor ( n41490 , n40288 , n40609 );
nor ( n41491 , n26326 , n41439 );
and ( n41492 , n41490 , n41491 );
xor ( n41493 , n41490 , n41491 );
xor ( n41494 , n40292 , n40607 );
nor ( n41495 , n25272 , n41439 );
and ( n41496 , n41494 , n41495 );
xor ( n41497 , n41494 , n41495 );
xor ( n41498 , n40296 , n40605 );
nor ( n41499 , n24242 , n41439 );
and ( n41500 , n41498 , n41499 );
xor ( n41501 , n41498 , n41499 );
xor ( n41502 , n40300 , n40603 );
nor ( n41503 , n23225 , n41439 );
and ( n41504 , n41502 , n41503 );
xor ( n41505 , n41502 , n41503 );
xor ( n41506 , n40304 , n40601 );
nor ( n41507 , n22231 , n41439 );
and ( n41508 , n41506 , n41507 );
xor ( n41509 , n41506 , n41507 );
xor ( n41510 , n40308 , n40599 );
nor ( n41511 , n21258 , n41439 );
and ( n41512 , n41510 , n41511 );
xor ( n41513 , n41510 , n41511 );
xor ( n41514 , n40312 , n40597 );
nor ( n41515 , n20303 , n41439 );
and ( n41516 , n41514 , n41515 );
xor ( n41517 , n41514 , n41515 );
xor ( n41518 , n40316 , n40595 );
nor ( n41519 , n19365 , n41439 );
and ( n41520 , n41518 , n41519 );
xor ( n41521 , n41518 , n41519 );
xor ( n41522 , n40320 , n40593 );
nor ( n41523 , n18448 , n41439 );
and ( n41524 , n41522 , n41523 );
xor ( n41525 , n41522 , n41523 );
xor ( n41526 , n40324 , n40591 );
nor ( n41527 , n17548 , n41439 );
and ( n41528 , n41526 , n41527 );
xor ( n41529 , n41526 , n41527 );
xor ( n41530 , n40328 , n40589 );
nor ( n41531 , n16669 , n41439 );
and ( n41532 , n41530 , n41531 );
xor ( n41533 , n41530 , n41531 );
xor ( n41534 , n40332 , n40587 );
nor ( n41535 , n15809 , n41439 );
and ( n41536 , n41534 , n41535 );
xor ( n41537 , n41534 , n41535 );
xor ( n41538 , n40336 , n40585 );
nor ( n41539 , n14968 , n41439 );
and ( n41540 , n41538 , n41539 );
xor ( n41541 , n41538 , n41539 );
xor ( n41542 , n40340 , n40583 );
nor ( n41543 , n14147 , n41439 );
and ( n41544 , n41542 , n41543 );
xor ( n41545 , n41542 , n41543 );
xor ( n41546 , n40344 , n40581 );
nor ( n41547 , n13349 , n41439 );
and ( n41548 , n41546 , n41547 );
xor ( n41549 , n41546 , n41547 );
xor ( n41550 , n40348 , n40579 );
nor ( n41551 , n12564 , n41439 );
and ( n41552 , n41550 , n41551 );
xor ( n41553 , n41550 , n41551 );
xor ( n41554 , n40352 , n40577 );
nor ( n41555 , n11799 , n41439 );
and ( n41556 , n41554 , n41555 );
xor ( n41557 , n41554 , n41555 );
xor ( n41558 , n40356 , n40575 );
nor ( n41559 , n11050 , n41439 );
and ( n41560 , n41558 , n41559 );
xor ( n41561 , n41558 , n41559 );
xor ( n41562 , n40360 , n40573 );
nor ( n41563 , n10321 , n41439 );
and ( n41564 , n41562 , n41563 );
xor ( n41565 , n41562 , n41563 );
xor ( n41566 , n40364 , n40571 );
nor ( n41567 , n9429 , n41439 );
and ( n41568 , n41566 , n41567 );
xor ( n41569 , n41566 , n41567 );
xor ( n41570 , n40368 , n40569 );
nor ( n41571 , n8949 , n41439 );
and ( n41572 , n41570 , n41571 );
xor ( n41573 , n41570 , n41571 );
xor ( n41574 , n40372 , n40567 );
nor ( n41575 , n9437 , n41439 );
and ( n41576 , n41574 , n41575 );
xor ( n41577 , n41574 , n41575 );
xor ( n41578 , n40376 , n40565 );
nor ( n41579 , n9446 , n41439 );
and ( n41580 , n41578 , n41579 );
xor ( n41581 , n41578 , n41579 );
xor ( n41582 , n40380 , n40563 );
nor ( n41583 , n9455 , n41439 );
and ( n41584 , n41582 , n41583 );
xor ( n41585 , n41582 , n41583 );
xor ( n41586 , n40384 , n40561 );
nor ( n41587 , n9464 , n41439 );
and ( n41588 , n41586 , n41587 );
xor ( n41589 , n41586 , n41587 );
xor ( n41590 , n40388 , n40559 );
nor ( n41591 , n9473 , n41439 );
and ( n41592 , n41590 , n41591 );
xor ( n41593 , n41590 , n41591 );
xor ( n41594 , n40392 , n40557 );
nor ( n41595 , n9482 , n41439 );
and ( n41596 , n41594 , n41595 );
xor ( n41597 , n41594 , n41595 );
xor ( n41598 , n40396 , n40555 );
nor ( n41599 , n9491 , n41439 );
and ( n41600 , n41598 , n41599 );
xor ( n41601 , n41598 , n41599 );
xor ( n41602 , n40400 , n40553 );
nor ( n41603 , n9500 , n41439 );
and ( n41604 , n41602 , n41603 );
xor ( n41605 , n41602 , n41603 );
xor ( n41606 , n40404 , n40551 );
nor ( n41607 , n9509 , n41439 );
and ( n41608 , n41606 , n41607 );
xor ( n41609 , n41606 , n41607 );
xor ( n41610 , n40408 , n40549 );
nor ( n41611 , n9518 , n41439 );
and ( n41612 , n41610 , n41611 );
xor ( n41613 , n41610 , n41611 );
xor ( n41614 , n40412 , n40547 );
nor ( n41615 , n9527 , n41439 );
and ( n41616 , n41614 , n41615 );
xor ( n41617 , n41614 , n41615 );
xor ( n41618 , n40416 , n40545 );
nor ( n41619 , n9536 , n41439 );
and ( n41620 , n41618 , n41619 );
xor ( n41621 , n41618 , n41619 );
xor ( n41622 , n40420 , n40543 );
nor ( n41623 , n9545 , n41439 );
and ( n41624 , n41622 , n41623 );
xor ( n41625 , n41622 , n41623 );
xor ( n41626 , n40424 , n40541 );
nor ( n41627 , n9554 , n41439 );
and ( n41628 , n41626 , n41627 );
xor ( n41629 , n41626 , n41627 );
xor ( n41630 , n40428 , n40539 );
nor ( n41631 , n9563 , n41439 );
and ( n41632 , n41630 , n41631 );
xor ( n41633 , n41630 , n41631 );
xor ( n41634 , n40432 , n40537 );
nor ( n41635 , n9572 , n41439 );
and ( n41636 , n41634 , n41635 );
xor ( n41637 , n41634 , n41635 );
xor ( n41638 , n40436 , n40535 );
nor ( n41639 , n9581 , n41439 );
and ( n41640 , n41638 , n41639 );
xor ( n41641 , n41638 , n41639 );
xor ( n41642 , n40440 , n40533 );
nor ( n41643 , n9590 , n41439 );
and ( n41644 , n41642 , n41643 );
xor ( n41645 , n41642 , n41643 );
xor ( n41646 , n40444 , n40531 );
nor ( n41647 , n9599 , n41439 );
and ( n41648 , n41646 , n41647 );
xor ( n41649 , n41646 , n41647 );
xor ( n41650 , n40448 , n40529 );
nor ( n41651 , n9608 , n41439 );
and ( n41652 , n41650 , n41651 );
xor ( n41653 , n41650 , n41651 );
xor ( n41654 , n40452 , n40527 );
nor ( n41655 , n9617 , n41439 );
and ( n41656 , n41654 , n41655 );
xor ( n41657 , n41654 , n41655 );
xor ( n41658 , n40456 , n40525 );
nor ( n41659 , n9626 , n41439 );
and ( n41660 , n41658 , n41659 );
xor ( n41661 , n41658 , n41659 );
xor ( n41662 , n40460 , n40523 );
nor ( n41663 , n9635 , n41439 );
and ( n41664 , n41662 , n41663 );
xor ( n41665 , n41662 , n41663 );
xor ( n41666 , n40464 , n40521 );
nor ( n41667 , n9644 , n41439 );
and ( n41668 , n41666 , n41667 );
xor ( n41669 , n41666 , n41667 );
xor ( n41670 , n40468 , n40519 );
nor ( n41671 , n9653 , n41439 );
and ( n41672 , n41670 , n41671 );
xor ( n41673 , n41670 , n41671 );
xor ( n41674 , n40472 , n40517 );
nor ( n41675 , n9662 , n41439 );
and ( n41676 , n41674 , n41675 );
xor ( n41677 , n41674 , n41675 );
xor ( n41678 , n40476 , n40515 );
nor ( n41679 , n9671 , n41439 );
and ( n41680 , n41678 , n41679 );
xor ( n41681 , n41678 , n41679 );
xor ( n41682 , n40480 , n40513 );
nor ( n41683 , n9680 , n41439 );
and ( n41684 , n41682 , n41683 );
xor ( n41685 , n41682 , n41683 );
xor ( n41686 , n40484 , n40511 );
nor ( n41687 , n9689 , n41439 );
and ( n41688 , n41686 , n41687 );
xor ( n41689 , n41686 , n41687 );
xor ( n41690 , n40488 , n40509 );
nor ( n41691 , n9698 , n41439 );
and ( n41692 , n41690 , n41691 );
xor ( n41693 , n41690 , n41691 );
xor ( n41694 , n40492 , n40507 );
nor ( n41695 , n9707 , n41439 );
and ( n41696 , n41694 , n41695 );
xor ( n41697 , n41694 , n41695 );
xor ( n41698 , n40496 , n40505 );
nor ( n41699 , n9716 , n41439 );
and ( n41700 , n41698 , n41699 );
xor ( n41701 , n41698 , n41699 );
xor ( n41702 , n40500 , n40503 );
nor ( n41703 , n9725 , n41439 );
and ( n41704 , n41702 , n41703 );
xor ( n41705 , n41702 , n41703 );
xor ( n41706 , n40501 , n40502 );
nor ( n41707 , n9734 , n41439 );
and ( n41708 , n41706 , n41707 );
xor ( n41709 , n41706 , n41707 );
nor ( n41710 , n9752 , n40234 );
nor ( n41711 , n9743 , n41439 );
and ( n41712 , n41710 , n41711 );
and ( n41713 , n41709 , n41712 );
or ( n41714 , n41708 , n41713 );
and ( n41715 , n41705 , n41714 );
or ( n41716 , n41704 , n41715 );
and ( n41717 , n41701 , n41716 );
or ( n41718 , n41700 , n41717 );
and ( n41719 , n41697 , n41718 );
or ( n41720 , n41696 , n41719 );
and ( n41721 , n41693 , n41720 );
or ( n41722 , n41692 , n41721 );
and ( n41723 , n41689 , n41722 );
or ( n41724 , n41688 , n41723 );
and ( n41725 , n41685 , n41724 );
or ( n41726 , n41684 , n41725 );
and ( n41727 , n41681 , n41726 );
or ( n41728 , n41680 , n41727 );
and ( n41729 , n41677 , n41728 );
or ( n41730 , n41676 , n41729 );
and ( n41731 , n41673 , n41730 );
or ( n41732 , n41672 , n41731 );
and ( n41733 , n41669 , n41732 );
or ( n41734 , n41668 , n41733 );
and ( n41735 , n41665 , n41734 );
or ( n41736 , n41664 , n41735 );
and ( n41737 , n41661 , n41736 );
or ( n41738 , n41660 , n41737 );
and ( n41739 , n41657 , n41738 );
or ( n41740 , n41656 , n41739 );
and ( n41741 , n41653 , n41740 );
or ( n41742 , n41652 , n41741 );
and ( n41743 , n41649 , n41742 );
or ( n41744 , n41648 , n41743 );
and ( n41745 , n41645 , n41744 );
or ( n41746 , n41644 , n41745 );
and ( n41747 , n41641 , n41746 );
or ( n41748 , n41640 , n41747 );
and ( n41749 , n41637 , n41748 );
or ( n41750 , n41636 , n41749 );
and ( n41751 , n41633 , n41750 );
or ( n41752 , n41632 , n41751 );
and ( n41753 , n41629 , n41752 );
or ( n41754 , n41628 , n41753 );
and ( n41755 , n41625 , n41754 );
or ( n41756 , n41624 , n41755 );
and ( n41757 , n41621 , n41756 );
or ( n41758 , n41620 , n41757 );
and ( n41759 , n41617 , n41758 );
or ( n41760 , n41616 , n41759 );
and ( n41761 , n41613 , n41760 );
or ( n41762 , n41612 , n41761 );
and ( n41763 , n41609 , n41762 );
or ( n41764 , n41608 , n41763 );
and ( n41765 , n41605 , n41764 );
or ( n41766 , n41604 , n41765 );
and ( n41767 , n41601 , n41766 );
or ( n41768 , n41600 , n41767 );
and ( n41769 , n41597 , n41768 );
or ( n41770 , n41596 , n41769 );
and ( n41771 , n41593 , n41770 );
or ( n41772 , n41592 , n41771 );
and ( n41773 , n41589 , n41772 );
or ( n41774 , n41588 , n41773 );
and ( n41775 , n41585 , n41774 );
or ( n41776 , n41584 , n41775 );
and ( n41777 , n41581 , n41776 );
or ( n41778 , n41580 , n41777 );
and ( n41779 , n41577 , n41778 );
or ( n41780 , n41576 , n41779 );
and ( n41781 , n41573 , n41780 );
or ( n41782 , n41572 , n41781 );
and ( n41783 , n41569 , n41782 );
or ( n41784 , n41568 , n41783 );
and ( n41785 , n41565 , n41784 );
or ( n41786 , n41564 , n41785 );
and ( n41787 , n41561 , n41786 );
or ( n41788 , n41560 , n41787 );
and ( n41789 , n41557 , n41788 );
or ( n41790 , n41556 , n41789 );
and ( n41791 , n41553 , n41790 );
or ( n41792 , n41552 , n41791 );
and ( n41793 , n41549 , n41792 );
or ( n41794 , n41548 , n41793 );
and ( n41795 , n41545 , n41794 );
or ( n41796 , n41544 , n41795 );
and ( n41797 , n41541 , n41796 );
or ( n41798 , n41540 , n41797 );
and ( n41799 , n41537 , n41798 );
or ( n41800 , n41536 , n41799 );
and ( n41801 , n41533 , n41800 );
or ( n41802 , n41532 , n41801 );
and ( n41803 , n41529 , n41802 );
or ( n41804 , n41528 , n41803 );
and ( n41805 , n41525 , n41804 );
or ( n41806 , n41524 , n41805 );
and ( n41807 , n41521 , n41806 );
or ( n41808 , n41520 , n41807 );
and ( n41809 , n41517 , n41808 );
or ( n41810 , n41516 , n41809 );
and ( n41811 , n41513 , n41810 );
or ( n41812 , n41512 , n41811 );
and ( n41813 , n41509 , n41812 );
or ( n41814 , n41508 , n41813 );
and ( n41815 , n41505 , n41814 );
or ( n41816 , n41504 , n41815 );
and ( n41817 , n41501 , n41816 );
or ( n41818 , n41500 , n41817 );
and ( n41819 , n41497 , n41818 );
or ( n41820 , n41496 , n41819 );
and ( n41821 , n41493 , n41820 );
or ( n41822 , n41492 , n41821 );
and ( n41823 , n41489 , n41822 );
or ( n41824 , n41488 , n41823 );
and ( n41825 , n41485 , n41824 );
or ( n41826 , n41484 , n41825 );
and ( n41827 , n41481 , n41826 );
or ( n41828 , n41480 , n41827 );
and ( n41829 , n41477 , n41828 );
or ( n41830 , n41476 , n41829 );
and ( n41831 , n41473 , n41830 );
or ( n41832 , n41472 , n41831 );
and ( n41833 , n41469 , n41832 );
or ( n41834 , n41468 , n41833 );
and ( n41835 , n41465 , n41834 );
or ( n41836 , n41464 , n41835 );
and ( n41837 , n41461 , n41836 );
or ( n41838 , n41460 , n41837 );
and ( n41839 , n41457 , n41838 );
or ( n41840 , n41456 , n41839 );
and ( n41841 , n41453 , n41840 );
or ( n41842 , n41452 , n41841 );
and ( n41843 , n41449 , n41842 );
or ( n41844 , n41448 , n41843 );
and ( n41845 , n41445 , n41844 );
or ( n41846 , n41444 , n41845 );
xor ( n41847 , n41441 , n41846 );
and ( n41848 , n33403 , n867 );
nor ( n41849 , n868 , n41848 );
nor ( n41850 , n958 , n32231 );
xor ( n41851 , n41849 , n41850 );
and ( n41852 , n40638 , n40639 );
and ( n41853 , n40640 , n40643 );
or ( n41854 , n41852 , n41853 );
xor ( n41855 , n41851 , n41854 );
nor ( n41856 , n1062 , n31083 );
xor ( n41857 , n41855 , n41856 );
and ( n41858 , n40644 , n40645 );
and ( n41859 , n40646 , n40649 );
or ( n41860 , n41858 , n41859 );
xor ( n41861 , n41857 , n41860 );
nor ( n41862 , n1176 , n29948 );
xor ( n41863 , n41861 , n41862 );
and ( n41864 , n40650 , n40651 );
and ( n41865 , n40652 , n40655 );
or ( n41866 , n41864 , n41865 );
xor ( n41867 , n41863 , n41866 );
nor ( n41868 , n1303 , n28833 );
xor ( n41869 , n41867 , n41868 );
and ( n41870 , n40656 , n40657 );
and ( n41871 , n40658 , n40661 );
or ( n41872 , n41870 , n41871 );
xor ( n41873 , n41869 , n41872 );
nor ( n41874 , n1445 , n27737 );
xor ( n41875 , n41873 , n41874 );
and ( n41876 , n40662 , n40663 );
and ( n41877 , n40664 , n40667 );
or ( n41878 , n41876 , n41877 );
xor ( n41879 , n41875 , n41878 );
nor ( n41880 , n1598 , n26660 );
xor ( n41881 , n41879 , n41880 );
and ( n41882 , n40668 , n40669 );
and ( n41883 , n40670 , n40673 );
or ( n41884 , n41882 , n41883 );
xor ( n41885 , n41881 , n41884 );
nor ( n41886 , n1766 , n25600 );
xor ( n41887 , n41885 , n41886 );
and ( n41888 , n40674 , n40675 );
and ( n41889 , n40676 , n40679 );
or ( n41890 , n41888 , n41889 );
xor ( n41891 , n41887 , n41890 );
nor ( n41892 , n1945 , n24564 );
xor ( n41893 , n41891 , n41892 );
and ( n41894 , n40680 , n40681 );
and ( n41895 , n40682 , n40685 );
or ( n41896 , n41894 , n41895 );
xor ( n41897 , n41893 , n41896 );
nor ( n41898 , n2137 , n23541 );
xor ( n41899 , n41897 , n41898 );
and ( n41900 , n40686 , n40687 );
and ( n41901 , n40688 , n40691 );
or ( n41902 , n41900 , n41901 );
xor ( n41903 , n41899 , n41902 );
nor ( n41904 , n2343 , n22541 );
xor ( n41905 , n41903 , n41904 );
and ( n41906 , n40692 , n40693 );
and ( n41907 , n40694 , n40697 );
or ( n41908 , n41906 , n41907 );
xor ( n41909 , n41905 , n41908 );
nor ( n41910 , n2566 , n21562 );
xor ( n41911 , n41909 , n41910 );
and ( n41912 , n40698 , n40699 );
and ( n41913 , n40700 , n40703 );
or ( n41914 , n41912 , n41913 );
xor ( n41915 , n41911 , n41914 );
nor ( n41916 , n2797 , n20601 );
xor ( n41917 , n41915 , n41916 );
and ( n41918 , n40704 , n40705 );
and ( n41919 , n40706 , n40709 );
or ( n41920 , n41918 , n41919 );
xor ( n41921 , n41917 , n41920 );
nor ( n41922 , n3043 , n19657 );
xor ( n41923 , n41921 , n41922 );
and ( n41924 , n40710 , n40711 );
and ( n41925 , n40712 , n40715 );
or ( n41926 , n41924 , n41925 );
xor ( n41927 , n41923 , n41926 );
nor ( n41928 , n3300 , n18734 );
xor ( n41929 , n41927 , n41928 );
and ( n41930 , n40716 , n40717 );
and ( n41931 , n40718 , n40721 );
or ( n41932 , n41930 , n41931 );
xor ( n41933 , n41929 , n41932 );
nor ( n41934 , n3570 , n17828 );
xor ( n41935 , n41933 , n41934 );
and ( n41936 , n40722 , n40723 );
and ( n41937 , n40724 , n40727 );
or ( n41938 , n41936 , n41937 );
xor ( n41939 , n41935 , n41938 );
nor ( n41940 , n3853 , n16943 );
xor ( n41941 , n41939 , n41940 );
and ( n41942 , n40728 , n40729 );
and ( n41943 , n40730 , n40733 );
or ( n41944 , n41942 , n41943 );
xor ( n41945 , n41941 , n41944 );
nor ( n41946 , n4151 , n16077 );
xor ( n41947 , n41945 , n41946 );
and ( n41948 , n40734 , n40735 );
and ( n41949 , n40736 , n40739 );
or ( n41950 , n41948 , n41949 );
xor ( n41951 , n41947 , n41950 );
nor ( n41952 , n4458 , n15230 );
xor ( n41953 , n41951 , n41952 );
and ( n41954 , n40740 , n40741 );
and ( n41955 , n40742 , n40745 );
or ( n41956 , n41954 , n41955 );
xor ( n41957 , n41953 , n41956 );
nor ( n41958 , n4786 , n14403 );
xor ( n41959 , n41957 , n41958 );
and ( n41960 , n40746 , n40747 );
and ( n41961 , n40748 , n40751 );
or ( n41962 , n41960 , n41961 );
xor ( n41963 , n41959 , n41962 );
nor ( n41964 , n5126 , n13599 );
xor ( n41965 , n41963 , n41964 );
and ( n41966 , n40752 , n40753 );
and ( n41967 , n40754 , n40757 );
or ( n41968 , n41966 , n41967 );
xor ( n41969 , n41965 , n41968 );
nor ( n41970 , n5477 , n12808 );
xor ( n41971 , n41969 , n41970 );
and ( n41972 , n40758 , n40759 );
and ( n41973 , n40760 , n40763 );
or ( n41974 , n41972 , n41973 );
xor ( n41975 , n41971 , n41974 );
nor ( n41976 , n5838 , n12037 );
xor ( n41977 , n41975 , n41976 );
and ( n41978 , n40764 , n40765 );
and ( n41979 , n40766 , n40769 );
or ( n41980 , n41978 , n41979 );
xor ( n41981 , n41977 , n41980 );
nor ( n41982 , n6212 , n11282 );
xor ( n41983 , n41981 , n41982 );
and ( n41984 , n40770 , n40771 );
and ( n41985 , n40772 , n40775 );
or ( n41986 , n41984 , n41985 );
xor ( n41987 , n41983 , n41986 );
nor ( n41988 , n6596 , n10547 );
xor ( n41989 , n41987 , n41988 );
and ( n41990 , n40776 , n40777 );
and ( n41991 , n40778 , n40781 );
or ( n41992 , n41990 , n41991 );
xor ( n41993 , n41989 , n41992 );
nor ( n41994 , n6997 , n9829 );
xor ( n41995 , n41993 , n41994 );
and ( n41996 , n40782 , n40783 );
and ( n41997 , n40784 , n40787 );
or ( n41998 , n41996 , n41997 );
xor ( n41999 , n41995 , n41998 );
nor ( n42000 , n7413 , n8955 );
xor ( n42001 , n41999 , n42000 );
and ( n42002 , n40788 , n40789 );
and ( n42003 , n40790 , n40793 );
or ( n42004 , n42002 , n42003 );
xor ( n42005 , n42001 , n42004 );
nor ( n42006 , n7841 , n603 );
xor ( n42007 , n42005 , n42006 );
and ( n42008 , n40794 , n40795 );
and ( n42009 , n40796 , n40799 );
or ( n42010 , n42008 , n42009 );
xor ( n42011 , n42007 , n42010 );
nor ( n42012 , n8281 , n652 );
xor ( n42013 , n42011 , n42012 );
and ( n42014 , n40800 , n40801 );
and ( n42015 , n40802 , n40805 );
or ( n42016 , n42014 , n42015 );
xor ( n42017 , n42013 , n42016 );
nor ( n42018 , n8737 , n624 );
xor ( n42019 , n42017 , n42018 );
and ( n42020 , n40806 , n40807 );
and ( n42021 , n40808 , n40811 );
or ( n42022 , n42020 , n42021 );
xor ( n42023 , n42019 , n42022 );
nor ( n42024 , n9420 , n648 );
xor ( n42025 , n42023 , n42024 );
and ( n42026 , n40812 , n40813 );
and ( n42027 , n40814 , n40817 );
or ( n42028 , n42026 , n42027 );
xor ( n42029 , n42025 , n42028 );
nor ( n42030 , n10312 , n686 );
xor ( n42031 , n42029 , n42030 );
and ( n42032 , n40818 , n40819 );
and ( n42033 , n40820 , n40823 );
or ( n42034 , n42032 , n42033 );
xor ( n42035 , n42031 , n42034 );
nor ( n42036 , n11041 , n735 );
xor ( n42037 , n42035 , n42036 );
and ( n42038 , n40824 , n40825 );
and ( n42039 , n40826 , n40829 );
or ( n42040 , n42038 , n42039 );
xor ( n42041 , n42037 , n42040 );
nor ( n42042 , n11790 , n798 );
xor ( n42043 , n42041 , n42042 );
and ( n42044 , n40830 , n40831 );
and ( n42045 , n40832 , n40835 );
or ( n42046 , n42044 , n42045 );
xor ( n42047 , n42043 , n42046 );
nor ( n42048 , n12555 , n870 );
xor ( n42049 , n42047 , n42048 );
and ( n42050 , n40836 , n40837 );
and ( n42051 , n40838 , n40841 );
or ( n42052 , n42050 , n42051 );
xor ( n42053 , n42049 , n42052 );
nor ( n42054 , n13340 , n960 );
xor ( n42055 , n42053 , n42054 );
and ( n42056 , n40842 , n40843 );
and ( n42057 , n40844 , n40847 );
or ( n42058 , n42056 , n42057 );
xor ( n42059 , n42055 , n42058 );
nor ( n42060 , n14138 , n1064 );
xor ( n42061 , n42059 , n42060 );
and ( n42062 , n40848 , n40849 );
and ( n42063 , n40850 , n40853 );
or ( n42064 , n42062 , n42063 );
xor ( n42065 , n42061 , n42064 );
nor ( n42066 , n14959 , n1178 );
xor ( n42067 , n42065 , n42066 );
and ( n42068 , n40854 , n40855 );
and ( n42069 , n40856 , n40859 );
or ( n42070 , n42068 , n42069 );
xor ( n42071 , n42067 , n42070 );
nor ( n42072 , n15800 , n1305 );
xor ( n42073 , n42071 , n42072 );
and ( n42074 , n40860 , n40861 );
and ( n42075 , n40862 , n40865 );
or ( n42076 , n42074 , n42075 );
xor ( n42077 , n42073 , n42076 );
nor ( n42078 , n16660 , n1447 );
xor ( n42079 , n42077 , n42078 );
and ( n42080 , n40866 , n40867 );
and ( n42081 , n40868 , n40871 );
or ( n42082 , n42080 , n42081 );
xor ( n42083 , n42079 , n42082 );
nor ( n42084 , n17539 , n1600 );
xor ( n42085 , n42083 , n42084 );
and ( n42086 , n40872 , n40873 );
and ( n42087 , n40874 , n40877 );
or ( n42088 , n42086 , n42087 );
xor ( n42089 , n42085 , n42088 );
nor ( n42090 , n18439 , n1768 );
xor ( n42091 , n42089 , n42090 );
and ( n42092 , n40878 , n40879 );
and ( n42093 , n40880 , n40883 );
or ( n42094 , n42092 , n42093 );
xor ( n42095 , n42091 , n42094 );
nor ( n42096 , n19356 , n1947 );
xor ( n42097 , n42095 , n42096 );
and ( n42098 , n40884 , n40885 );
and ( n42099 , n40886 , n40889 );
or ( n42100 , n42098 , n42099 );
xor ( n42101 , n42097 , n42100 );
nor ( n42102 , n20294 , n2139 );
xor ( n42103 , n42101 , n42102 );
and ( n42104 , n40890 , n40891 );
and ( n42105 , n40892 , n40895 );
or ( n42106 , n42104 , n42105 );
xor ( n42107 , n42103 , n42106 );
nor ( n42108 , n21249 , n2345 );
xor ( n42109 , n42107 , n42108 );
and ( n42110 , n40896 , n40897 );
and ( n42111 , n40898 , n40901 );
or ( n42112 , n42110 , n42111 );
xor ( n42113 , n42109 , n42112 );
nor ( n42114 , n22222 , n2568 );
xor ( n42115 , n42113 , n42114 );
and ( n42116 , n40902 , n40903 );
and ( n42117 , n40904 , n40907 );
or ( n42118 , n42116 , n42117 );
xor ( n42119 , n42115 , n42118 );
nor ( n42120 , n23216 , n2799 );
xor ( n42121 , n42119 , n42120 );
and ( n42122 , n40908 , n40909 );
and ( n42123 , n40910 , n40913 );
or ( n42124 , n42122 , n42123 );
xor ( n42125 , n42121 , n42124 );
nor ( n42126 , n24233 , n3045 );
xor ( n42127 , n42125 , n42126 );
and ( n42128 , n40914 , n40915 );
and ( n42129 , n40916 , n40919 );
or ( n42130 , n42128 , n42129 );
xor ( n42131 , n42127 , n42130 );
nor ( n42132 , n25263 , n3302 );
xor ( n42133 , n42131 , n42132 );
and ( n42134 , n40920 , n40921 );
and ( n42135 , n40922 , n40925 );
or ( n42136 , n42134 , n42135 );
xor ( n42137 , n42133 , n42136 );
nor ( n42138 , n26317 , n3572 );
xor ( n42139 , n42137 , n42138 );
and ( n42140 , n40926 , n40927 );
and ( n42141 , n40928 , n40931 );
or ( n42142 , n42140 , n42141 );
xor ( n42143 , n42139 , n42142 );
nor ( n42144 , n27388 , n3855 );
xor ( n42145 , n42143 , n42144 );
and ( n42146 , n40932 , n40933 );
and ( n42147 , n40934 , n40937 );
or ( n42148 , n42146 , n42147 );
xor ( n42149 , n42145 , n42148 );
nor ( n42150 , n28478 , n4153 );
xor ( n42151 , n42149 , n42150 );
and ( n42152 , n40938 , n40939 );
and ( n42153 , n40940 , n40943 );
or ( n42154 , n42152 , n42153 );
xor ( n42155 , n42151 , n42154 );
nor ( n42156 , n29587 , n4460 );
xor ( n42157 , n42155 , n42156 );
and ( n42158 , n40944 , n40945 );
and ( n42159 , n40946 , n40949 );
or ( n42160 , n42158 , n42159 );
xor ( n42161 , n42157 , n42160 );
nor ( n42162 , n30716 , n4788 );
xor ( n42163 , n42161 , n42162 );
and ( n42164 , n40950 , n40951 );
and ( n42165 , n40952 , n40955 );
or ( n42166 , n42164 , n42165 );
xor ( n42167 , n42163 , n42166 );
nor ( n42168 , n31858 , n5128 );
xor ( n42169 , n42167 , n42168 );
and ( n42170 , n40956 , n40957 );
and ( n42171 , n40958 , n40961 );
or ( n42172 , n42170 , n42171 );
xor ( n42173 , n42169 , n42172 );
nor ( n42174 , n33024 , n5479 );
xor ( n42175 , n42173 , n42174 );
and ( n42176 , n40962 , n40963 );
and ( n42177 , n40964 , n40967 );
or ( n42178 , n42176 , n42177 );
xor ( n42179 , n42175 , n42178 );
nor ( n42180 , n34215 , n5840 );
xor ( n42181 , n42179 , n42180 );
and ( n42182 , n40968 , n40969 );
and ( n42183 , n40970 , n40973 );
or ( n42184 , n42182 , n42183 );
xor ( n42185 , n42181 , n42184 );
nor ( n42186 , n35410 , n6214 );
xor ( n42187 , n42185 , n42186 );
and ( n42188 , n40974 , n40975 );
and ( n42189 , n40976 , n40979 );
or ( n42190 , n42188 , n42189 );
xor ( n42191 , n42187 , n42190 );
nor ( n42192 , n36611 , n6598 );
xor ( n42193 , n42191 , n42192 );
and ( n42194 , n40980 , n40981 );
and ( n42195 , n40982 , n40985 );
or ( n42196 , n42194 , n42195 );
xor ( n42197 , n42193 , n42196 );
nor ( n42198 , n37816 , n6999 );
xor ( n42199 , n42197 , n42198 );
and ( n42200 , n40986 , n40987 );
and ( n42201 , n40988 , n40991 );
or ( n42202 , n42200 , n42201 );
xor ( n42203 , n42199 , n42202 );
nor ( n42204 , n39018 , n7415 );
xor ( n42205 , n42203 , n42204 );
and ( n42206 , n40992 , n40993 );
and ( n42207 , n40994 , n40997 );
or ( n42208 , n42206 , n42207 );
xor ( n42209 , n42205 , n42208 );
nor ( n42210 , n40223 , n7843 );
xor ( n42211 , n42209 , n42210 );
and ( n42212 , n40998 , n40999 );
and ( n42213 , n41000 , n41003 );
or ( n42214 , n42212 , n42213 );
xor ( n42215 , n42211 , n42214 );
nor ( n42216 , n41428 , n8283 );
xor ( n42217 , n42215 , n42216 );
and ( n42218 , n41004 , n41005 );
and ( n42219 , n41006 , n41009 );
or ( n42220 , n42218 , n42219 );
xor ( n42221 , n42217 , n42220 );
and ( n42222 , n41022 , n41026 );
and ( n42223 , n41026 , n41414 );
and ( n42224 , n41022 , n41414 );
or ( n42225 , n42222 , n42223 , n42224 );
and ( n42226 , n33774 , n840 );
not ( n42227 , n840 );
nor ( n42228 , n42226 , n42227 );
xor ( n42229 , n42225 , n42228 );
and ( n42230 , n41035 , n41039 );
and ( n42231 , n41039 , n41107 );
and ( n42232 , n41035 , n41107 );
or ( n42233 , n42230 , n42231 , n42232 );
and ( n42234 , n41031 , n41108 );
and ( n42235 , n41108 , n41413 );
and ( n42236 , n41031 , n41413 );
or ( n42237 , n42234 , n42235 , n42236 );
xor ( n42238 , n42233 , n42237 );
and ( n42239 , n41113 , n41233 );
and ( n42240 , n41233 , n41412 );
and ( n42241 , n41113 , n41412 );
or ( n42242 , n42239 , n42240 , n42241 );
and ( n42243 , n41044 , n41048 );
and ( n42244 , n41048 , n41106 );
and ( n42245 , n41044 , n41106 );
or ( n42246 , n42243 , n42244 , n42245 );
and ( n42247 , n41117 , n41121 );
and ( n42248 , n41121 , n41232 );
and ( n42249 , n41117 , n41232 );
or ( n42250 , n42247 , n42248 , n42249 );
xor ( n42251 , n42246 , n42250 );
and ( n42252 , n41075 , n41079 );
and ( n42253 , n41079 , n41085 );
and ( n42254 , n41075 , n41085 );
or ( n42255 , n42252 , n42253 , n42254 );
and ( n42256 , n41053 , n41057 );
and ( n42257 , n41057 , n41105 );
and ( n42258 , n41053 , n41105 );
or ( n42259 , n42256 , n42257 , n42258 );
xor ( n42260 , n42255 , n42259 );
and ( n42261 , n41062 , n41066 );
and ( n42262 , n41066 , n41104 );
and ( n42263 , n41062 , n41104 );
or ( n42264 , n42261 , n42262 , n42263 );
and ( n42265 , n41130 , n41155 );
and ( n42266 , n41155 , n41193 );
and ( n42267 , n41130 , n41193 );
or ( n42268 , n42265 , n42266 , n42267 );
xor ( n42269 , n42264 , n42268 );
and ( n42270 , n41071 , n41086 );
and ( n42271 , n41086 , n41103 );
and ( n42272 , n41071 , n41103 );
or ( n42273 , n42270 , n42271 , n42272 );
and ( n42274 , n41134 , n41138 );
and ( n42275 , n41138 , n41154 );
and ( n42276 , n41134 , n41154 );
or ( n42277 , n42274 , n42275 , n42276 );
xor ( n42278 , n42273 , n42277 );
and ( n42279 , n41091 , n41096 );
and ( n42280 , n41096 , n41102 );
and ( n42281 , n41091 , n41102 );
or ( n42282 , n42279 , n42280 , n42281 );
and ( n42283 , n41081 , n41082 );
and ( n42284 , n41082 , n41084 );
and ( n42285 , n41081 , n41084 );
or ( n42286 , n42283 , n42284 , n42285 );
and ( n42287 , n41092 , n41093 );
and ( n42288 , n41093 , n41095 );
and ( n42289 , n41092 , n41095 );
or ( n42290 , n42287 , n42288 , n42289 );
xor ( n42291 , n42286 , n42290 );
and ( n42292 , n30695 , n1134 );
and ( n42293 , n31836 , n1034 );
xor ( n42294 , n42292 , n42293 );
and ( n42295 , n32649 , n940 );
xor ( n42296 , n42294 , n42295 );
xor ( n42297 , n42291 , n42296 );
xor ( n42298 , n42282 , n42297 );
and ( n42299 , n41098 , n41099 );
and ( n42300 , n41099 , n41101 );
and ( n42301 , n41098 , n41101 );
or ( n42302 , n42299 , n42300 , n42301 );
and ( n42303 , n27361 , n1551 );
and ( n42304 , n28456 , n1424 );
xor ( n42305 , n42303 , n42304 );
and ( n42306 , n29559 , n1254 );
xor ( n42307 , n42305 , n42306 );
xor ( n42308 , n42302 , n42307 );
and ( n42309 , n24214 , n2100 );
and ( n42310 , n25243 , n1882 );
xor ( n42311 , n42309 , n42310 );
and ( n42312 , n26296 , n1738 );
xor ( n42313 , n42311 , n42312 );
xor ( n42314 , n42308 , n42313 );
xor ( n42315 , n42298 , n42314 );
xor ( n42316 , n42278 , n42315 );
xor ( n42317 , n42269 , n42316 );
xor ( n42318 , n42260 , n42317 );
xor ( n42319 , n42251 , n42318 );
xor ( n42320 , n42242 , n42319 );
and ( n42321 , n41238 , n41316 );
and ( n42322 , n41316 , n41411 );
and ( n42323 , n41238 , n41411 );
or ( n42324 , n42321 , n42322 , n42323 );
and ( n42325 , n41126 , n41194 );
and ( n42326 , n41194 , n41231 );
and ( n42327 , n41126 , n41231 );
or ( n42328 , n42325 , n42326 , n42327 );
and ( n42329 , n41242 , n41246 );
and ( n42330 , n41246 , n41315 );
and ( n42331 , n41242 , n41315 );
or ( n42332 , n42329 , n42330 , n42331 );
xor ( n42333 , n42328 , n42332 );
and ( n42334 , n41199 , n41203 );
and ( n42335 , n41203 , n41230 );
and ( n42336 , n41199 , n41230 );
or ( n42337 , n42334 , n42335 , n42336 );
and ( n42338 , n41160 , n41176 );
and ( n42339 , n41176 , n41192 );
and ( n42340 , n41160 , n41192 );
or ( n42341 , n42338 , n42339 , n42340 );
and ( n42342 , n41143 , n41147 );
and ( n42343 , n41147 , n41153 );
and ( n42344 , n41143 , n41153 );
or ( n42345 , n42342 , n42343 , n42344 );
and ( n42346 , n41164 , n41169 );
and ( n42347 , n41169 , n41175 );
and ( n42348 , n41164 , n41175 );
or ( n42349 , n42346 , n42347 , n42348 );
xor ( n42350 , n42345 , n42349 );
and ( n42351 , n41149 , n41150 );
and ( n42352 , n41150 , n41152 );
and ( n42353 , n41149 , n41152 );
or ( n42354 , n42351 , n42352 , n42353 );
and ( n42355 , n41165 , n41166 );
and ( n42356 , n41166 , n41168 );
and ( n42357 , n41165 , n41168 );
or ( n42358 , n42355 , n42356 , n42357 );
xor ( n42359 , n42354 , n42358 );
and ( n42360 , n21216 , n2739 );
and ( n42361 , n22186 , n2544 );
xor ( n42362 , n42360 , n42361 );
and ( n42363 , n22892 , n2298 );
xor ( n42364 , n42362 , n42363 );
xor ( n42365 , n42359 , n42364 );
xor ( n42366 , n42350 , n42365 );
xor ( n42367 , n42341 , n42366 );
and ( n42368 , n41181 , n41185 );
and ( n42369 , n41185 , n41191 );
and ( n42370 , n41181 , n41191 );
or ( n42371 , n42368 , n42369 , n42370 );
and ( n42372 , n41171 , n41172 );
and ( n42373 , n41172 , n41174 );
and ( n42374 , n41171 , n41174 );
or ( n42375 , n42372 , n42373 , n42374 );
and ( n42376 , n18144 , n3495 );
and ( n42377 , n19324 , n3271 );
xor ( n42378 , n42376 , n42377 );
and ( n42379 , n20233 , n2981 );
xor ( n42380 , n42378 , n42379 );
xor ( n42381 , n42375 , n42380 );
and ( n42382 , n15758 , n4403 );
and ( n42383 , n16637 , n4102 );
xor ( n42384 , n42382 , n42383 );
and ( n42385 , n17512 , n3749 );
xor ( n42386 , n42384 , n42385 );
xor ( n42387 , n42381 , n42386 );
xor ( n42388 , n42371 , n42387 );
and ( n42389 , n41187 , n41188 );
and ( n42390 , n41188 , n41190 );
and ( n42391 , n41187 , n41190 );
or ( n42392 , n42389 , n42390 , n42391 );
and ( n42393 , n41218 , n41219 );
and ( n42394 , n41219 , n41221 );
and ( n42395 , n41218 , n41221 );
or ( n42396 , n42393 , n42394 , n42395 );
xor ( n42397 , n42392 , n42396 );
and ( n42398 , n13322 , n5408 );
and ( n42399 , n14118 , n5103 );
xor ( n42400 , n42398 , n42399 );
and ( n42401 , n14938 , n4730 );
xor ( n42402 , n42400 , n42401 );
xor ( n42403 , n42397 , n42402 );
xor ( n42404 , n42388 , n42403 );
xor ( n42405 , n42367 , n42404 );
xor ( n42406 , n42337 , n42405 );
and ( n42407 , n41208 , n41212 );
and ( n42408 , n41212 , n41229 );
and ( n42409 , n41208 , n41229 );
or ( n42410 , n42407 , n42408 , n42409 );
and ( n42411 , n41255 , n41270 );
and ( n42412 , n41270 , n41287 );
and ( n42413 , n41255 , n41287 );
or ( n42414 , n42411 , n42412 , n42413 );
xor ( n42415 , n42410 , n42414 );
and ( n42416 , n41217 , n41222 );
and ( n42417 , n41222 , n41228 );
and ( n42418 , n41217 , n41228 );
or ( n42419 , n42416 , n42417 , n42418 );
and ( n42420 , n41259 , n41263 );
and ( n42421 , n41263 , n41269 );
and ( n42422 , n41259 , n41269 );
or ( n42423 , n42420 , n42421 , n42422 );
xor ( n42424 , n42419 , n42423 );
and ( n42425 , n41224 , n41225 );
and ( n42426 , n41225 , n41227 );
and ( n42427 , n41224 , n41227 );
or ( n42428 , n42425 , n42426 , n42427 );
and ( n42429 , n11015 , n6504 );
and ( n42430 , n11769 , n6132 );
xor ( n42431 , n42429 , n42430 );
and ( n42432 , n12320 , n5765 );
xor ( n42433 , n42431 , n42432 );
xor ( n42434 , n42428 , n42433 );
and ( n42435 , n8718 , n7662 );
and ( n42436 , n9400 , n7310 );
xor ( n42437 , n42435 , n42436 );
and ( n42438 , n10291 , n6971 );
xor ( n42439 , n42437 , n42438 );
xor ( n42440 , n42434 , n42439 );
xor ( n42441 , n42424 , n42440 );
xor ( n42442 , n42415 , n42441 );
xor ( n42443 , n42406 , n42442 );
xor ( n42444 , n42333 , n42443 );
xor ( n42445 , n42324 , n42444 );
and ( n42446 , n41321 , n41368 );
and ( n42447 , n41368 , n41410 );
and ( n42448 , n41321 , n41410 );
or ( n42449 , n42446 , n42447 , n42448 );
and ( n42450 , n41251 , n41288 );
and ( n42451 , n41288 , n41314 );
and ( n42452 , n41251 , n41314 );
or ( n42453 , n42450 , n42451 , n42452 );
and ( n42454 , n41325 , n41329 );
and ( n42455 , n41329 , n41367 );
and ( n42456 , n41325 , n41367 );
or ( n42457 , n42454 , n42455 , n42456 );
xor ( n42458 , n42453 , n42457 );
and ( n42459 , n41293 , n41297 );
and ( n42460 , n41297 , n41313 );
and ( n42461 , n41293 , n41313 );
or ( n42462 , n42459 , n42460 , n42461 );
and ( n42463 , n41275 , n41280 );
and ( n42464 , n41280 , n41286 );
and ( n42465 , n41275 , n41286 );
or ( n42466 , n42463 , n42464 , n42465 );
and ( n42467 , n41265 , n41266 );
and ( n42468 , n41266 , n41268 );
and ( n42469 , n41265 , n41268 );
or ( n42470 , n42467 , n42468 , n42469 );
and ( n42471 , n41276 , n41277 );
and ( n42472 , n41277 , n41279 );
and ( n42473 , n41276 , n41279 );
or ( n42474 , n42471 , n42472 , n42473 );
xor ( n42475 , n42470 , n42474 );
and ( n42476 , n7385 , n9348 );
and ( n42477 , n7808 , n8669 );
xor ( n42478 , n42476 , n42477 );
buf ( n42479 , n8079 );
xor ( n42480 , n42478 , n42479 );
xor ( n42481 , n42475 , n42480 );
xor ( n42482 , n42466 , n42481 );
and ( n42483 , n41282 , n41283 );
and ( n42484 , n41283 , n41285 );
and ( n42485 , n41282 , n41285 );
or ( n42486 , n42483 , n42484 , n42485 );
and ( n42487 , n6187 , n11718 );
and ( n42488 , n6569 , n10977 );
xor ( n42489 , n42487 , n42488 );
and ( n42490 , n6816 , n10239 );
xor ( n42491 , n42489 , n42490 );
xor ( n42492 , n42486 , n42491 );
and ( n42493 , n4959 , n14044 );
and ( n42494 , n5459 , n13256 );
xor ( n42495 , n42493 , n42494 );
and ( n42496 , n5819 , n12531 );
xor ( n42497 , n42495 , n42496 );
xor ( n42498 , n42492 , n42497 );
xor ( n42499 , n42482 , n42498 );
xor ( n42500 , n42462 , n42499 );
and ( n42501 , n41302 , n41306 );
and ( n42502 , n41306 , n41312 );
and ( n42503 , n41302 , n41312 );
or ( n42504 , n42501 , n42502 , n42503 );
and ( n42505 , n41338 , n41343 );
and ( n42506 , n41343 , n41349 );
and ( n42507 , n41338 , n41349 );
or ( n42508 , n42505 , n42506 , n42507 );
xor ( n42509 , n42504 , n42508 );
and ( n42510 , n41308 , n41309 );
and ( n42511 , n41309 , n41311 );
and ( n42512 , n41308 , n41311 );
or ( n42513 , n42510 , n42511 , n42512 );
and ( n42514 , n41339 , n41340 );
and ( n42515 , n41340 , n41342 );
and ( n42516 , n41339 , n41342 );
or ( n42517 , n42514 , n42515 , n42516 );
xor ( n42518 , n42513 , n42517 );
and ( n42519 , n4132 , n16550 );
and ( n42520 , n4438 , n15691 );
xor ( n42521 , n42519 , n42520 );
and ( n42522 , n4766 , n14838 );
xor ( n42523 , n42521 , n42522 );
xor ( n42524 , n42518 , n42523 );
xor ( n42525 , n42509 , n42524 );
xor ( n42526 , n42500 , n42525 );
xor ( n42527 , n42458 , n42526 );
xor ( n42528 , n42449 , n42527 );
and ( n42529 , n41370 , n41396 );
and ( n42530 , n41396 , n41409 );
and ( n42531 , n41370 , n41409 );
or ( n42532 , n42529 , n42530 , n42531 );
and ( n42533 , n41334 , n41350 );
and ( n42534 , n41350 , n41366 );
and ( n42535 , n41334 , n41366 );
or ( n42536 , n42533 , n42534 , n42535 );
and ( n42537 , n41374 , n41378 );
and ( n42538 , n41378 , n41395 );
and ( n42539 , n41374 , n41395 );
or ( n42540 , n42537 , n42538 , n42539 );
xor ( n42541 , n42536 , n42540 );
and ( n42542 , n41355 , n41359 );
and ( n42543 , n41359 , n41365 );
and ( n42544 , n41355 , n41365 );
or ( n42545 , n42542 , n42543 , n42544 );
and ( n42546 , n41345 , n41346 );
and ( n42547 , n41346 , n41348 );
and ( n42548 , n41345 , n41348 );
or ( n42549 , n42546 , n42547 , n42548 );
and ( n42550 , n3182 , n19222 );
and ( n42551 , n3545 , n18407 );
xor ( n42552 , n42550 , n42551 );
and ( n42553 , n3801 , n17422 );
xor ( n42554 , n42552 , n42553 );
xor ( n42555 , n42549 , n42554 );
and ( n42556 , n2462 , n22065 );
and ( n42557 , n2779 , n20976 );
xor ( n42558 , n42556 , n42557 );
and ( n42559 , n3024 , n20156 );
xor ( n42560 , n42558 , n42559 );
xor ( n42561 , n42555 , n42560 );
xor ( n42562 , n42545 , n42561 );
and ( n42563 , n41361 , n41362 );
and ( n42564 , n41362 , n41364 );
and ( n42565 , n41361 , n41364 );
or ( n42566 , n42563 , n42564 , n42565 );
and ( n42567 , n41384 , n41385 );
and ( n42568 , n41385 , n41387 );
and ( n42569 , n41384 , n41387 );
or ( n42570 , n42567 , n42568 , n42569 );
xor ( n42571 , n42566 , n42570 );
and ( n42572 , n1933 , n25163 );
and ( n42573 , n2120 , n24137 );
xor ( n42574 , n42572 , n42573 );
and ( n42575 , n2324 , n23075 );
xor ( n42576 , n42574 , n42575 );
xor ( n42577 , n42571 , n42576 );
xor ( n42578 , n42562 , n42577 );
xor ( n42579 , n42541 , n42578 );
xor ( n42580 , n42532 , n42579 );
and ( n42581 , n41383 , n41388 );
and ( n42582 , n41388 , n41394 );
and ( n42583 , n41383 , n41394 );
or ( n42584 , n42581 , n42582 , n42583 );
and ( n42585 , n41401 , n41408 );
xor ( n42586 , n42584 , n42585 );
and ( n42587 , n41390 , n41391 );
and ( n42588 , n41391 , n41393 );
and ( n42589 , n41390 , n41393 );
or ( n42590 , n42587 , n42588 , n42589 );
and ( n42591 , n1047 , n31761 );
and ( n42592 , n1164 , n30629 );
xor ( n42593 , n42591 , n42592 );
and ( n42594 , n1287 , n29508 );
xor ( n42595 , n42593 , n42594 );
xor ( n42596 , n42590 , n42595 );
and ( n42597 , n1383 , n28406 );
and ( n42598 , n1580 , n27296 );
xor ( n42599 , n42597 , n42598 );
and ( n42600 , n1694 , n26216 );
xor ( n42601 , n42599 , n42600 );
xor ( n42602 , n42596 , n42601 );
xor ( n42603 , n42586 , n42602 );
and ( n42604 , n41404 , n41405 );
and ( n42605 , n41405 , n41407 );
and ( n42606 , n41404 , n41407 );
or ( n42607 , n42604 , n42605 , n42606 );
not ( n42608 , n856 );
and ( n42609 , n34193 , n856 );
nor ( n42610 , n42608 , n42609 );
and ( n42611 , n925 , n32999 );
xor ( n42612 , n42610 , n42611 );
xor ( n42613 , n42607 , n42612 );
xor ( n42614 , n42603 , n42613 );
xor ( n42615 , n42580 , n42614 );
xor ( n42616 , n42528 , n42615 );
xor ( n42617 , n42445 , n42616 );
xor ( n42618 , n42320 , n42617 );
xor ( n42619 , n42238 , n42618 );
xor ( n42620 , n42229 , n42619 );
and ( n42621 , n41014 , n41017 );
and ( n42622 , n41017 , n41415 );
and ( n42623 , n41014 , n41415 );
or ( n42624 , n42621 , n42622 , n42623 );
xor ( n42625 , n42620 , n42624 );
and ( n42626 , n41416 , n41420 );
and ( n42627 , n41421 , n41424 );
or ( n42628 , n42626 , n42627 );
xor ( n42629 , n42625 , n42628 );
buf ( n42630 , n42629 );
buf ( n42631 , n42630 );
not ( n42632 , n42631 );
nor ( n42633 , n42632 , n8739 );
xor ( n42634 , n42221 , n42633 );
and ( n42635 , n41010 , n41429 );
and ( n42636 , n41430 , n41433 );
or ( n42637 , n42635 , n42636 );
xor ( n42638 , n42634 , n42637 );
buf ( n42639 , n42638 );
buf ( n42640 , n42639 );
not ( n42641 , n42640 );
buf ( n42642 , n569 );
not ( n42643 , n42642 );
nor ( n42644 , n42641 , n42643 );
xor ( n42645 , n41847 , n42644 );
xor ( n42646 , n41445 , n41844 );
nor ( n42647 , n41437 , n42643 );
and ( n42648 , n42646 , n42647 );
xor ( n42649 , n42646 , n42647 );
xor ( n42650 , n41449 , n41842 );
nor ( n42651 , n40232 , n42643 );
and ( n42652 , n42650 , n42651 );
xor ( n42653 , n42650 , n42651 );
xor ( n42654 , n41453 , n41840 );
nor ( n42655 , n39027 , n42643 );
and ( n42656 , n42654 , n42655 );
xor ( n42657 , n42654 , n42655 );
xor ( n42658 , n41457 , n41838 );
nor ( n42659 , n37825 , n42643 );
and ( n42660 , n42658 , n42659 );
xor ( n42661 , n42658 , n42659 );
xor ( n42662 , n41461 , n41836 );
nor ( n42663 , n36620 , n42643 );
and ( n42664 , n42662 , n42663 );
xor ( n42665 , n42662 , n42663 );
xor ( n42666 , n41465 , n41834 );
nor ( n42667 , n35419 , n42643 );
and ( n42668 , n42666 , n42667 );
xor ( n42669 , n42666 , n42667 );
xor ( n42670 , n41469 , n41832 );
nor ( n42671 , n34224 , n42643 );
and ( n42672 , n42670 , n42671 );
xor ( n42673 , n42670 , n42671 );
xor ( n42674 , n41473 , n41830 );
nor ( n42675 , n33033 , n42643 );
and ( n42676 , n42674 , n42675 );
xor ( n42677 , n42674 , n42675 );
xor ( n42678 , n41477 , n41828 );
nor ( n42679 , n31867 , n42643 );
and ( n42680 , n42678 , n42679 );
xor ( n42681 , n42678 , n42679 );
xor ( n42682 , n41481 , n41826 );
nor ( n42683 , n30725 , n42643 );
and ( n42684 , n42682 , n42683 );
xor ( n42685 , n42682 , n42683 );
xor ( n42686 , n41485 , n41824 );
nor ( n42687 , n29596 , n42643 );
and ( n42688 , n42686 , n42687 );
xor ( n42689 , n42686 , n42687 );
xor ( n42690 , n41489 , n41822 );
nor ( n42691 , n28487 , n42643 );
and ( n42692 , n42690 , n42691 );
xor ( n42693 , n42690 , n42691 );
xor ( n42694 , n41493 , n41820 );
nor ( n42695 , n27397 , n42643 );
and ( n42696 , n42694 , n42695 );
xor ( n42697 , n42694 , n42695 );
xor ( n42698 , n41497 , n41818 );
nor ( n42699 , n26326 , n42643 );
and ( n42700 , n42698 , n42699 );
xor ( n42701 , n42698 , n42699 );
xor ( n42702 , n41501 , n41816 );
nor ( n42703 , n25272 , n42643 );
and ( n42704 , n42702 , n42703 );
xor ( n42705 , n42702 , n42703 );
xor ( n42706 , n41505 , n41814 );
nor ( n42707 , n24242 , n42643 );
and ( n42708 , n42706 , n42707 );
xor ( n42709 , n42706 , n42707 );
xor ( n42710 , n41509 , n41812 );
nor ( n42711 , n23225 , n42643 );
and ( n42712 , n42710 , n42711 );
xor ( n42713 , n42710 , n42711 );
xor ( n42714 , n41513 , n41810 );
nor ( n42715 , n22231 , n42643 );
and ( n42716 , n42714 , n42715 );
xor ( n42717 , n42714 , n42715 );
xor ( n42718 , n41517 , n41808 );
nor ( n42719 , n21258 , n42643 );
and ( n42720 , n42718 , n42719 );
xor ( n42721 , n42718 , n42719 );
xor ( n42722 , n41521 , n41806 );
nor ( n42723 , n20303 , n42643 );
and ( n42724 , n42722 , n42723 );
xor ( n42725 , n42722 , n42723 );
xor ( n42726 , n41525 , n41804 );
nor ( n42727 , n19365 , n42643 );
and ( n42728 , n42726 , n42727 );
xor ( n42729 , n42726 , n42727 );
xor ( n42730 , n41529 , n41802 );
nor ( n42731 , n18448 , n42643 );
and ( n42732 , n42730 , n42731 );
xor ( n42733 , n42730 , n42731 );
xor ( n42734 , n41533 , n41800 );
nor ( n42735 , n17548 , n42643 );
and ( n42736 , n42734 , n42735 );
xor ( n42737 , n42734 , n42735 );
xor ( n42738 , n41537 , n41798 );
nor ( n42739 , n16669 , n42643 );
and ( n42740 , n42738 , n42739 );
xor ( n42741 , n42738 , n42739 );
xor ( n42742 , n41541 , n41796 );
nor ( n42743 , n15809 , n42643 );
and ( n42744 , n42742 , n42743 );
xor ( n42745 , n42742 , n42743 );
xor ( n42746 , n41545 , n41794 );
nor ( n42747 , n14968 , n42643 );
and ( n42748 , n42746 , n42747 );
xor ( n42749 , n42746 , n42747 );
xor ( n42750 , n41549 , n41792 );
nor ( n42751 , n14147 , n42643 );
and ( n42752 , n42750 , n42751 );
xor ( n42753 , n42750 , n42751 );
xor ( n42754 , n41553 , n41790 );
nor ( n42755 , n13349 , n42643 );
and ( n42756 , n42754 , n42755 );
xor ( n42757 , n42754 , n42755 );
xor ( n42758 , n41557 , n41788 );
nor ( n42759 , n12564 , n42643 );
and ( n42760 , n42758 , n42759 );
xor ( n42761 , n42758 , n42759 );
xor ( n42762 , n41561 , n41786 );
nor ( n42763 , n11799 , n42643 );
and ( n42764 , n42762 , n42763 );
xor ( n42765 , n42762 , n42763 );
xor ( n42766 , n41565 , n41784 );
nor ( n42767 , n11050 , n42643 );
and ( n42768 , n42766 , n42767 );
xor ( n42769 , n42766 , n42767 );
xor ( n42770 , n41569 , n41782 );
nor ( n42771 , n10321 , n42643 );
and ( n42772 , n42770 , n42771 );
xor ( n42773 , n42770 , n42771 );
xor ( n42774 , n41573 , n41780 );
nor ( n42775 , n9429 , n42643 );
and ( n42776 , n42774 , n42775 );
xor ( n42777 , n42774 , n42775 );
xor ( n42778 , n41577 , n41778 );
nor ( n42779 , n8949 , n42643 );
and ( n42780 , n42778 , n42779 );
xor ( n42781 , n42778 , n42779 );
xor ( n42782 , n41581 , n41776 );
nor ( n42783 , n9437 , n42643 );
and ( n42784 , n42782 , n42783 );
xor ( n42785 , n42782 , n42783 );
xor ( n42786 , n41585 , n41774 );
nor ( n42787 , n9446 , n42643 );
and ( n42788 , n42786 , n42787 );
xor ( n42789 , n42786 , n42787 );
xor ( n42790 , n41589 , n41772 );
nor ( n42791 , n9455 , n42643 );
and ( n42792 , n42790 , n42791 );
xor ( n42793 , n42790 , n42791 );
xor ( n42794 , n41593 , n41770 );
nor ( n42795 , n9464 , n42643 );
and ( n42796 , n42794 , n42795 );
xor ( n42797 , n42794 , n42795 );
xor ( n42798 , n41597 , n41768 );
nor ( n42799 , n9473 , n42643 );
and ( n42800 , n42798 , n42799 );
xor ( n42801 , n42798 , n42799 );
xor ( n42802 , n41601 , n41766 );
nor ( n42803 , n9482 , n42643 );
and ( n42804 , n42802 , n42803 );
xor ( n42805 , n42802 , n42803 );
xor ( n42806 , n41605 , n41764 );
nor ( n42807 , n9491 , n42643 );
and ( n42808 , n42806 , n42807 );
xor ( n42809 , n42806 , n42807 );
xor ( n42810 , n41609 , n41762 );
nor ( n42811 , n9500 , n42643 );
and ( n42812 , n42810 , n42811 );
xor ( n42813 , n42810 , n42811 );
xor ( n42814 , n41613 , n41760 );
nor ( n42815 , n9509 , n42643 );
and ( n42816 , n42814 , n42815 );
xor ( n42817 , n42814 , n42815 );
xor ( n42818 , n41617 , n41758 );
nor ( n42819 , n9518 , n42643 );
and ( n42820 , n42818 , n42819 );
xor ( n42821 , n42818 , n42819 );
xor ( n42822 , n41621 , n41756 );
nor ( n42823 , n9527 , n42643 );
and ( n42824 , n42822 , n42823 );
xor ( n42825 , n42822 , n42823 );
xor ( n42826 , n41625 , n41754 );
nor ( n42827 , n9536 , n42643 );
and ( n42828 , n42826 , n42827 );
xor ( n42829 , n42826 , n42827 );
xor ( n42830 , n41629 , n41752 );
nor ( n42831 , n9545 , n42643 );
and ( n42832 , n42830 , n42831 );
xor ( n42833 , n42830 , n42831 );
xor ( n42834 , n41633 , n41750 );
nor ( n42835 , n9554 , n42643 );
and ( n42836 , n42834 , n42835 );
xor ( n42837 , n42834 , n42835 );
xor ( n42838 , n41637 , n41748 );
nor ( n42839 , n9563 , n42643 );
and ( n42840 , n42838 , n42839 );
xor ( n42841 , n42838 , n42839 );
xor ( n42842 , n41641 , n41746 );
nor ( n42843 , n9572 , n42643 );
and ( n42844 , n42842 , n42843 );
xor ( n42845 , n42842 , n42843 );
xor ( n42846 , n41645 , n41744 );
nor ( n42847 , n9581 , n42643 );
and ( n42848 , n42846 , n42847 );
xor ( n42849 , n42846 , n42847 );
xor ( n42850 , n41649 , n41742 );
nor ( n42851 , n9590 , n42643 );
and ( n42852 , n42850 , n42851 );
xor ( n42853 , n42850 , n42851 );
xor ( n42854 , n41653 , n41740 );
nor ( n42855 , n9599 , n42643 );
and ( n42856 , n42854 , n42855 );
xor ( n42857 , n42854 , n42855 );
xor ( n42858 , n41657 , n41738 );
nor ( n42859 , n9608 , n42643 );
and ( n42860 , n42858 , n42859 );
xor ( n42861 , n42858 , n42859 );
xor ( n42862 , n41661 , n41736 );
nor ( n42863 , n9617 , n42643 );
and ( n42864 , n42862 , n42863 );
xor ( n42865 , n42862 , n42863 );
xor ( n42866 , n41665 , n41734 );
nor ( n42867 , n9626 , n42643 );
and ( n42868 , n42866 , n42867 );
xor ( n42869 , n42866 , n42867 );
xor ( n42870 , n41669 , n41732 );
nor ( n42871 , n9635 , n42643 );
and ( n42872 , n42870 , n42871 );
xor ( n42873 , n42870 , n42871 );
xor ( n42874 , n41673 , n41730 );
nor ( n42875 , n9644 , n42643 );
and ( n42876 , n42874 , n42875 );
xor ( n42877 , n42874 , n42875 );
xor ( n42878 , n41677 , n41728 );
nor ( n42879 , n9653 , n42643 );
and ( n42880 , n42878 , n42879 );
xor ( n42881 , n42878 , n42879 );
xor ( n42882 , n41681 , n41726 );
nor ( n42883 , n9662 , n42643 );
and ( n42884 , n42882 , n42883 );
xor ( n42885 , n42882 , n42883 );
xor ( n42886 , n41685 , n41724 );
nor ( n42887 , n9671 , n42643 );
and ( n42888 , n42886 , n42887 );
xor ( n42889 , n42886 , n42887 );
xor ( n42890 , n41689 , n41722 );
nor ( n42891 , n9680 , n42643 );
and ( n42892 , n42890 , n42891 );
xor ( n42893 , n42890 , n42891 );
xor ( n42894 , n41693 , n41720 );
nor ( n42895 , n9689 , n42643 );
and ( n42896 , n42894 , n42895 );
xor ( n42897 , n42894 , n42895 );
xor ( n42898 , n41697 , n41718 );
nor ( n42899 , n9698 , n42643 );
and ( n42900 , n42898 , n42899 );
xor ( n42901 , n42898 , n42899 );
xor ( n42902 , n41701 , n41716 );
nor ( n42903 , n9707 , n42643 );
and ( n42904 , n42902 , n42903 );
xor ( n42905 , n42902 , n42903 );
xor ( n42906 , n41705 , n41714 );
nor ( n42907 , n9716 , n42643 );
and ( n42908 , n42906 , n42907 );
xor ( n42909 , n42906 , n42907 );
xor ( n42910 , n41709 , n41712 );
nor ( n42911 , n9725 , n42643 );
and ( n42912 , n42910 , n42911 );
xor ( n42913 , n42910 , n42911 );
xor ( n42914 , n41710 , n41711 );
nor ( n42915 , n9734 , n42643 );
and ( n42916 , n42914 , n42915 );
xor ( n42917 , n42914 , n42915 );
nor ( n42918 , n9752 , n41439 );
nor ( n42919 , n9743 , n42643 );
and ( n42920 , n42918 , n42919 );
and ( n42921 , n42917 , n42920 );
or ( n42922 , n42916 , n42921 );
and ( n42923 , n42913 , n42922 );
or ( n42924 , n42912 , n42923 );
and ( n42925 , n42909 , n42924 );
or ( n42926 , n42908 , n42925 );
and ( n42927 , n42905 , n42926 );
or ( n42928 , n42904 , n42927 );
and ( n42929 , n42901 , n42928 );
or ( n42930 , n42900 , n42929 );
and ( n42931 , n42897 , n42930 );
or ( n42932 , n42896 , n42931 );
and ( n42933 , n42893 , n42932 );
or ( n42934 , n42892 , n42933 );
and ( n42935 , n42889 , n42934 );
or ( n42936 , n42888 , n42935 );
and ( n42937 , n42885 , n42936 );
or ( n42938 , n42884 , n42937 );
and ( n42939 , n42881 , n42938 );
or ( n42940 , n42880 , n42939 );
and ( n42941 , n42877 , n42940 );
or ( n42942 , n42876 , n42941 );
and ( n42943 , n42873 , n42942 );
or ( n42944 , n42872 , n42943 );
and ( n42945 , n42869 , n42944 );
or ( n42946 , n42868 , n42945 );
and ( n42947 , n42865 , n42946 );
or ( n42948 , n42864 , n42947 );
and ( n42949 , n42861 , n42948 );
or ( n42950 , n42860 , n42949 );
and ( n42951 , n42857 , n42950 );
or ( n42952 , n42856 , n42951 );
and ( n42953 , n42853 , n42952 );
or ( n42954 , n42852 , n42953 );
and ( n42955 , n42849 , n42954 );
or ( n42956 , n42848 , n42955 );
and ( n42957 , n42845 , n42956 );
or ( n42958 , n42844 , n42957 );
and ( n42959 , n42841 , n42958 );
or ( n42960 , n42840 , n42959 );
and ( n42961 , n42837 , n42960 );
or ( n42962 , n42836 , n42961 );
and ( n42963 , n42833 , n42962 );
or ( n42964 , n42832 , n42963 );
and ( n42965 , n42829 , n42964 );
or ( n42966 , n42828 , n42965 );
and ( n42967 , n42825 , n42966 );
or ( n42968 , n42824 , n42967 );
and ( n42969 , n42821 , n42968 );
or ( n42970 , n42820 , n42969 );
and ( n42971 , n42817 , n42970 );
or ( n42972 , n42816 , n42971 );
and ( n42973 , n42813 , n42972 );
or ( n42974 , n42812 , n42973 );
and ( n42975 , n42809 , n42974 );
or ( n42976 , n42808 , n42975 );
and ( n42977 , n42805 , n42976 );
or ( n42978 , n42804 , n42977 );
and ( n42979 , n42801 , n42978 );
or ( n42980 , n42800 , n42979 );
and ( n42981 , n42797 , n42980 );
or ( n42982 , n42796 , n42981 );
and ( n42983 , n42793 , n42982 );
or ( n42984 , n42792 , n42983 );
and ( n42985 , n42789 , n42984 );
or ( n42986 , n42788 , n42985 );
and ( n42987 , n42785 , n42986 );
or ( n42988 , n42784 , n42987 );
and ( n42989 , n42781 , n42988 );
or ( n42990 , n42780 , n42989 );
and ( n42991 , n42777 , n42990 );
or ( n42992 , n42776 , n42991 );
and ( n42993 , n42773 , n42992 );
or ( n42994 , n42772 , n42993 );
and ( n42995 , n42769 , n42994 );
or ( n42996 , n42768 , n42995 );
and ( n42997 , n42765 , n42996 );
or ( n42998 , n42764 , n42997 );
and ( n42999 , n42761 , n42998 );
or ( n43000 , n42760 , n42999 );
and ( n43001 , n42757 , n43000 );
or ( n43002 , n42756 , n43001 );
and ( n43003 , n42753 , n43002 );
or ( n43004 , n42752 , n43003 );
and ( n43005 , n42749 , n43004 );
or ( n43006 , n42748 , n43005 );
and ( n43007 , n42745 , n43006 );
or ( n43008 , n42744 , n43007 );
and ( n43009 , n42741 , n43008 );
or ( n43010 , n42740 , n43009 );
and ( n43011 , n42737 , n43010 );
or ( n43012 , n42736 , n43011 );
and ( n43013 , n42733 , n43012 );
or ( n43014 , n42732 , n43013 );
and ( n43015 , n42729 , n43014 );
or ( n43016 , n42728 , n43015 );
and ( n43017 , n42725 , n43016 );
or ( n43018 , n42724 , n43017 );
and ( n43019 , n42721 , n43018 );
or ( n43020 , n42720 , n43019 );
and ( n43021 , n42717 , n43020 );
or ( n43022 , n42716 , n43021 );
and ( n43023 , n42713 , n43022 );
or ( n43024 , n42712 , n43023 );
and ( n43025 , n42709 , n43024 );
or ( n43026 , n42708 , n43025 );
and ( n43027 , n42705 , n43026 );
or ( n43028 , n42704 , n43027 );
and ( n43029 , n42701 , n43028 );
or ( n43030 , n42700 , n43029 );
and ( n43031 , n42697 , n43030 );
or ( n43032 , n42696 , n43031 );
and ( n43033 , n42693 , n43032 );
or ( n43034 , n42692 , n43033 );
and ( n43035 , n42689 , n43034 );
or ( n43036 , n42688 , n43035 );
and ( n43037 , n42685 , n43036 );
or ( n43038 , n42684 , n43037 );
and ( n43039 , n42681 , n43038 );
or ( n43040 , n42680 , n43039 );
and ( n43041 , n42677 , n43040 );
or ( n43042 , n42676 , n43041 );
and ( n43043 , n42673 , n43042 );
or ( n43044 , n42672 , n43043 );
and ( n43045 , n42669 , n43044 );
or ( n43046 , n42668 , n43045 );
and ( n43047 , n42665 , n43046 );
or ( n43048 , n42664 , n43047 );
and ( n43049 , n42661 , n43048 );
or ( n43050 , n42660 , n43049 );
and ( n43051 , n42657 , n43050 );
or ( n43052 , n42656 , n43051 );
and ( n43053 , n42653 , n43052 );
or ( n43054 , n42652 , n43053 );
and ( n43055 , n42649 , n43054 );
or ( n43056 , n42648 , n43055 );
xor ( n43057 , n42645 , n43056 );
and ( n43058 , n33403 , n957 );
nor ( n43059 , n958 , n43058 );
nor ( n43060 , n1062 , n32231 );
xor ( n43061 , n43059 , n43060 );
and ( n43062 , n41849 , n41850 );
and ( n43063 , n41851 , n41854 );
or ( n43064 , n43062 , n43063 );
xor ( n43065 , n43061 , n43064 );
nor ( n43066 , n1176 , n31083 );
xor ( n43067 , n43065 , n43066 );
and ( n43068 , n41855 , n41856 );
and ( n43069 , n41857 , n41860 );
or ( n43070 , n43068 , n43069 );
xor ( n43071 , n43067 , n43070 );
nor ( n43072 , n1303 , n29948 );
xor ( n43073 , n43071 , n43072 );
and ( n43074 , n41861 , n41862 );
and ( n43075 , n41863 , n41866 );
or ( n43076 , n43074 , n43075 );
xor ( n43077 , n43073 , n43076 );
nor ( n43078 , n1445 , n28833 );
xor ( n43079 , n43077 , n43078 );
and ( n43080 , n41867 , n41868 );
and ( n43081 , n41869 , n41872 );
or ( n43082 , n43080 , n43081 );
xor ( n43083 , n43079 , n43082 );
nor ( n43084 , n1598 , n27737 );
xor ( n43085 , n43083 , n43084 );
and ( n43086 , n41873 , n41874 );
and ( n43087 , n41875 , n41878 );
or ( n43088 , n43086 , n43087 );
xor ( n43089 , n43085 , n43088 );
nor ( n43090 , n1766 , n26660 );
xor ( n43091 , n43089 , n43090 );
and ( n43092 , n41879 , n41880 );
and ( n43093 , n41881 , n41884 );
or ( n43094 , n43092 , n43093 );
xor ( n43095 , n43091 , n43094 );
nor ( n43096 , n1945 , n25600 );
xor ( n43097 , n43095 , n43096 );
and ( n43098 , n41885 , n41886 );
and ( n43099 , n41887 , n41890 );
or ( n43100 , n43098 , n43099 );
xor ( n43101 , n43097 , n43100 );
nor ( n43102 , n2137 , n24564 );
xor ( n43103 , n43101 , n43102 );
and ( n43104 , n41891 , n41892 );
and ( n43105 , n41893 , n41896 );
or ( n43106 , n43104 , n43105 );
xor ( n43107 , n43103 , n43106 );
nor ( n43108 , n2343 , n23541 );
xor ( n43109 , n43107 , n43108 );
and ( n43110 , n41897 , n41898 );
and ( n43111 , n41899 , n41902 );
or ( n43112 , n43110 , n43111 );
xor ( n43113 , n43109 , n43112 );
nor ( n43114 , n2566 , n22541 );
xor ( n43115 , n43113 , n43114 );
and ( n43116 , n41903 , n41904 );
and ( n43117 , n41905 , n41908 );
or ( n43118 , n43116 , n43117 );
xor ( n43119 , n43115 , n43118 );
nor ( n43120 , n2797 , n21562 );
xor ( n43121 , n43119 , n43120 );
and ( n43122 , n41909 , n41910 );
and ( n43123 , n41911 , n41914 );
or ( n43124 , n43122 , n43123 );
xor ( n43125 , n43121 , n43124 );
nor ( n43126 , n3043 , n20601 );
xor ( n43127 , n43125 , n43126 );
and ( n43128 , n41915 , n41916 );
and ( n43129 , n41917 , n41920 );
or ( n43130 , n43128 , n43129 );
xor ( n43131 , n43127 , n43130 );
nor ( n43132 , n3300 , n19657 );
xor ( n43133 , n43131 , n43132 );
and ( n43134 , n41921 , n41922 );
and ( n43135 , n41923 , n41926 );
or ( n43136 , n43134 , n43135 );
xor ( n43137 , n43133 , n43136 );
nor ( n43138 , n3570 , n18734 );
xor ( n43139 , n43137 , n43138 );
and ( n43140 , n41927 , n41928 );
and ( n43141 , n41929 , n41932 );
or ( n43142 , n43140 , n43141 );
xor ( n43143 , n43139 , n43142 );
nor ( n43144 , n3853 , n17828 );
xor ( n43145 , n43143 , n43144 );
and ( n43146 , n41933 , n41934 );
and ( n43147 , n41935 , n41938 );
or ( n43148 , n43146 , n43147 );
xor ( n43149 , n43145 , n43148 );
nor ( n43150 , n4151 , n16943 );
xor ( n43151 , n43149 , n43150 );
and ( n43152 , n41939 , n41940 );
and ( n43153 , n41941 , n41944 );
or ( n43154 , n43152 , n43153 );
xor ( n43155 , n43151 , n43154 );
nor ( n43156 , n4458 , n16077 );
xor ( n43157 , n43155 , n43156 );
and ( n43158 , n41945 , n41946 );
and ( n43159 , n41947 , n41950 );
or ( n43160 , n43158 , n43159 );
xor ( n43161 , n43157 , n43160 );
nor ( n43162 , n4786 , n15230 );
xor ( n43163 , n43161 , n43162 );
and ( n43164 , n41951 , n41952 );
and ( n43165 , n41953 , n41956 );
or ( n43166 , n43164 , n43165 );
xor ( n43167 , n43163 , n43166 );
nor ( n43168 , n5126 , n14403 );
xor ( n43169 , n43167 , n43168 );
and ( n43170 , n41957 , n41958 );
and ( n43171 , n41959 , n41962 );
or ( n43172 , n43170 , n43171 );
xor ( n43173 , n43169 , n43172 );
nor ( n43174 , n5477 , n13599 );
xor ( n43175 , n43173 , n43174 );
and ( n43176 , n41963 , n41964 );
and ( n43177 , n41965 , n41968 );
or ( n43178 , n43176 , n43177 );
xor ( n43179 , n43175 , n43178 );
nor ( n43180 , n5838 , n12808 );
xor ( n43181 , n43179 , n43180 );
and ( n43182 , n41969 , n41970 );
and ( n43183 , n41971 , n41974 );
or ( n43184 , n43182 , n43183 );
xor ( n43185 , n43181 , n43184 );
nor ( n43186 , n6212 , n12037 );
xor ( n43187 , n43185 , n43186 );
and ( n43188 , n41975 , n41976 );
and ( n43189 , n41977 , n41980 );
or ( n43190 , n43188 , n43189 );
xor ( n43191 , n43187 , n43190 );
nor ( n43192 , n6596 , n11282 );
xor ( n43193 , n43191 , n43192 );
and ( n43194 , n41981 , n41982 );
and ( n43195 , n41983 , n41986 );
or ( n43196 , n43194 , n43195 );
xor ( n43197 , n43193 , n43196 );
nor ( n43198 , n6997 , n10547 );
xor ( n43199 , n43197 , n43198 );
and ( n43200 , n41987 , n41988 );
and ( n43201 , n41989 , n41992 );
or ( n43202 , n43200 , n43201 );
xor ( n43203 , n43199 , n43202 );
nor ( n43204 , n7413 , n9829 );
xor ( n43205 , n43203 , n43204 );
and ( n43206 , n41993 , n41994 );
and ( n43207 , n41995 , n41998 );
or ( n43208 , n43206 , n43207 );
xor ( n43209 , n43205 , n43208 );
nor ( n43210 , n7841 , n8955 );
xor ( n43211 , n43209 , n43210 );
and ( n43212 , n41999 , n42000 );
and ( n43213 , n42001 , n42004 );
or ( n43214 , n43212 , n43213 );
xor ( n43215 , n43211 , n43214 );
nor ( n43216 , n8281 , n603 );
xor ( n43217 , n43215 , n43216 );
and ( n43218 , n42005 , n42006 );
and ( n43219 , n42007 , n42010 );
or ( n43220 , n43218 , n43219 );
xor ( n43221 , n43217 , n43220 );
nor ( n43222 , n8737 , n652 );
xor ( n43223 , n43221 , n43222 );
and ( n43224 , n42011 , n42012 );
and ( n43225 , n42013 , n42016 );
or ( n43226 , n43224 , n43225 );
xor ( n43227 , n43223 , n43226 );
nor ( n43228 , n9420 , n624 );
xor ( n43229 , n43227 , n43228 );
and ( n43230 , n42017 , n42018 );
and ( n43231 , n42019 , n42022 );
or ( n43232 , n43230 , n43231 );
xor ( n43233 , n43229 , n43232 );
nor ( n43234 , n10312 , n648 );
xor ( n43235 , n43233 , n43234 );
and ( n43236 , n42023 , n42024 );
and ( n43237 , n42025 , n42028 );
or ( n43238 , n43236 , n43237 );
xor ( n43239 , n43235 , n43238 );
nor ( n43240 , n11041 , n686 );
xor ( n43241 , n43239 , n43240 );
and ( n43242 , n42029 , n42030 );
and ( n43243 , n42031 , n42034 );
or ( n43244 , n43242 , n43243 );
xor ( n43245 , n43241 , n43244 );
nor ( n43246 , n11790 , n735 );
xor ( n43247 , n43245 , n43246 );
and ( n43248 , n42035 , n42036 );
and ( n43249 , n42037 , n42040 );
or ( n43250 , n43248 , n43249 );
xor ( n43251 , n43247 , n43250 );
nor ( n43252 , n12555 , n798 );
xor ( n43253 , n43251 , n43252 );
and ( n43254 , n42041 , n42042 );
and ( n43255 , n42043 , n42046 );
or ( n43256 , n43254 , n43255 );
xor ( n43257 , n43253 , n43256 );
nor ( n43258 , n13340 , n870 );
xor ( n43259 , n43257 , n43258 );
and ( n43260 , n42047 , n42048 );
and ( n43261 , n42049 , n42052 );
or ( n43262 , n43260 , n43261 );
xor ( n43263 , n43259 , n43262 );
nor ( n43264 , n14138 , n960 );
xor ( n43265 , n43263 , n43264 );
and ( n43266 , n42053 , n42054 );
and ( n43267 , n42055 , n42058 );
or ( n43268 , n43266 , n43267 );
xor ( n43269 , n43265 , n43268 );
nor ( n43270 , n14959 , n1064 );
xor ( n43271 , n43269 , n43270 );
and ( n43272 , n42059 , n42060 );
and ( n43273 , n42061 , n42064 );
or ( n43274 , n43272 , n43273 );
xor ( n43275 , n43271 , n43274 );
nor ( n43276 , n15800 , n1178 );
xor ( n43277 , n43275 , n43276 );
and ( n43278 , n42065 , n42066 );
and ( n43279 , n42067 , n42070 );
or ( n43280 , n43278 , n43279 );
xor ( n43281 , n43277 , n43280 );
nor ( n43282 , n16660 , n1305 );
xor ( n43283 , n43281 , n43282 );
and ( n43284 , n42071 , n42072 );
and ( n43285 , n42073 , n42076 );
or ( n43286 , n43284 , n43285 );
xor ( n43287 , n43283 , n43286 );
nor ( n43288 , n17539 , n1447 );
xor ( n43289 , n43287 , n43288 );
and ( n43290 , n42077 , n42078 );
and ( n43291 , n42079 , n42082 );
or ( n43292 , n43290 , n43291 );
xor ( n43293 , n43289 , n43292 );
nor ( n43294 , n18439 , n1600 );
xor ( n43295 , n43293 , n43294 );
and ( n43296 , n42083 , n42084 );
and ( n43297 , n42085 , n42088 );
or ( n43298 , n43296 , n43297 );
xor ( n43299 , n43295 , n43298 );
nor ( n43300 , n19356 , n1768 );
xor ( n43301 , n43299 , n43300 );
and ( n43302 , n42089 , n42090 );
and ( n43303 , n42091 , n42094 );
or ( n43304 , n43302 , n43303 );
xor ( n43305 , n43301 , n43304 );
nor ( n43306 , n20294 , n1947 );
xor ( n43307 , n43305 , n43306 );
and ( n43308 , n42095 , n42096 );
and ( n43309 , n42097 , n42100 );
or ( n43310 , n43308 , n43309 );
xor ( n43311 , n43307 , n43310 );
nor ( n43312 , n21249 , n2139 );
xor ( n43313 , n43311 , n43312 );
and ( n43314 , n42101 , n42102 );
and ( n43315 , n42103 , n42106 );
or ( n43316 , n43314 , n43315 );
xor ( n43317 , n43313 , n43316 );
nor ( n43318 , n22222 , n2345 );
xor ( n43319 , n43317 , n43318 );
and ( n43320 , n42107 , n42108 );
and ( n43321 , n42109 , n42112 );
or ( n43322 , n43320 , n43321 );
xor ( n43323 , n43319 , n43322 );
nor ( n43324 , n23216 , n2568 );
xor ( n43325 , n43323 , n43324 );
and ( n43326 , n42113 , n42114 );
and ( n43327 , n42115 , n42118 );
or ( n43328 , n43326 , n43327 );
xor ( n43329 , n43325 , n43328 );
nor ( n43330 , n24233 , n2799 );
xor ( n43331 , n43329 , n43330 );
and ( n43332 , n42119 , n42120 );
and ( n43333 , n42121 , n42124 );
or ( n43334 , n43332 , n43333 );
xor ( n43335 , n43331 , n43334 );
nor ( n43336 , n25263 , n3045 );
xor ( n43337 , n43335 , n43336 );
and ( n43338 , n42125 , n42126 );
and ( n43339 , n42127 , n42130 );
or ( n43340 , n43338 , n43339 );
xor ( n43341 , n43337 , n43340 );
nor ( n43342 , n26317 , n3302 );
xor ( n43343 , n43341 , n43342 );
and ( n43344 , n42131 , n42132 );
and ( n43345 , n42133 , n42136 );
or ( n43346 , n43344 , n43345 );
xor ( n43347 , n43343 , n43346 );
nor ( n43348 , n27388 , n3572 );
xor ( n43349 , n43347 , n43348 );
and ( n43350 , n42137 , n42138 );
and ( n43351 , n42139 , n42142 );
or ( n43352 , n43350 , n43351 );
xor ( n43353 , n43349 , n43352 );
nor ( n43354 , n28478 , n3855 );
xor ( n43355 , n43353 , n43354 );
and ( n43356 , n42143 , n42144 );
and ( n43357 , n42145 , n42148 );
or ( n43358 , n43356 , n43357 );
xor ( n43359 , n43355 , n43358 );
nor ( n43360 , n29587 , n4153 );
xor ( n43361 , n43359 , n43360 );
and ( n43362 , n42149 , n42150 );
and ( n43363 , n42151 , n42154 );
or ( n43364 , n43362 , n43363 );
xor ( n43365 , n43361 , n43364 );
nor ( n43366 , n30716 , n4460 );
xor ( n43367 , n43365 , n43366 );
and ( n43368 , n42155 , n42156 );
and ( n43369 , n42157 , n42160 );
or ( n43370 , n43368 , n43369 );
xor ( n43371 , n43367 , n43370 );
nor ( n43372 , n31858 , n4788 );
xor ( n43373 , n43371 , n43372 );
and ( n43374 , n42161 , n42162 );
and ( n43375 , n42163 , n42166 );
or ( n43376 , n43374 , n43375 );
xor ( n43377 , n43373 , n43376 );
nor ( n43378 , n33024 , n5128 );
xor ( n43379 , n43377 , n43378 );
and ( n43380 , n42167 , n42168 );
and ( n43381 , n42169 , n42172 );
or ( n43382 , n43380 , n43381 );
xor ( n43383 , n43379 , n43382 );
nor ( n43384 , n34215 , n5479 );
xor ( n43385 , n43383 , n43384 );
and ( n43386 , n42173 , n42174 );
and ( n43387 , n42175 , n42178 );
or ( n43388 , n43386 , n43387 );
xor ( n43389 , n43385 , n43388 );
nor ( n43390 , n35410 , n5840 );
xor ( n43391 , n43389 , n43390 );
and ( n43392 , n42179 , n42180 );
and ( n43393 , n42181 , n42184 );
or ( n43394 , n43392 , n43393 );
xor ( n43395 , n43391 , n43394 );
nor ( n43396 , n36611 , n6214 );
xor ( n43397 , n43395 , n43396 );
and ( n43398 , n42185 , n42186 );
and ( n43399 , n42187 , n42190 );
or ( n43400 , n43398 , n43399 );
xor ( n43401 , n43397 , n43400 );
nor ( n43402 , n37816 , n6598 );
xor ( n43403 , n43401 , n43402 );
and ( n43404 , n42191 , n42192 );
and ( n43405 , n42193 , n42196 );
or ( n43406 , n43404 , n43405 );
xor ( n43407 , n43403 , n43406 );
nor ( n43408 , n39018 , n6999 );
xor ( n43409 , n43407 , n43408 );
and ( n43410 , n42197 , n42198 );
and ( n43411 , n42199 , n42202 );
or ( n43412 , n43410 , n43411 );
xor ( n43413 , n43409 , n43412 );
nor ( n43414 , n40223 , n7415 );
xor ( n43415 , n43413 , n43414 );
and ( n43416 , n42203 , n42204 );
and ( n43417 , n42205 , n42208 );
or ( n43418 , n43416 , n43417 );
xor ( n43419 , n43415 , n43418 );
nor ( n43420 , n41428 , n7843 );
xor ( n43421 , n43419 , n43420 );
and ( n43422 , n42209 , n42210 );
and ( n43423 , n42211 , n42214 );
or ( n43424 , n43422 , n43423 );
xor ( n43425 , n43421 , n43424 );
nor ( n43426 , n42632 , n8283 );
xor ( n43427 , n43425 , n43426 );
and ( n43428 , n42215 , n42216 );
and ( n43429 , n42217 , n42220 );
or ( n43430 , n43428 , n43429 );
xor ( n43431 , n43427 , n43430 );
and ( n43432 , n42233 , n42237 );
and ( n43433 , n42237 , n42618 );
and ( n43434 , n42233 , n42618 );
or ( n43435 , n43432 , n43433 , n43434 );
and ( n43436 , n33774 , n940 );
not ( n43437 , n940 );
nor ( n43438 , n43436 , n43437 );
xor ( n43439 , n43435 , n43438 );
and ( n43440 , n42246 , n42250 );
and ( n43441 , n42250 , n42318 );
and ( n43442 , n42246 , n42318 );
or ( n43443 , n43440 , n43441 , n43442 );
and ( n43444 , n42242 , n42319 );
and ( n43445 , n42319 , n42617 );
and ( n43446 , n42242 , n42617 );
or ( n43447 , n43444 , n43445 , n43446 );
xor ( n43448 , n43443 , n43447 );
and ( n43449 , n42324 , n42444 );
and ( n43450 , n42444 , n42616 );
and ( n43451 , n42324 , n42616 );
or ( n43452 , n43449 , n43450 , n43451 );
and ( n43453 , n42255 , n42259 );
and ( n43454 , n42259 , n42317 );
and ( n43455 , n42255 , n42317 );
or ( n43456 , n43453 , n43454 , n43455 );
and ( n43457 , n42328 , n42332 );
and ( n43458 , n42332 , n42443 );
and ( n43459 , n42328 , n42443 );
or ( n43460 , n43457 , n43458 , n43459 );
xor ( n43461 , n43456 , n43460 );
and ( n43462 , n42286 , n42290 );
and ( n43463 , n42290 , n42296 );
and ( n43464 , n42286 , n42296 );
or ( n43465 , n43462 , n43463 , n43464 );
and ( n43466 , n42264 , n42268 );
and ( n43467 , n42268 , n42316 );
and ( n43468 , n42264 , n42316 );
or ( n43469 , n43466 , n43467 , n43468 );
xor ( n43470 , n43465 , n43469 );
and ( n43471 , n42273 , n42277 );
and ( n43472 , n42277 , n42315 );
and ( n43473 , n42273 , n42315 );
or ( n43474 , n43471 , n43472 , n43473 );
and ( n43475 , n42341 , n42366 );
and ( n43476 , n42366 , n42404 );
and ( n43477 , n42341 , n42404 );
or ( n43478 , n43475 , n43476 , n43477 );
xor ( n43479 , n43474 , n43478 );
and ( n43480 , n42282 , n42297 );
and ( n43481 , n42297 , n42314 );
and ( n43482 , n42282 , n42314 );
or ( n43483 , n43480 , n43481 , n43482 );
and ( n43484 , n42345 , n42349 );
and ( n43485 , n42349 , n42365 );
and ( n43486 , n42345 , n42365 );
or ( n43487 , n43484 , n43485 , n43486 );
xor ( n43488 , n43483 , n43487 );
and ( n43489 , n42302 , n42307 );
and ( n43490 , n42307 , n42313 );
and ( n43491 , n42302 , n42313 );
or ( n43492 , n43489 , n43490 , n43491 );
and ( n43493 , n42292 , n42293 );
and ( n43494 , n42293 , n42295 );
and ( n43495 , n42292 , n42295 );
or ( n43496 , n43493 , n43494 , n43495 );
and ( n43497 , n42303 , n42304 );
and ( n43498 , n42304 , n42306 );
and ( n43499 , n42303 , n42306 );
or ( n43500 , n43497 , n43498 , n43499 );
xor ( n43501 , n43496 , n43500 );
and ( n43502 , n30695 , n1254 );
and ( n43503 , n31836 , n1134 );
xor ( n43504 , n43502 , n43503 );
and ( n43505 , n32649 , n1034 );
xor ( n43506 , n43504 , n43505 );
xor ( n43507 , n43501 , n43506 );
xor ( n43508 , n43492 , n43507 );
and ( n43509 , n42309 , n42310 );
and ( n43510 , n42310 , n42312 );
and ( n43511 , n42309 , n42312 );
or ( n43512 , n43509 , n43510 , n43511 );
and ( n43513 , n27361 , n1738 );
and ( n43514 , n28456 , n1551 );
xor ( n43515 , n43513 , n43514 );
and ( n43516 , n29559 , n1424 );
xor ( n43517 , n43515 , n43516 );
xor ( n43518 , n43512 , n43517 );
and ( n43519 , n24214 , n2298 );
and ( n43520 , n25243 , n2100 );
xor ( n43521 , n43519 , n43520 );
and ( n43522 , n26296 , n1882 );
xor ( n43523 , n43521 , n43522 );
xor ( n43524 , n43518 , n43523 );
xor ( n43525 , n43508 , n43524 );
xor ( n43526 , n43488 , n43525 );
xor ( n43527 , n43479 , n43526 );
xor ( n43528 , n43470 , n43527 );
xor ( n43529 , n43461 , n43528 );
xor ( n43530 , n43452 , n43529 );
and ( n43531 , n42449 , n42527 );
and ( n43532 , n42527 , n42615 );
and ( n43533 , n42449 , n42615 );
or ( n43534 , n43531 , n43532 , n43533 );
and ( n43535 , n42337 , n42405 );
and ( n43536 , n42405 , n42442 );
and ( n43537 , n42337 , n42442 );
or ( n43538 , n43535 , n43536 , n43537 );
and ( n43539 , n42453 , n42457 );
and ( n43540 , n42457 , n42526 );
and ( n43541 , n42453 , n42526 );
or ( n43542 , n43539 , n43540 , n43541 );
xor ( n43543 , n43538 , n43542 );
and ( n43544 , n42410 , n42414 );
and ( n43545 , n42414 , n42441 );
and ( n43546 , n42410 , n42441 );
or ( n43547 , n43544 , n43545 , n43546 );
and ( n43548 , n42371 , n42387 );
and ( n43549 , n42387 , n42403 );
and ( n43550 , n42371 , n42403 );
or ( n43551 , n43548 , n43549 , n43550 );
and ( n43552 , n42354 , n42358 );
and ( n43553 , n42358 , n42364 );
and ( n43554 , n42354 , n42364 );
or ( n43555 , n43552 , n43553 , n43554 );
and ( n43556 , n42375 , n42380 );
and ( n43557 , n42380 , n42386 );
and ( n43558 , n42375 , n42386 );
or ( n43559 , n43556 , n43557 , n43558 );
xor ( n43560 , n43555 , n43559 );
and ( n43561 , n42360 , n42361 );
and ( n43562 , n42361 , n42363 );
and ( n43563 , n42360 , n42363 );
or ( n43564 , n43561 , n43562 , n43563 );
and ( n43565 , n42376 , n42377 );
and ( n43566 , n42377 , n42379 );
and ( n43567 , n42376 , n42379 );
or ( n43568 , n43565 , n43566 , n43567 );
xor ( n43569 , n43564 , n43568 );
and ( n43570 , n21216 , n2981 );
and ( n43571 , n22186 , n2739 );
xor ( n43572 , n43570 , n43571 );
and ( n43573 , n22892 , n2544 );
xor ( n43574 , n43572 , n43573 );
xor ( n43575 , n43569 , n43574 );
xor ( n43576 , n43560 , n43575 );
xor ( n43577 , n43551 , n43576 );
and ( n43578 , n42392 , n42396 );
and ( n43579 , n42396 , n42402 );
and ( n43580 , n42392 , n42402 );
or ( n43581 , n43578 , n43579 , n43580 );
and ( n43582 , n42382 , n42383 );
and ( n43583 , n42383 , n42385 );
and ( n43584 , n42382 , n42385 );
or ( n43585 , n43582 , n43583 , n43584 );
and ( n43586 , n18144 , n3749 );
and ( n43587 , n19324 , n3495 );
xor ( n43588 , n43586 , n43587 );
and ( n43589 , n20233 , n3271 );
xor ( n43590 , n43588 , n43589 );
xor ( n43591 , n43585 , n43590 );
and ( n43592 , n15758 , n4730 );
and ( n43593 , n16637 , n4403 );
xor ( n43594 , n43592 , n43593 );
and ( n43595 , n17512 , n4102 );
xor ( n43596 , n43594 , n43595 );
xor ( n43597 , n43591 , n43596 );
xor ( n43598 , n43581 , n43597 );
and ( n43599 , n42398 , n42399 );
and ( n43600 , n42399 , n42401 );
and ( n43601 , n42398 , n42401 );
or ( n43602 , n43599 , n43600 , n43601 );
and ( n43603 , n42429 , n42430 );
and ( n43604 , n42430 , n42432 );
and ( n43605 , n42429 , n42432 );
or ( n43606 , n43603 , n43604 , n43605 );
xor ( n43607 , n43602 , n43606 );
and ( n43608 , n13322 , n5765 );
and ( n43609 , n14118 , n5408 );
xor ( n43610 , n43608 , n43609 );
and ( n43611 , n14938 , n5103 );
xor ( n43612 , n43610 , n43611 );
xor ( n43613 , n43607 , n43612 );
xor ( n43614 , n43598 , n43613 );
xor ( n43615 , n43577 , n43614 );
xor ( n43616 , n43547 , n43615 );
and ( n43617 , n42419 , n42423 );
and ( n43618 , n42423 , n42440 );
and ( n43619 , n42419 , n42440 );
or ( n43620 , n43617 , n43618 , n43619 );
and ( n43621 , n42466 , n42481 );
and ( n43622 , n42481 , n42498 );
and ( n43623 , n42466 , n42498 );
or ( n43624 , n43621 , n43622 , n43623 );
xor ( n43625 , n43620 , n43624 );
and ( n43626 , n42428 , n42433 );
and ( n43627 , n42433 , n42439 );
and ( n43628 , n42428 , n42439 );
or ( n43629 , n43626 , n43627 , n43628 );
and ( n43630 , n42470 , n42474 );
and ( n43631 , n42474 , n42480 );
and ( n43632 , n42470 , n42480 );
or ( n43633 , n43630 , n43631 , n43632 );
xor ( n43634 , n43629 , n43633 );
and ( n43635 , n42435 , n42436 );
and ( n43636 , n42436 , n42438 );
and ( n43637 , n42435 , n42438 );
or ( n43638 , n43635 , n43636 , n43637 );
and ( n43639 , n11015 , n6971 );
and ( n43640 , n11769 , n6504 );
xor ( n43641 , n43639 , n43640 );
and ( n43642 , n12320 , n6132 );
xor ( n43643 , n43641 , n43642 );
xor ( n43644 , n43638 , n43643 );
and ( n43645 , n8718 , n8243 );
and ( n43646 , n9400 , n7662 );
xor ( n43647 , n43645 , n43646 );
and ( n43648 , n10291 , n7310 );
xor ( n43649 , n43647 , n43648 );
xor ( n43650 , n43644 , n43649 );
xor ( n43651 , n43634 , n43650 );
xor ( n43652 , n43625 , n43651 );
xor ( n43653 , n43616 , n43652 );
xor ( n43654 , n43543 , n43653 );
xor ( n43655 , n43534 , n43654 );
and ( n43656 , n42532 , n42579 );
and ( n43657 , n42579 , n42614 );
and ( n43658 , n42532 , n42614 );
or ( n43659 , n43656 , n43657 , n43658 );
and ( n43660 , n42462 , n42499 );
and ( n43661 , n42499 , n42525 );
and ( n43662 , n42462 , n42525 );
or ( n43663 , n43660 , n43661 , n43662 );
and ( n43664 , n42536 , n42540 );
and ( n43665 , n42540 , n42578 );
and ( n43666 , n42536 , n42578 );
or ( n43667 , n43664 , n43665 , n43666 );
xor ( n43668 , n43663 , n43667 );
and ( n43669 , n42504 , n42508 );
and ( n43670 , n42508 , n42524 );
and ( n43671 , n42504 , n42524 );
or ( n43672 , n43669 , n43670 , n43671 );
and ( n43673 , n42486 , n42491 );
and ( n43674 , n42491 , n42497 );
and ( n43675 , n42486 , n42497 );
or ( n43676 , n43673 , n43674 , n43675 );
and ( n43677 , n42476 , n42477 );
and ( n43678 , n42477 , n42479 );
and ( n43679 , n42476 , n42479 );
or ( n43680 , n43677 , n43678 , n43679 );
and ( n43681 , n42487 , n42488 );
and ( n43682 , n42488 , n42490 );
and ( n43683 , n42487 , n42490 );
or ( n43684 , n43681 , n43682 , n43683 );
xor ( n43685 , n43680 , n43684 );
and ( n43686 , n7385 , n10239 );
and ( n43687 , n7808 , n9348 );
xor ( n43688 , n43686 , n43687 );
and ( n43689 , n8079 , n8669 );
xor ( n43690 , n43688 , n43689 );
xor ( n43691 , n43685 , n43690 );
xor ( n43692 , n43676 , n43691 );
and ( n43693 , n42493 , n42494 );
and ( n43694 , n42494 , n42496 );
and ( n43695 , n42493 , n42496 );
or ( n43696 , n43693 , n43694 , n43695 );
and ( n43697 , n6187 , n12531 );
and ( n43698 , n6569 , n11718 );
xor ( n43699 , n43697 , n43698 );
and ( n43700 , n6816 , n10977 );
xor ( n43701 , n43699 , n43700 );
xor ( n43702 , n43696 , n43701 );
and ( n43703 , n4959 , n14838 );
and ( n43704 , n5459 , n14044 );
xor ( n43705 , n43703 , n43704 );
and ( n43706 , n5819 , n13256 );
xor ( n43707 , n43705 , n43706 );
xor ( n43708 , n43702 , n43707 );
xor ( n43709 , n43692 , n43708 );
xor ( n43710 , n43672 , n43709 );
and ( n43711 , n42513 , n42517 );
and ( n43712 , n42517 , n42523 );
and ( n43713 , n42513 , n42523 );
or ( n43714 , n43711 , n43712 , n43713 );
and ( n43715 , n42549 , n42554 );
and ( n43716 , n42554 , n42560 );
and ( n43717 , n42549 , n42560 );
or ( n43718 , n43715 , n43716 , n43717 );
xor ( n43719 , n43714 , n43718 );
and ( n43720 , n42519 , n42520 );
and ( n43721 , n42520 , n42522 );
and ( n43722 , n42519 , n42522 );
or ( n43723 , n43720 , n43721 , n43722 );
and ( n43724 , n42550 , n42551 );
and ( n43725 , n42551 , n42553 );
and ( n43726 , n42550 , n42553 );
or ( n43727 , n43724 , n43725 , n43726 );
xor ( n43728 , n43723 , n43727 );
and ( n43729 , n4132 , n17422 );
and ( n43730 , n4438 , n16550 );
xor ( n43731 , n43729 , n43730 );
and ( n43732 , n4766 , n15691 );
xor ( n43733 , n43731 , n43732 );
xor ( n43734 , n43728 , n43733 );
xor ( n43735 , n43719 , n43734 );
xor ( n43736 , n43710 , n43735 );
xor ( n43737 , n43668 , n43736 );
xor ( n43738 , n43659 , n43737 );
and ( n43739 , n42603 , n42613 );
and ( n43740 , n42584 , n42585 );
and ( n43741 , n42585 , n42602 );
and ( n43742 , n42584 , n42602 );
or ( n43743 , n43740 , n43741 , n43742 );
and ( n43744 , n42545 , n42561 );
and ( n43745 , n42561 , n42577 );
and ( n43746 , n42545 , n42577 );
or ( n43747 , n43744 , n43745 , n43746 );
xor ( n43748 , n43743 , n43747 );
and ( n43749 , n42566 , n42570 );
and ( n43750 , n42570 , n42576 );
and ( n43751 , n42566 , n42576 );
or ( n43752 , n43749 , n43750 , n43751 );
and ( n43753 , n42556 , n42557 );
and ( n43754 , n42557 , n42559 );
and ( n43755 , n42556 , n42559 );
or ( n43756 , n43753 , n43754 , n43755 );
and ( n43757 , n3182 , n20156 );
and ( n43758 , n3545 , n19222 );
xor ( n43759 , n43757 , n43758 );
and ( n43760 , n3801 , n18407 );
xor ( n43761 , n43759 , n43760 );
xor ( n43762 , n43756 , n43761 );
and ( n43763 , n2462 , n23075 );
and ( n43764 , n2779 , n22065 );
xor ( n43765 , n43763 , n43764 );
and ( n43766 , n3024 , n20976 );
xor ( n43767 , n43765 , n43766 );
xor ( n43768 , n43762 , n43767 );
xor ( n43769 , n43752 , n43768 );
and ( n43770 , n42572 , n42573 );
and ( n43771 , n42573 , n42575 );
and ( n43772 , n42572 , n42575 );
or ( n43773 , n43770 , n43771 , n43772 );
and ( n43774 , n42597 , n42598 );
and ( n43775 , n42598 , n42600 );
and ( n43776 , n42597 , n42600 );
or ( n43777 , n43774 , n43775 , n43776 );
xor ( n43778 , n43773 , n43777 );
and ( n43779 , n1933 , n26216 );
and ( n43780 , n2120 , n25163 );
xor ( n43781 , n43779 , n43780 );
and ( n43782 , n2324 , n24137 );
xor ( n43783 , n43781 , n43782 );
xor ( n43784 , n43778 , n43783 );
xor ( n43785 , n43769 , n43784 );
xor ( n43786 , n43748 , n43785 );
xor ( n43787 , n43739 , n43786 );
and ( n43788 , n42590 , n42595 );
and ( n43789 , n42595 , n42601 );
and ( n43790 , n42590 , n42601 );
or ( n43791 , n43788 , n43789 , n43790 );
and ( n43792 , n42607 , n42612 );
xor ( n43793 , n43791 , n43792 );
and ( n43794 , n42591 , n42592 );
and ( n43795 , n42592 , n42594 );
and ( n43796 , n42591 , n42594 );
or ( n43797 , n43794 , n43795 , n43796 );
and ( n43798 , n1383 , n29508 );
and ( n43799 , n1580 , n28406 );
xor ( n43800 , n43798 , n43799 );
and ( n43801 , n1694 , n27296 );
xor ( n43802 , n43800 , n43801 );
xor ( n43803 , n43797 , n43802 );
and ( n43804 , n1047 , n32999 );
and ( n43805 , n1164 , n31761 );
xor ( n43806 , n43804 , n43805 );
and ( n43807 , n1287 , n30629 );
xor ( n43808 , n43806 , n43807 );
xor ( n43809 , n43803 , n43808 );
xor ( n43810 , n43793 , n43809 );
and ( n43811 , n42610 , n42611 );
not ( n43812 , n925 );
and ( n43813 , n34193 , n925 );
nor ( n43814 , n43812 , n43813 );
xor ( n43815 , n43811 , n43814 );
xor ( n43816 , n43810 , n43815 );
xor ( n43817 , n43787 , n43816 );
xor ( n43818 , n43738 , n43817 );
xor ( n43819 , n43655 , n43818 );
xor ( n43820 , n43530 , n43819 );
xor ( n43821 , n43448 , n43820 );
xor ( n43822 , n43439 , n43821 );
and ( n43823 , n42225 , n42228 );
and ( n43824 , n42228 , n42619 );
and ( n43825 , n42225 , n42619 );
or ( n43826 , n43823 , n43824 , n43825 );
xor ( n43827 , n43822 , n43826 );
and ( n43828 , n42620 , n42624 );
and ( n43829 , n42625 , n42628 );
or ( n43830 , n43828 , n43829 );
xor ( n43831 , n43827 , n43830 );
buf ( n43832 , n43831 );
buf ( n43833 , n43832 );
not ( n43834 , n43833 );
nor ( n43835 , n43834 , n8739 );
xor ( n43836 , n43431 , n43835 );
and ( n43837 , n42221 , n42633 );
and ( n43838 , n42634 , n42637 );
or ( n43839 , n43837 , n43838 );
xor ( n43840 , n43836 , n43839 );
buf ( n43841 , n43840 );
buf ( n43842 , n43841 );
not ( n43843 , n43842 );
buf ( n43844 , n570 );
not ( n43845 , n43844 );
nor ( n43846 , n43843 , n43845 );
xor ( n43847 , n43057 , n43846 );
xor ( n43848 , n42649 , n43054 );
nor ( n43849 , n42641 , n43845 );
and ( n43850 , n43848 , n43849 );
xor ( n43851 , n43848 , n43849 );
xor ( n43852 , n42653 , n43052 );
nor ( n43853 , n41437 , n43845 );
and ( n43854 , n43852 , n43853 );
xor ( n43855 , n43852 , n43853 );
xor ( n43856 , n42657 , n43050 );
nor ( n43857 , n40232 , n43845 );
and ( n43858 , n43856 , n43857 );
xor ( n43859 , n43856 , n43857 );
xor ( n43860 , n42661 , n43048 );
nor ( n43861 , n39027 , n43845 );
and ( n43862 , n43860 , n43861 );
xor ( n43863 , n43860 , n43861 );
xor ( n43864 , n42665 , n43046 );
nor ( n43865 , n37825 , n43845 );
and ( n43866 , n43864 , n43865 );
xor ( n43867 , n43864 , n43865 );
xor ( n43868 , n42669 , n43044 );
nor ( n43869 , n36620 , n43845 );
and ( n43870 , n43868 , n43869 );
xor ( n43871 , n43868 , n43869 );
xor ( n43872 , n42673 , n43042 );
nor ( n43873 , n35419 , n43845 );
and ( n43874 , n43872 , n43873 );
xor ( n43875 , n43872 , n43873 );
xor ( n43876 , n42677 , n43040 );
nor ( n43877 , n34224 , n43845 );
and ( n43878 , n43876 , n43877 );
xor ( n43879 , n43876 , n43877 );
xor ( n43880 , n42681 , n43038 );
nor ( n43881 , n33033 , n43845 );
and ( n43882 , n43880 , n43881 );
xor ( n43883 , n43880 , n43881 );
xor ( n43884 , n42685 , n43036 );
nor ( n43885 , n31867 , n43845 );
and ( n43886 , n43884 , n43885 );
xor ( n43887 , n43884 , n43885 );
xor ( n43888 , n42689 , n43034 );
nor ( n43889 , n30725 , n43845 );
and ( n43890 , n43888 , n43889 );
xor ( n43891 , n43888 , n43889 );
xor ( n43892 , n42693 , n43032 );
nor ( n43893 , n29596 , n43845 );
and ( n43894 , n43892 , n43893 );
xor ( n43895 , n43892 , n43893 );
xor ( n43896 , n42697 , n43030 );
nor ( n43897 , n28487 , n43845 );
and ( n43898 , n43896 , n43897 );
xor ( n43899 , n43896 , n43897 );
xor ( n43900 , n42701 , n43028 );
nor ( n43901 , n27397 , n43845 );
and ( n43902 , n43900 , n43901 );
xor ( n43903 , n43900 , n43901 );
xor ( n43904 , n42705 , n43026 );
nor ( n43905 , n26326 , n43845 );
and ( n43906 , n43904 , n43905 );
xor ( n43907 , n43904 , n43905 );
xor ( n43908 , n42709 , n43024 );
nor ( n43909 , n25272 , n43845 );
and ( n43910 , n43908 , n43909 );
xor ( n43911 , n43908 , n43909 );
xor ( n43912 , n42713 , n43022 );
nor ( n43913 , n24242 , n43845 );
and ( n43914 , n43912 , n43913 );
xor ( n43915 , n43912 , n43913 );
xor ( n43916 , n42717 , n43020 );
nor ( n43917 , n23225 , n43845 );
and ( n43918 , n43916 , n43917 );
xor ( n43919 , n43916 , n43917 );
xor ( n43920 , n42721 , n43018 );
nor ( n43921 , n22231 , n43845 );
and ( n43922 , n43920 , n43921 );
xor ( n43923 , n43920 , n43921 );
xor ( n43924 , n42725 , n43016 );
nor ( n43925 , n21258 , n43845 );
and ( n43926 , n43924 , n43925 );
xor ( n43927 , n43924 , n43925 );
xor ( n43928 , n42729 , n43014 );
nor ( n43929 , n20303 , n43845 );
and ( n43930 , n43928 , n43929 );
xor ( n43931 , n43928 , n43929 );
xor ( n43932 , n42733 , n43012 );
nor ( n43933 , n19365 , n43845 );
and ( n43934 , n43932 , n43933 );
xor ( n43935 , n43932 , n43933 );
xor ( n43936 , n42737 , n43010 );
nor ( n43937 , n18448 , n43845 );
and ( n43938 , n43936 , n43937 );
xor ( n43939 , n43936 , n43937 );
xor ( n43940 , n42741 , n43008 );
nor ( n43941 , n17548 , n43845 );
and ( n43942 , n43940 , n43941 );
xor ( n43943 , n43940 , n43941 );
xor ( n43944 , n42745 , n43006 );
nor ( n43945 , n16669 , n43845 );
and ( n43946 , n43944 , n43945 );
xor ( n43947 , n43944 , n43945 );
xor ( n43948 , n42749 , n43004 );
nor ( n43949 , n15809 , n43845 );
and ( n43950 , n43948 , n43949 );
xor ( n43951 , n43948 , n43949 );
xor ( n43952 , n42753 , n43002 );
nor ( n43953 , n14968 , n43845 );
and ( n43954 , n43952 , n43953 );
xor ( n43955 , n43952 , n43953 );
xor ( n43956 , n42757 , n43000 );
nor ( n43957 , n14147 , n43845 );
and ( n43958 , n43956 , n43957 );
xor ( n43959 , n43956 , n43957 );
xor ( n43960 , n42761 , n42998 );
nor ( n43961 , n13349 , n43845 );
and ( n43962 , n43960 , n43961 );
xor ( n43963 , n43960 , n43961 );
xor ( n43964 , n42765 , n42996 );
nor ( n43965 , n12564 , n43845 );
and ( n43966 , n43964 , n43965 );
xor ( n43967 , n43964 , n43965 );
xor ( n43968 , n42769 , n42994 );
nor ( n43969 , n11799 , n43845 );
and ( n43970 , n43968 , n43969 );
xor ( n43971 , n43968 , n43969 );
xor ( n43972 , n42773 , n42992 );
nor ( n43973 , n11050 , n43845 );
and ( n43974 , n43972 , n43973 );
xor ( n43975 , n43972 , n43973 );
xor ( n43976 , n42777 , n42990 );
nor ( n43977 , n10321 , n43845 );
and ( n43978 , n43976 , n43977 );
xor ( n43979 , n43976 , n43977 );
xor ( n43980 , n42781 , n42988 );
nor ( n43981 , n9429 , n43845 );
and ( n43982 , n43980 , n43981 );
xor ( n43983 , n43980 , n43981 );
xor ( n43984 , n42785 , n42986 );
nor ( n43985 , n8949 , n43845 );
and ( n43986 , n43984 , n43985 );
xor ( n43987 , n43984 , n43985 );
xor ( n43988 , n42789 , n42984 );
nor ( n43989 , n9437 , n43845 );
and ( n43990 , n43988 , n43989 );
xor ( n43991 , n43988 , n43989 );
xor ( n43992 , n42793 , n42982 );
nor ( n43993 , n9446 , n43845 );
and ( n43994 , n43992 , n43993 );
xor ( n43995 , n43992 , n43993 );
xor ( n43996 , n42797 , n42980 );
nor ( n43997 , n9455 , n43845 );
and ( n43998 , n43996 , n43997 );
xor ( n43999 , n43996 , n43997 );
xor ( n44000 , n42801 , n42978 );
nor ( n44001 , n9464 , n43845 );
and ( n44002 , n44000 , n44001 );
xor ( n44003 , n44000 , n44001 );
xor ( n44004 , n42805 , n42976 );
nor ( n44005 , n9473 , n43845 );
and ( n44006 , n44004 , n44005 );
xor ( n44007 , n44004 , n44005 );
xor ( n44008 , n42809 , n42974 );
nor ( n44009 , n9482 , n43845 );
and ( n44010 , n44008 , n44009 );
xor ( n44011 , n44008 , n44009 );
xor ( n44012 , n42813 , n42972 );
nor ( n44013 , n9491 , n43845 );
and ( n44014 , n44012 , n44013 );
xor ( n44015 , n44012 , n44013 );
xor ( n44016 , n42817 , n42970 );
nor ( n44017 , n9500 , n43845 );
and ( n44018 , n44016 , n44017 );
xor ( n44019 , n44016 , n44017 );
xor ( n44020 , n42821 , n42968 );
nor ( n44021 , n9509 , n43845 );
and ( n44022 , n44020 , n44021 );
xor ( n44023 , n44020 , n44021 );
xor ( n44024 , n42825 , n42966 );
nor ( n44025 , n9518 , n43845 );
and ( n44026 , n44024 , n44025 );
xor ( n44027 , n44024 , n44025 );
xor ( n44028 , n42829 , n42964 );
nor ( n44029 , n9527 , n43845 );
and ( n44030 , n44028 , n44029 );
xor ( n44031 , n44028 , n44029 );
xor ( n44032 , n42833 , n42962 );
nor ( n44033 , n9536 , n43845 );
and ( n44034 , n44032 , n44033 );
xor ( n44035 , n44032 , n44033 );
xor ( n44036 , n42837 , n42960 );
nor ( n44037 , n9545 , n43845 );
and ( n44038 , n44036 , n44037 );
xor ( n44039 , n44036 , n44037 );
xor ( n44040 , n42841 , n42958 );
nor ( n44041 , n9554 , n43845 );
and ( n44042 , n44040 , n44041 );
xor ( n44043 , n44040 , n44041 );
xor ( n44044 , n42845 , n42956 );
nor ( n44045 , n9563 , n43845 );
and ( n44046 , n44044 , n44045 );
xor ( n44047 , n44044 , n44045 );
xor ( n44048 , n42849 , n42954 );
nor ( n44049 , n9572 , n43845 );
and ( n44050 , n44048 , n44049 );
xor ( n44051 , n44048 , n44049 );
xor ( n44052 , n42853 , n42952 );
nor ( n44053 , n9581 , n43845 );
and ( n44054 , n44052 , n44053 );
xor ( n44055 , n44052 , n44053 );
xor ( n44056 , n42857 , n42950 );
nor ( n44057 , n9590 , n43845 );
and ( n44058 , n44056 , n44057 );
xor ( n44059 , n44056 , n44057 );
xor ( n44060 , n42861 , n42948 );
nor ( n44061 , n9599 , n43845 );
and ( n44062 , n44060 , n44061 );
xor ( n44063 , n44060 , n44061 );
xor ( n44064 , n42865 , n42946 );
nor ( n44065 , n9608 , n43845 );
and ( n44066 , n44064 , n44065 );
xor ( n44067 , n44064 , n44065 );
xor ( n44068 , n42869 , n42944 );
nor ( n44069 , n9617 , n43845 );
and ( n44070 , n44068 , n44069 );
xor ( n44071 , n44068 , n44069 );
xor ( n44072 , n42873 , n42942 );
nor ( n44073 , n9626 , n43845 );
and ( n44074 , n44072 , n44073 );
xor ( n44075 , n44072 , n44073 );
xor ( n44076 , n42877 , n42940 );
nor ( n44077 , n9635 , n43845 );
and ( n44078 , n44076 , n44077 );
xor ( n44079 , n44076 , n44077 );
xor ( n44080 , n42881 , n42938 );
nor ( n44081 , n9644 , n43845 );
and ( n44082 , n44080 , n44081 );
xor ( n44083 , n44080 , n44081 );
xor ( n44084 , n42885 , n42936 );
nor ( n44085 , n9653 , n43845 );
and ( n44086 , n44084 , n44085 );
xor ( n44087 , n44084 , n44085 );
xor ( n44088 , n42889 , n42934 );
nor ( n44089 , n9662 , n43845 );
and ( n44090 , n44088 , n44089 );
xor ( n44091 , n44088 , n44089 );
xor ( n44092 , n42893 , n42932 );
nor ( n44093 , n9671 , n43845 );
and ( n44094 , n44092 , n44093 );
xor ( n44095 , n44092 , n44093 );
xor ( n44096 , n42897 , n42930 );
nor ( n44097 , n9680 , n43845 );
and ( n44098 , n44096 , n44097 );
xor ( n44099 , n44096 , n44097 );
xor ( n44100 , n42901 , n42928 );
nor ( n44101 , n9689 , n43845 );
and ( n44102 , n44100 , n44101 );
xor ( n44103 , n44100 , n44101 );
xor ( n44104 , n42905 , n42926 );
nor ( n44105 , n9698 , n43845 );
and ( n44106 , n44104 , n44105 );
xor ( n44107 , n44104 , n44105 );
xor ( n44108 , n42909 , n42924 );
nor ( n44109 , n9707 , n43845 );
and ( n44110 , n44108 , n44109 );
xor ( n44111 , n44108 , n44109 );
xor ( n44112 , n42913 , n42922 );
nor ( n44113 , n9716 , n43845 );
and ( n44114 , n44112 , n44113 );
xor ( n44115 , n44112 , n44113 );
xor ( n44116 , n42917 , n42920 );
nor ( n44117 , n9725 , n43845 );
and ( n44118 , n44116 , n44117 );
xor ( n44119 , n44116 , n44117 );
xor ( n44120 , n42918 , n42919 );
nor ( n44121 , n9734 , n43845 );
and ( n44122 , n44120 , n44121 );
xor ( n44123 , n44120 , n44121 );
nor ( n44124 , n9752 , n42643 );
nor ( n44125 , n9743 , n43845 );
and ( n44126 , n44124 , n44125 );
and ( n44127 , n44123 , n44126 );
or ( n44128 , n44122 , n44127 );
and ( n44129 , n44119 , n44128 );
or ( n44130 , n44118 , n44129 );
and ( n44131 , n44115 , n44130 );
or ( n44132 , n44114 , n44131 );
and ( n44133 , n44111 , n44132 );
or ( n44134 , n44110 , n44133 );
and ( n44135 , n44107 , n44134 );
or ( n44136 , n44106 , n44135 );
and ( n44137 , n44103 , n44136 );
or ( n44138 , n44102 , n44137 );
and ( n44139 , n44099 , n44138 );
or ( n44140 , n44098 , n44139 );
and ( n44141 , n44095 , n44140 );
or ( n44142 , n44094 , n44141 );
and ( n44143 , n44091 , n44142 );
or ( n44144 , n44090 , n44143 );
and ( n44145 , n44087 , n44144 );
or ( n44146 , n44086 , n44145 );
and ( n44147 , n44083 , n44146 );
or ( n44148 , n44082 , n44147 );
and ( n44149 , n44079 , n44148 );
or ( n44150 , n44078 , n44149 );
and ( n44151 , n44075 , n44150 );
or ( n44152 , n44074 , n44151 );
and ( n44153 , n44071 , n44152 );
or ( n44154 , n44070 , n44153 );
and ( n44155 , n44067 , n44154 );
or ( n44156 , n44066 , n44155 );
and ( n44157 , n44063 , n44156 );
or ( n44158 , n44062 , n44157 );
and ( n44159 , n44059 , n44158 );
or ( n44160 , n44058 , n44159 );
and ( n44161 , n44055 , n44160 );
or ( n44162 , n44054 , n44161 );
and ( n44163 , n44051 , n44162 );
or ( n44164 , n44050 , n44163 );
and ( n44165 , n44047 , n44164 );
or ( n44166 , n44046 , n44165 );
and ( n44167 , n44043 , n44166 );
or ( n44168 , n44042 , n44167 );
and ( n44169 , n44039 , n44168 );
or ( n44170 , n44038 , n44169 );
and ( n44171 , n44035 , n44170 );
or ( n44172 , n44034 , n44171 );
and ( n44173 , n44031 , n44172 );
or ( n44174 , n44030 , n44173 );
and ( n44175 , n44027 , n44174 );
or ( n44176 , n44026 , n44175 );
and ( n44177 , n44023 , n44176 );
or ( n44178 , n44022 , n44177 );
and ( n44179 , n44019 , n44178 );
or ( n44180 , n44018 , n44179 );
and ( n44181 , n44015 , n44180 );
or ( n44182 , n44014 , n44181 );
and ( n44183 , n44011 , n44182 );
or ( n44184 , n44010 , n44183 );
and ( n44185 , n44007 , n44184 );
or ( n44186 , n44006 , n44185 );
and ( n44187 , n44003 , n44186 );
or ( n44188 , n44002 , n44187 );
and ( n44189 , n43999 , n44188 );
or ( n44190 , n43998 , n44189 );
and ( n44191 , n43995 , n44190 );
or ( n44192 , n43994 , n44191 );
and ( n44193 , n43991 , n44192 );
or ( n44194 , n43990 , n44193 );
and ( n44195 , n43987 , n44194 );
or ( n44196 , n43986 , n44195 );
and ( n44197 , n43983 , n44196 );
or ( n44198 , n43982 , n44197 );
and ( n44199 , n43979 , n44198 );
or ( n44200 , n43978 , n44199 );
and ( n44201 , n43975 , n44200 );
or ( n44202 , n43974 , n44201 );
and ( n44203 , n43971 , n44202 );
or ( n44204 , n43970 , n44203 );
and ( n44205 , n43967 , n44204 );
or ( n44206 , n43966 , n44205 );
and ( n44207 , n43963 , n44206 );
or ( n44208 , n43962 , n44207 );
and ( n44209 , n43959 , n44208 );
or ( n44210 , n43958 , n44209 );
and ( n44211 , n43955 , n44210 );
or ( n44212 , n43954 , n44211 );
and ( n44213 , n43951 , n44212 );
or ( n44214 , n43950 , n44213 );
and ( n44215 , n43947 , n44214 );
or ( n44216 , n43946 , n44215 );
and ( n44217 , n43943 , n44216 );
or ( n44218 , n43942 , n44217 );
and ( n44219 , n43939 , n44218 );
or ( n44220 , n43938 , n44219 );
and ( n44221 , n43935 , n44220 );
or ( n44222 , n43934 , n44221 );
and ( n44223 , n43931 , n44222 );
or ( n44224 , n43930 , n44223 );
and ( n44225 , n43927 , n44224 );
or ( n44226 , n43926 , n44225 );
and ( n44227 , n43923 , n44226 );
or ( n44228 , n43922 , n44227 );
and ( n44229 , n43919 , n44228 );
or ( n44230 , n43918 , n44229 );
and ( n44231 , n43915 , n44230 );
or ( n44232 , n43914 , n44231 );
and ( n44233 , n43911 , n44232 );
or ( n44234 , n43910 , n44233 );
and ( n44235 , n43907 , n44234 );
or ( n44236 , n43906 , n44235 );
and ( n44237 , n43903 , n44236 );
or ( n44238 , n43902 , n44237 );
and ( n44239 , n43899 , n44238 );
or ( n44240 , n43898 , n44239 );
and ( n44241 , n43895 , n44240 );
or ( n44242 , n43894 , n44241 );
and ( n44243 , n43891 , n44242 );
or ( n44244 , n43890 , n44243 );
and ( n44245 , n43887 , n44244 );
or ( n44246 , n43886 , n44245 );
and ( n44247 , n43883 , n44246 );
or ( n44248 , n43882 , n44247 );
and ( n44249 , n43879 , n44248 );
or ( n44250 , n43878 , n44249 );
and ( n44251 , n43875 , n44250 );
or ( n44252 , n43874 , n44251 );
and ( n44253 , n43871 , n44252 );
or ( n44254 , n43870 , n44253 );
and ( n44255 , n43867 , n44254 );
or ( n44256 , n43866 , n44255 );
and ( n44257 , n43863 , n44256 );
or ( n44258 , n43862 , n44257 );
and ( n44259 , n43859 , n44258 );
or ( n44260 , n43858 , n44259 );
and ( n44261 , n43855 , n44260 );
or ( n44262 , n43854 , n44261 );
and ( n44263 , n43851 , n44262 );
or ( n44264 , n43850 , n44263 );
xor ( n44265 , n43847 , n44264 );
and ( n44266 , n33403 , n1061 );
nor ( n44267 , n1062 , n44266 );
nor ( n44268 , n1176 , n32231 );
xor ( n44269 , n44267 , n44268 );
and ( n44270 , n43059 , n43060 );
and ( n44271 , n43061 , n43064 );
or ( n44272 , n44270 , n44271 );
xor ( n44273 , n44269 , n44272 );
nor ( n44274 , n1303 , n31083 );
xor ( n44275 , n44273 , n44274 );
and ( n44276 , n43065 , n43066 );
and ( n44277 , n43067 , n43070 );
or ( n44278 , n44276 , n44277 );
xor ( n44279 , n44275 , n44278 );
nor ( n44280 , n1445 , n29948 );
xor ( n44281 , n44279 , n44280 );
and ( n44282 , n43071 , n43072 );
and ( n44283 , n43073 , n43076 );
or ( n44284 , n44282 , n44283 );
xor ( n44285 , n44281 , n44284 );
nor ( n44286 , n1598 , n28833 );
xor ( n44287 , n44285 , n44286 );
and ( n44288 , n43077 , n43078 );
and ( n44289 , n43079 , n43082 );
or ( n44290 , n44288 , n44289 );
xor ( n44291 , n44287 , n44290 );
nor ( n44292 , n1766 , n27737 );
xor ( n44293 , n44291 , n44292 );
and ( n44294 , n43083 , n43084 );
and ( n44295 , n43085 , n43088 );
or ( n44296 , n44294 , n44295 );
xor ( n44297 , n44293 , n44296 );
nor ( n44298 , n1945 , n26660 );
xor ( n44299 , n44297 , n44298 );
and ( n44300 , n43089 , n43090 );
and ( n44301 , n43091 , n43094 );
or ( n44302 , n44300 , n44301 );
xor ( n44303 , n44299 , n44302 );
nor ( n44304 , n2137 , n25600 );
xor ( n44305 , n44303 , n44304 );
and ( n44306 , n43095 , n43096 );
and ( n44307 , n43097 , n43100 );
or ( n44308 , n44306 , n44307 );
xor ( n44309 , n44305 , n44308 );
nor ( n44310 , n2343 , n24564 );
xor ( n44311 , n44309 , n44310 );
and ( n44312 , n43101 , n43102 );
and ( n44313 , n43103 , n43106 );
or ( n44314 , n44312 , n44313 );
xor ( n44315 , n44311 , n44314 );
nor ( n44316 , n2566 , n23541 );
xor ( n44317 , n44315 , n44316 );
and ( n44318 , n43107 , n43108 );
and ( n44319 , n43109 , n43112 );
or ( n44320 , n44318 , n44319 );
xor ( n44321 , n44317 , n44320 );
nor ( n44322 , n2797 , n22541 );
xor ( n44323 , n44321 , n44322 );
and ( n44324 , n43113 , n43114 );
and ( n44325 , n43115 , n43118 );
or ( n44326 , n44324 , n44325 );
xor ( n44327 , n44323 , n44326 );
nor ( n44328 , n3043 , n21562 );
xor ( n44329 , n44327 , n44328 );
and ( n44330 , n43119 , n43120 );
and ( n44331 , n43121 , n43124 );
or ( n44332 , n44330 , n44331 );
xor ( n44333 , n44329 , n44332 );
nor ( n44334 , n3300 , n20601 );
xor ( n44335 , n44333 , n44334 );
and ( n44336 , n43125 , n43126 );
and ( n44337 , n43127 , n43130 );
or ( n44338 , n44336 , n44337 );
xor ( n44339 , n44335 , n44338 );
nor ( n44340 , n3570 , n19657 );
xor ( n44341 , n44339 , n44340 );
and ( n44342 , n43131 , n43132 );
and ( n44343 , n43133 , n43136 );
or ( n44344 , n44342 , n44343 );
xor ( n44345 , n44341 , n44344 );
nor ( n44346 , n3853 , n18734 );
xor ( n44347 , n44345 , n44346 );
and ( n44348 , n43137 , n43138 );
and ( n44349 , n43139 , n43142 );
or ( n44350 , n44348 , n44349 );
xor ( n44351 , n44347 , n44350 );
nor ( n44352 , n4151 , n17828 );
xor ( n44353 , n44351 , n44352 );
and ( n44354 , n43143 , n43144 );
and ( n44355 , n43145 , n43148 );
or ( n44356 , n44354 , n44355 );
xor ( n44357 , n44353 , n44356 );
nor ( n44358 , n4458 , n16943 );
xor ( n44359 , n44357 , n44358 );
and ( n44360 , n43149 , n43150 );
and ( n44361 , n43151 , n43154 );
or ( n44362 , n44360 , n44361 );
xor ( n44363 , n44359 , n44362 );
nor ( n44364 , n4786 , n16077 );
xor ( n44365 , n44363 , n44364 );
and ( n44366 , n43155 , n43156 );
and ( n44367 , n43157 , n43160 );
or ( n44368 , n44366 , n44367 );
xor ( n44369 , n44365 , n44368 );
nor ( n44370 , n5126 , n15230 );
xor ( n44371 , n44369 , n44370 );
and ( n44372 , n43161 , n43162 );
and ( n44373 , n43163 , n43166 );
or ( n44374 , n44372 , n44373 );
xor ( n44375 , n44371 , n44374 );
nor ( n44376 , n5477 , n14403 );
xor ( n44377 , n44375 , n44376 );
and ( n44378 , n43167 , n43168 );
and ( n44379 , n43169 , n43172 );
or ( n44380 , n44378 , n44379 );
xor ( n44381 , n44377 , n44380 );
nor ( n44382 , n5838 , n13599 );
xor ( n44383 , n44381 , n44382 );
and ( n44384 , n43173 , n43174 );
and ( n44385 , n43175 , n43178 );
or ( n44386 , n44384 , n44385 );
xor ( n44387 , n44383 , n44386 );
nor ( n44388 , n6212 , n12808 );
xor ( n44389 , n44387 , n44388 );
and ( n44390 , n43179 , n43180 );
and ( n44391 , n43181 , n43184 );
or ( n44392 , n44390 , n44391 );
xor ( n44393 , n44389 , n44392 );
nor ( n44394 , n6596 , n12037 );
xor ( n44395 , n44393 , n44394 );
and ( n44396 , n43185 , n43186 );
and ( n44397 , n43187 , n43190 );
or ( n44398 , n44396 , n44397 );
xor ( n44399 , n44395 , n44398 );
nor ( n44400 , n6997 , n11282 );
xor ( n44401 , n44399 , n44400 );
and ( n44402 , n43191 , n43192 );
and ( n44403 , n43193 , n43196 );
or ( n44404 , n44402 , n44403 );
xor ( n44405 , n44401 , n44404 );
nor ( n44406 , n7413 , n10547 );
xor ( n44407 , n44405 , n44406 );
and ( n44408 , n43197 , n43198 );
and ( n44409 , n43199 , n43202 );
or ( n44410 , n44408 , n44409 );
xor ( n44411 , n44407 , n44410 );
nor ( n44412 , n7841 , n9829 );
xor ( n44413 , n44411 , n44412 );
and ( n44414 , n43203 , n43204 );
and ( n44415 , n43205 , n43208 );
or ( n44416 , n44414 , n44415 );
xor ( n44417 , n44413 , n44416 );
nor ( n44418 , n8281 , n8955 );
xor ( n44419 , n44417 , n44418 );
and ( n44420 , n43209 , n43210 );
and ( n44421 , n43211 , n43214 );
or ( n44422 , n44420 , n44421 );
xor ( n44423 , n44419 , n44422 );
nor ( n44424 , n8737 , n603 );
xor ( n44425 , n44423 , n44424 );
and ( n44426 , n43215 , n43216 );
and ( n44427 , n43217 , n43220 );
or ( n44428 , n44426 , n44427 );
xor ( n44429 , n44425 , n44428 );
nor ( n44430 , n9420 , n652 );
xor ( n44431 , n44429 , n44430 );
and ( n44432 , n43221 , n43222 );
and ( n44433 , n43223 , n43226 );
or ( n44434 , n44432 , n44433 );
xor ( n44435 , n44431 , n44434 );
nor ( n44436 , n10312 , n624 );
xor ( n44437 , n44435 , n44436 );
and ( n44438 , n43227 , n43228 );
and ( n44439 , n43229 , n43232 );
or ( n44440 , n44438 , n44439 );
xor ( n44441 , n44437 , n44440 );
nor ( n44442 , n11041 , n648 );
xor ( n44443 , n44441 , n44442 );
and ( n44444 , n43233 , n43234 );
and ( n44445 , n43235 , n43238 );
or ( n44446 , n44444 , n44445 );
xor ( n44447 , n44443 , n44446 );
nor ( n44448 , n11790 , n686 );
xor ( n44449 , n44447 , n44448 );
and ( n44450 , n43239 , n43240 );
and ( n44451 , n43241 , n43244 );
or ( n44452 , n44450 , n44451 );
xor ( n44453 , n44449 , n44452 );
nor ( n44454 , n12555 , n735 );
xor ( n44455 , n44453 , n44454 );
and ( n44456 , n43245 , n43246 );
and ( n44457 , n43247 , n43250 );
or ( n44458 , n44456 , n44457 );
xor ( n44459 , n44455 , n44458 );
nor ( n44460 , n13340 , n798 );
xor ( n44461 , n44459 , n44460 );
and ( n44462 , n43251 , n43252 );
and ( n44463 , n43253 , n43256 );
or ( n44464 , n44462 , n44463 );
xor ( n44465 , n44461 , n44464 );
nor ( n44466 , n14138 , n870 );
xor ( n44467 , n44465 , n44466 );
and ( n44468 , n43257 , n43258 );
and ( n44469 , n43259 , n43262 );
or ( n44470 , n44468 , n44469 );
xor ( n44471 , n44467 , n44470 );
nor ( n44472 , n14959 , n960 );
xor ( n44473 , n44471 , n44472 );
and ( n44474 , n43263 , n43264 );
and ( n44475 , n43265 , n43268 );
or ( n44476 , n44474 , n44475 );
xor ( n44477 , n44473 , n44476 );
nor ( n44478 , n15800 , n1064 );
xor ( n44479 , n44477 , n44478 );
and ( n44480 , n43269 , n43270 );
and ( n44481 , n43271 , n43274 );
or ( n44482 , n44480 , n44481 );
xor ( n44483 , n44479 , n44482 );
nor ( n44484 , n16660 , n1178 );
xor ( n44485 , n44483 , n44484 );
and ( n44486 , n43275 , n43276 );
and ( n44487 , n43277 , n43280 );
or ( n44488 , n44486 , n44487 );
xor ( n44489 , n44485 , n44488 );
nor ( n44490 , n17539 , n1305 );
xor ( n44491 , n44489 , n44490 );
and ( n44492 , n43281 , n43282 );
and ( n44493 , n43283 , n43286 );
or ( n44494 , n44492 , n44493 );
xor ( n44495 , n44491 , n44494 );
nor ( n44496 , n18439 , n1447 );
xor ( n44497 , n44495 , n44496 );
and ( n44498 , n43287 , n43288 );
and ( n44499 , n43289 , n43292 );
or ( n44500 , n44498 , n44499 );
xor ( n44501 , n44497 , n44500 );
nor ( n44502 , n19356 , n1600 );
xor ( n44503 , n44501 , n44502 );
and ( n44504 , n43293 , n43294 );
and ( n44505 , n43295 , n43298 );
or ( n44506 , n44504 , n44505 );
xor ( n44507 , n44503 , n44506 );
nor ( n44508 , n20294 , n1768 );
xor ( n44509 , n44507 , n44508 );
and ( n44510 , n43299 , n43300 );
and ( n44511 , n43301 , n43304 );
or ( n44512 , n44510 , n44511 );
xor ( n44513 , n44509 , n44512 );
nor ( n44514 , n21249 , n1947 );
xor ( n44515 , n44513 , n44514 );
and ( n44516 , n43305 , n43306 );
and ( n44517 , n43307 , n43310 );
or ( n44518 , n44516 , n44517 );
xor ( n44519 , n44515 , n44518 );
nor ( n44520 , n22222 , n2139 );
xor ( n44521 , n44519 , n44520 );
and ( n44522 , n43311 , n43312 );
and ( n44523 , n43313 , n43316 );
or ( n44524 , n44522 , n44523 );
xor ( n44525 , n44521 , n44524 );
nor ( n44526 , n23216 , n2345 );
xor ( n44527 , n44525 , n44526 );
and ( n44528 , n43317 , n43318 );
and ( n44529 , n43319 , n43322 );
or ( n44530 , n44528 , n44529 );
xor ( n44531 , n44527 , n44530 );
nor ( n44532 , n24233 , n2568 );
xor ( n44533 , n44531 , n44532 );
and ( n44534 , n43323 , n43324 );
and ( n44535 , n43325 , n43328 );
or ( n44536 , n44534 , n44535 );
xor ( n44537 , n44533 , n44536 );
nor ( n44538 , n25263 , n2799 );
xor ( n44539 , n44537 , n44538 );
and ( n44540 , n43329 , n43330 );
and ( n44541 , n43331 , n43334 );
or ( n44542 , n44540 , n44541 );
xor ( n44543 , n44539 , n44542 );
nor ( n44544 , n26317 , n3045 );
xor ( n44545 , n44543 , n44544 );
and ( n44546 , n43335 , n43336 );
and ( n44547 , n43337 , n43340 );
or ( n44548 , n44546 , n44547 );
xor ( n44549 , n44545 , n44548 );
nor ( n44550 , n27388 , n3302 );
xor ( n44551 , n44549 , n44550 );
and ( n44552 , n43341 , n43342 );
and ( n44553 , n43343 , n43346 );
or ( n44554 , n44552 , n44553 );
xor ( n44555 , n44551 , n44554 );
nor ( n44556 , n28478 , n3572 );
xor ( n44557 , n44555 , n44556 );
and ( n44558 , n43347 , n43348 );
and ( n44559 , n43349 , n43352 );
or ( n44560 , n44558 , n44559 );
xor ( n44561 , n44557 , n44560 );
nor ( n44562 , n29587 , n3855 );
xor ( n44563 , n44561 , n44562 );
and ( n44564 , n43353 , n43354 );
and ( n44565 , n43355 , n43358 );
or ( n44566 , n44564 , n44565 );
xor ( n44567 , n44563 , n44566 );
nor ( n44568 , n30716 , n4153 );
xor ( n44569 , n44567 , n44568 );
and ( n44570 , n43359 , n43360 );
and ( n44571 , n43361 , n43364 );
or ( n44572 , n44570 , n44571 );
xor ( n44573 , n44569 , n44572 );
nor ( n44574 , n31858 , n4460 );
xor ( n44575 , n44573 , n44574 );
and ( n44576 , n43365 , n43366 );
and ( n44577 , n43367 , n43370 );
or ( n44578 , n44576 , n44577 );
xor ( n44579 , n44575 , n44578 );
nor ( n44580 , n33024 , n4788 );
xor ( n44581 , n44579 , n44580 );
and ( n44582 , n43371 , n43372 );
and ( n44583 , n43373 , n43376 );
or ( n44584 , n44582 , n44583 );
xor ( n44585 , n44581 , n44584 );
nor ( n44586 , n34215 , n5128 );
xor ( n44587 , n44585 , n44586 );
and ( n44588 , n43377 , n43378 );
and ( n44589 , n43379 , n43382 );
or ( n44590 , n44588 , n44589 );
xor ( n44591 , n44587 , n44590 );
nor ( n44592 , n35410 , n5479 );
xor ( n44593 , n44591 , n44592 );
and ( n44594 , n43383 , n43384 );
and ( n44595 , n43385 , n43388 );
or ( n44596 , n44594 , n44595 );
xor ( n44597 , n44593 , n44596 );
nor ( n44598 , n36611 , n5840 );
xor ( n44599 , n44597 , n44598 );
and ( n44600 , n43389 , n43390 );
and ( n44601 , n43391 , n43394 );
or ( n44602 , n44600 , n44601 );
xor ( n44603 , n44599 , n44602 );
nor ( n44604 , n37816 , n6214 );
xor ( n44605 , n44603 , n44604 );
and ( n44606 , n43395 , n43396 );
and ( n44607 , n43397 , n43400 );
or ( n44608 , n44606 , n44607 );
xor ( n44609 , n44605 , n44608 );
nor ( n44610 , n39018 , n6598 );
xor ( n44611 , n44609 , n44610 );
and ( n44612 , n43401 , n43402 );
and ( n44613 , n43403 , n43406 );
or ( n44614 , n44612 , n44613 );
xor ( n44615 , n44611 , n44614 );
nor ( n44616 , n40223 , n6999 );
xor ( n44617 , n44615 , n44616 );
and ( n44618 , n43407 , n43408 );
and ( n44619 , n43409 , n43412 );
or ( n44620 , n44618 , n44619 );
xor ( n44621 , n44617 , n44620 );
nor ( n44622 , n41428 , n7415 );
xor ( n44623 , n44621 , n44622 );
and ( n44624 , n43413 , n43414 );
and ( n44625 , n43415 , n43418 );
or ( n44626 , n44624 , n44625 );
xor ( n44627 , n44623 , n44626 );
nor ( n44628 , n42632 , n7843 );
xor ( n44629 , n44627 , n44628 );
and ( n44630 , n43419 , n43420 );
and ( n44631 , n43421 , n43424 );
or ( n44632 , n44630 , n44631 );
xor ( n44633 , n44629 , n44632 );
nor ( n44634 , n43834 , n8283 );
xor ( n44635 , n44633 , n44634 );
and ( n44636 , n43425 , n43426 );
and ( n44637 , n43427 , n43430 );
or ( n44638 , n44636 , n44637 );
xor ( n44639 , n44635 , n44638 );
and ( n44640 , n43443 , n43447 );
and ( n44641 , n43447 , n43820 );
and ( n44642 , n43443 , n43820 );
or ( n44643 , n44640 , n44641 , n44642 );
and ( n44644 , n33774 , n1034 );
not ( n44645 , n1034 );
nor ( n44646 , n44644 , n44645 );
xor ( n44647 , n44643 , n44646 );
and ( n44648 , n43456 , n43460 );
and ( n44649 , n43460 , n43528 );
and ( n44650 , n43456 , n43528 );
or ( n44651 , n44648 , n44649 , n44650 );
and ( n44652 , n43452 , n43529 );
and ( n44653 , n43529 , n43819 );
and ( n44654 , n43452 , n43819 );
or ( n44655 , n44652 , n44653 , n44654 );
xor ( n44656 , n44651 , n44655 );
and ( n44657 , n43534 , n43654 );
and ( n44658 , n43654 , n43818 );
and ( n44659 , n43534 , n43818 );
or ( n44660 , n44657 , n44658 , n44659 );
and ( n44661 , n43465 , n43469 );
and ( n44662 , n43469 , n43527 );
and ( n44663 , n43465 , n43527 );
or ( n44664 , n44661 , n44662 , n44663 );
and ( n44665 , n43538 , n43542 );
and ( n44666 , n43542 , n43653 );
and ( n44667 , n43538 , n43653 );
or ( n44668 , n44665 , n44666 , n44667 );
xor ( n44669 , n44664 , n44668 );
and ( n44670 , n43496 , n43500 );
and ( n44671 , n43500 , n43506 );
and ( n44672 , n43496 , n43506 );
or ( n44673 , n44670 , n44671 , n44672 );
and ( n44674 , n43474 , n43478 );
and ( n44675 , n43478 , n43526 );
and ( n44676 , n43474 , n43526 );
or ( n44677 , n44674 , n44675 , n44676 );
xor ( n44678 , n44673 , n44677 );
and ( n44679 , n43483 , n43487 );
and ( n44680 , n43487 , n43525 );
and ( n44681 , n43483 , n43525 );
or ( n44682 , n44679 , n44680 , n44681 );
and ( n44683 , n43551 , n43576 );
and ( n44684 , n43576 , n43614 );
and ( n44685 , n43551 , n43614 );
or ( n44686 , n44683 , n44684 , n44685 );
xor ( n44687 , n44682 , n44686 );
and ( n44688 , n43492 , n43507 );
and ( n44689 , n43507 , n43524 );
and ( n44690 , n43492 , n43524 );
or ( n44691 , n44688 , n44689 , n44690 );
and ( n44692 , n43555 , n43559 );
and ( n44693 , n43559 , n43575 );
and ( n44694 , n43555 , n43575 );
or ( n44695 , n44692 , n44693 , n44694 );
xor ( n44696 , n44691 , n44695 );
and ( n44697 , n43512 , n43517 );
and ( n44698 , n43517 , n43523 );
and ( n44699 , n43512 , n43523 );
or ( n44700 , n44697 , n44698 , n44699 );
and ( n44701 , n43502 , n43503 );
and ( n44702 , n43503 , n43505 );
and ( n44703 , n43502 , n43505 );
or ( n44704 , n44701 , n44702 , n44703 );
and ( n44705 , n43513 , n43514 );
and ( n44706 , n43514 , n43516 );
and ( n44707 , n43513 , n43516 );
or ( n44708 , n44705 , n44706 , n44707 );
xor ( n44709 , n44704 , n44708 );
and ( n44710 , n30695 , n1424 );
and ( n44711 , n31836 , n1254 );
xor ( n44712 , n44710 , n44711 );
and ( n44713 , n32649 , n1134 );
xor ( n44714 , n44712 , n44713 );
xor ( n44715 , n44709 , n44714 );
xor ( n44716 , n44700 , n44715 );
and ( n44717 , n43519 , n43520 );
and ( n44718 , n43520 , n43522 );
and ( n44719 , n43519 , n43522 );
or ( n44720 , n44717 , n44718 , n44719 );
and ( n44721 , n27361 , n1882 );
and ( n44722 , n28456 , n1738 );
xor ( n44723 , n44721 , n44722 );
and ( n44724 , n29559 , n1551 );
xor ( n44725 , n44723 , n44724 );
xor ( n44726 , n44720 , n44725 );
and ( n44727 , n24214 , n2544 );
and ( n44728 , n25243 , n2298 );
xor ( n44729 , n44727 , n44728 );
and ( n44730 , n26296 , n2100 );
xor ( n44731 , n44729 , n44730 );
xor ( n44732 , n44726 , n44731 );
xor ( n44733 , n44716 , n44732 );
xor ( n44734 , n44696 , n44733 );
xor ( n44735 , n44687 , n44734 );
xor ( n44736 , n44678 , n44735 );
xor ( n44737 , n44669 , n44736 );
xor ( n44738 , n44660 , n44737 );
and ( n44739 , n43659 , n43737 );
and ( n44740 , n43737 , n43817 );
and ( n44741 , n43659 , n43817 );
or ( n44742 , n44739 , n44740 , n44741 );
and ( n44743 , n43547 , n43615 );
and ( n44744 , n43615 , n43652 );
and ( n44745 , n43547 , n43652 );
or ( n44746 , n44743 , n44744 , n44745 );
and ( n44747 , n43663 , n43667 );
and ( n44748 , n43667 , n43736 );
and ( n44749 , n43663 , n43736 );
or ( n44750 , n44747 , n44748 , n44749 );
xor ( n44751 , n44746 , n44750 );
and ( n44752 , n43620 , n43624 );
and ( n44753 , n43624 , n43651 );
and ( n44754 , n43620 , n43651 );
or ( n44755 , n44752 , n44753 , n44754 );
and ( n44756 , n43581 , n43597 );
and ( n44757 , n43597 , n43613 );
and ( n44758 , n43581 , n43613 );
or ( n44759 , n44756 , n44757 , n44758 );
and ( n44760 , n43564 , n43568 );
and ( n44761 , n43568 , n43574 );
and ( n44762 , n43564 , n43574 );
or ( n44763 , n44760 , n44761 , n44762 );
and ( n44764 , n43585 , n43590 );
and ( n44765 , n43590 , n43596 );
and ( n44766 , n43585 , n43596 );
or ( n44767 , n44764 , n44765 , n44766 );
xor ( n44768 , n44763 , n44767 );
and ( n44769 , n43570 , n43571 );
and ( n44770 , n43571 , n43573 );
and ( n44771 , n43570 , n43573 );
or ( n44772 , n44769 , n44770 , n44771 );
and ( n44773 , n43586 , n43587 );
and ( n44774 , n43587 , n43589 );
and ( n44775 , n43586 , n43589 );
or ( n44776 , n44773 , n44774 , n44775 );
xor ( n44777 , n44772 , n44776 );
and ( n44778 , n21216 , n3271 );
and ( n44779 , n22186 , n2981 );
xor ( n44780 , n44778 , n44779 );
and ( n44781 , n22892 , n2739 );
xor ( n44782 , n44780 , n44781 );
xor ( n44783 , n44777 , n44782 );
xor ( n44784 , n44768 , n44783 );
xor ( n44785 , n44759 , n44784 );
and ( n44786 , n43602 , n43606 );
and ( n44787 , n43606 , n43612 );
and ( n44788 , n43602 , n43612 );
or ( n44789 , n44786 , n44787 , n44788 );
and ( n44790 , n43592 , n43593 );
and ( n44791 , n43593 , n43595 );
and ( n44792 , n43592 , n43595 );
or ( n44793 , n44790 , n44791 , n44792 );
and ( n44794 , n18144 , n4102 );
and ( n44795 , n19324 , n3749 );
xor ( n44796 , n44794 , n44795 );
and ( n44797 , n20233 , n3495 );
xor ( n44798 , n44796 , n44797 );
xor ( n44799 , n44793 , n44798 );
and ( n44800 , n15758 , n5103 );
and ( n44801 , n16637 , n4730 );
xor ( n44802 , n44800 , n44801 );
and ( n44803 , n17512 , n4403 );
xor ( n44804 , n44802 , n44803 );
xor ( n44805 , n44799 , n44804 );
xor ( n44806 , n44789 , n44805 );
and ( n44807 , n43608 , n43609 );
and ( n44808 , n43609 , n43611 );
and ( n44809 , n43608 , n43611 );
or ( n44810 , n44807 , n44808 , n44809 );
and ( n44811 , n43639 , n43640 );
and ( n44812 , n43640 , n43642 );
and ( n44813 , n43639 , n43642 );
or ( n44814 , n44811 , n44812 , n44813 );
xor ( n44815 , n44810 , n44814 );
and ( n44816 , n13322 , n6132 );
and ( n44817 , n14118 , n5765 );
xor ( n44818 , n44816 , n44817 );
and ( n44819 , n14938 , n5408 );
xor ( n44820 , n44818 , n44819 );
xor ( n44821 , n44815 , n44820 );
xor ( n44822 , n44806 , n44821 );
xor ( n44823 , n44785 , n44822 );
xor ( n44824 , n44755 , n44823 );
and ( n44825 , n43629 , n43633 );
and ( n44826 , n43633 , n43650 );
and ( n44827 , n43629 , n43650 );
or ( n44828 , n44825 , n44826 , n44827 );
and ( n44829 , n43676 , n43691 );
and ( n44830 , n43691 , n43708 );
and ( n44831 , n43676 , n43708 );
or ( n44832 , n44829 , n44830 , n44831 );
xor ( n44833 , n44828 , n44832 );
and ( n44834 , n43638 , n43643 );
and ( n44835 , n43643 , n43649 );
and ( n44836 , n43638 , n43649 );
or ( n44837 , n44834 , n44835 , n44836 );
and ( n44838 , n43680 , n43684 );
and ( n44839 , n43684 , n43690 );
and ( n44840 , n43680 , n43690 );
or ( n44841 , n44838 , n44839 , n44840 );
xor ( n44842 , n44837 , n44841 );
and ( n44843 , n43645 , n43646 );
and ( n44844 , n43646 , n43648 );
and ( n44845 , n43645 , n43648 );
or ( n44846 , n44843 , n44844 , n44845 );
and ( n44847 , n11015 , n7310 );
and ( n44848 , n11769 , n6971 );
xor ( n44849 , n44847 , n44848 );
and ( n44850 , n12320 , n6504 );
xor ( n44851 , n44849 , n44850 );
xor ( n44852 , n44846 , n44851 );
buf ( n44853 , n8718 );
and ( n44854 , n9400 , n8243 );
xor ( n44855 , n44853 , n44854 );
and ( n44856 , n10291 , n7662 );
xor ( n44857 , n44855 , n44856 );
xor ( n44858 , n44852 , n44857 );
xor ( n44859 , n44842 , n44858 );
xor ( n44860 , n44833 , n44859 );
xor ( n44861 , n44824 , n44860 );
xor ( n44862 , n44751 , n44861 );
xor ( n44863 , n44742 , n44862 );
and ( n44864 , n43739 , n43786 );
and ( n44865 , n43786 , n43816 );
and ( n44866 , n43739 , n43816 );
or ( n44867 , n44864 , n44865 , n44866 );
and ( n44868 , n43672 , n43709 );
and ( n44869 , n43709 , n43735 );
and ( n44870 , n43672 , n43735 );
or ( n44871 , n44868 , n44869 , n44870 );
and ( n44872 , n43743 , n43747 );
and ( n44873 , n43747 , n43785 );
and ( n44874 , n43743 , n43785 );
or ( n44875 , n44872 , n44873 , n44874 );
xor ( n44876 , n44871 , n44875 );
and ( n44877 , n43714 , n43718 );
and ( n44878 , n43718 , n43734 );
and ( n44879 , n43714 , n43734 );
or ( n44880 , n44877 , n44878 , n44879 );
and ( n44881 , n43696 , n43701 );
and ( n44882 , n43701 , n43707 );
and ( n44883 , n43696 , n43707 );
or ( n44884 , n44881 , n44882 , n44883 );
and ( n44885 , n43686 , n43687 );
and ( n44886 , n43687 , n43689 );
and ( n44887 , n43686 , n43689 );
or ( n44888 , n44885 , n44886 , n44887 );
and ( n44889 , n43697 , n43698 );
and ( n44890 , n43698 , n43700 );
and ( n44891 , n43697 , n43700 );
or ( n44892 , n44889 , n44890 , n44891 );
xor ( n44893 , n44888 , n44892 );
and ( n44894 , n7385 , n10977 );
and ( n44895 , n7808 , n10239 );
xor ( n44896 , n44894 , n44895 );
and ( n44897 , n8079 , n9348 );
xor ( n44898 , n44896 , n44897 );
xor ( n44899 , n44893 , n44898 );
xor ( n44900 , n44884 , n44899 );
and ( n44901 , n43703 , n43704 );
and ( n44902 , n43704 , n43706 );
and ( n44903 , n43703 , n43706 );
or ( n44904 , n44901 , n44902 , n44903 );
and ( n44905 , n6187 , n13256 );
and ( n44906 , n6569 , n12531 );
xor ( n44907 , n44905 , n44906 );
and ( n44908 , n6816 , n11718 );
xor ( n44909 , n44907 , n44908 );
xor ( n44910 , n44904 , n44909 );
and ( n44911 , n4959 , n15691 );
and ( n44912 , n5459 , n14838 );
xor ( n44913 , n44911 , n44912 );
and ( n44914 , n5819 , n14044 );
xor ( n44915 , n44913 , n44914 );
xor ( n44916 , n44910 , n44915 );
xor ( n44917 , n44900 , n44916 );
xor ( n44918 , n44880 , n44917 );
and ( n44919 , n43723 , n43727 );
and ( n44920 , n43727 , n43733 );
and ( n44921 , n43723 , n43733 );
or ( n44922 , n44919 , n44920 , n44921 );
and ( n44923 , n43756 , n43761 );
and ( n44924 , n43761 , n43767 );
and ( n44925 , n43756 , n43767 );
or ( n44926 , n44923 , n44924 , n44925 );
xor ( n44927 , n44922 , n44926 );
and ( n44928 , n43729 , n43730 );
and ( n44929 , n43730 , n43732 );
and ( n44930 , n43729 , n43732 );
or ( n44931 , n44928 , n44929 , n44930 );
and ( n44932 , n43757 , n43758 );
and ( n44933 , n43758 , n43760 );
and ( n44934 , n43757 , n43760 );
or ( n44935 , n44932 , n44933 , n44934 );
xor ( n44936 , n44931 , n44935 );
and ( n44937 , n4132 , n18407 );
and ( n44938 , n4438 , n17422 );
xor ( n44939 , n44937 , n44938 );
and ( n44940 , n4766 , n16550 );
xor ( n44941 , n44939 , n44940 );
xor ( n44942 , n44936 , n44941 );
xor ( n44943 , n44927 , n44942 );
xor ( n44944 , n44918 , n44943 );
xor ( n44945 , n44876 , n44944 );
xor ( n44946 , n44867 , n44945 );
and ( n44947 , n43810 , n43815 );
and ( n44948 , n43797 , n43802 );
and ( n44949 , n43802 , n43808 );
and ( n44950 , n43797 , n43808 );
or ( n44951 , n44948 , n44949 , n44950 );
and ( n44952 , n43811 , n43814 );
xor ( n44953 , n44951 , n44952 );
and ( n44954 , n43804 , n43805 );
and ( n44955 , n43805 , n43807 );
and ( n44956 , n43804 , n43807 );
or ( n44957 , n44954 , n44955 , n44956 );
and ( n44958 , n1383 , n30629 );
and ( n44959 , n1580 , n29508 );
xor ( n44960 , n44958 , n44959 );
and ( n44961 , n1694 , n28406 );
xor ( n44962 , n44960 , n44961 );
xor ( n44963 , n44957 , n44962 );
not ( n44964 , n1047 );
and ( n44965 , n34193 , n1047 );
nor ( n44966 , n44964 , n44965 );
and ( n44967 , n1164 , n32999 );
xor ( n44968 , n44966 , n44967 );
and ( n44969 , n1287 , n31761 );
xor ( n44970 , n44968 , n44969 );
xor ( n44971 , n44963 , n44970 );
xor ( n44972 , n44953 , n44971 );
xor ( n44973 , n44947 , n44972 );
and ( n44974 , n43791 , n43792 );
and ( n44975 , n43792 , n43809 );
and ( n44976 , n43791 , n43809 );
or ( n44977 , n44974 , n44975 , n44976 );
and ( n44978 , n43752 , n43768 );
and ( n44979 , n43768 , n43784 );
and ( n44980 , n43752 , n43784 );
or ( n44981 , n44978 , n44979 , n44980 );
xor ( n44982 , n44977 , n44981 );
and ( n44983 , n43773 , n43777 );
and ( n44984 , n43777 , n43783 );
and ( n44985 , n43773 , n43783 );
or ( n44986 , n44983 , n44984 , n44985 );
and ( n44987 , n43763 , n43764 );
and ( n44988 , n43764 , n43766 );
and ( n44989 , n43763 , n43766 );
or ( n44990 , n44987 , n44988 , n44989 );
and ( n44991 , n3182 , n20976 );
and ( n44992 , n3545 , n20156 );
xor ( n44993 , n44991 , n44992 );
and ( n44994 , n3801 , n19222 );
xor ( n44995 , n44993 , n44994 );
xor ( n44996 , n44990 , n44995 );
and ( n44997 , n2462 , n24137 );
and ( n44998 , n2779 , n23075 );
xor ( n44999 , n44997 , n44998 );
and ( n45000 , n3024 , n22065 );
xor ( n45001 , n44999 , n45000 );
xor ( n45002 , n44996 , n45001 );
xor ( n45003 , n44986 , n45002 );
and ( n45004 , n43779 , n43780 );
and ( n45005 , n43780 , n43782 );
and ( n45006 , n43779 , n43782 );
or ( n45007 , n45004 , n45005 , n45006 );
and ( n45008 , n43798 , n43799 );
and ( n45009 , n43799 , n43801 );
and ( n45010 , n43798 , n43801 );
or ( n45011 , n45008 , n45009 , n45010 );
xor ( n45012 , n45007 , n45011 );
and ( n45013 , n1933 , n27296 );
and ( n45014 , n2120 , n26216 );
xor ( n45015 , n45013 , n45014 );
and ( n45016 , n2324 , n25163 );
xor ( n45017 , n45015 , n45016 );
xor ( n45018 , n45012 , n45017 );
xor ( n45019 , n45003 , n45018 );
xor ( n45020 , n44982 , n45019 );
xor ( n45021 , n44973 , n45020 );
xor ( n45022 , n44946 , n45021 );
xor ( n45023 , n44863 , n45022 );
xor ( n45024 , n44738 , n45023 );
xor ( n45025 , n44656 , n45024 );
xor ( n45026 , n44647 , n45025 );
and ( n45027 , n43435 , n43438 );
and ( n45028 , n43438 , n43821 );
and ( n45029 , n43435 , n43821 );
or ( n45030 , n45027 , n45028 , n45029 );
xor ( n45031 , n45026 , n45030 );
and ( n45032 , n43822 , n43826 );
and ( n45033 , n43827 , n43830 );
or ( n45034 , n45032 , n45033 );
xor ( n45035 , n45031 , n45034 );
buf ( n45036 , n45035 );
buf ( n45037 , n45036 );
not ( n45038 , n45037 );
nor ( n45039 , n45038 , n8739 );
xor ( n45040 , n44639 , n45039 );
and ( n45041 , n43431 , n43835 );
and ( n45042 , n43836 , n43839 );
or ( n45043 , n45041 , n45042 );
xor ( n45044 , n45040 , n45043 );
buf ( n45045 , n45044 );
buf ( n45046 , n45045 );
not ( n45047 , n45046 );
buf ( n45048 , n571 );
not ( n45049 , n45048 );
nor ( n45050 , n45047 , n45049 );
xor ( n45051 , n44265 , n45050 );
xor ( n45052 , n43851 , n44262 );
nor ( n45053 , n43843 , n45049 );
and ( n45054 , n45052 , n45053 );
xor ( n45055 , n45052 , n45053 );
xor ( n45056 , n43855 , n44260 );
nor ( n45057 , n42641 , n45049 );
and ( n45058 , n45056 , n45057 );
xor ( n45059 , n45056 , n45057 );
xor ( n45060 , n43859 , n44258 );
nor ( n45061 , n41437 , n45049 );
and ( n45062 , n45060 , n45061 );
xor ( n45063 , n45060 , n45061 );
xor ( n45064 , n43863 , n44256 );
nor ( n45065 , n40232 , n45049 );
and ( n45066 , n45064 , n45065 );
xor ( n45067 , n45064 , n45065 );
xor ( n45068 , n43867 , n44254 );
nor ( n45069 , n39027 , n45049 );
and ( n45070 , n45068 , n45069 );
xor ( n45071 , n45068 , n45069 );
xor ( n45072 , n43871 , n44252 );
nor ( n45073 , n37825 , n45049 );
and ( n45074 , n45072 , n45073 );
xor ( n45075 , n45072 , n45073 );
xor ( n45076 , n43875 , n44250 );
nor ( n45077 , n36620 , n45049 );
and ( n45078 , n45076 , n45077 );
xor ( n45079 , n45076 , n45077 );
xor ( n45080 , n43879 , n44248 );
nor ( n45081 , n35419 , n45049 );
and ( n45082 , n45080 , n45081 );
xor ( n45083 , n45080 , n45081 );
xor ( n45084 , n43883 , n44246 );
nor ( n45085 , n34224 , n45049 );
and ( n45086 , n45084 , n45085 );
xor ( n45087 , n45084 , n45085 );
xor ( n45088 , n43887 , n44244 );
nor ( n45089 , n33033 , n45049 );
and ( n45090 , n45088 , n45089 );
xor ( n45091 , n45088 , n45089 );
xor ( n45092 , n43891 , n44242 );
nor ( n45093 , n31867 , n45049 );
and ( n45094 , n45092 , n45093 );
xor ( n45095 , n45092 , n45093 );
xor ( n45096 , n43895 , n44240 );
nor ( n45097 , n30725 , n45049 );
and ( n45098 , n45096 , n45097 );
xor ( n45099 , n45096 , n45097 );
xor ( n45100 , n43899 , n44238 );
nor ( n45101 , n29596 , n45049 );
and ( n45102 , n45100 , n45101 );
xor ( n45103 , n45100 , n45101 );
xor ( n45104 , n43903 , n44236 );
nor ( n45105 , n28487 , n45049 );
and ( n45106 , n45104 , n45105 );
xor ( n45107 , n45104 , n45105 );
xor ( n45108 , n43907 , n44234 );
nor ( n45109 , n27397 , n45049 );
and ( n45110 , n45108 , n45109 );
xor ( n45111 , n45108 , n45109 );
xor ( n45112 , n43911 , n44232 );
nor ( n45113 , n26326 , n45049 );
and ( n45114 , n45112 , n45113 );
xor ( n45115 , n45112 , n45113 );
xor ( n45116 , n43915 , n44230 );
nor ( n45117 , n25272 , n45049 );
and ( n45118 , n45116 , n45117 );
xor ( n45119 , n45116 , n45117 );
xor ( n45120 , n43919 , n44228 );
nor ( n45121 , n24242 , n45049 );
and ( n45122 , n45120 , n45121 );
xor ( n45123 , n45120 , n45121 );
xor ( n45124 , n43923 , n44226 );
nor ( n45125 , n23225 , n45049 );
and ( n45126 , n45124 , n45125 );
xor ( n45127 , n45124 , n45125 );
xor ( n45128 , n43927 , n44224 );
nor ( n45129 , n22231 , n45049 );
and ( n45130 , n45128 , n45129 );
xor ( n45131 , n45128 , n45129 );
xor ( n45132 , n43931 , n44222 );
nor ( n45133 , n21258 , n45049 );
and ( n45134 , n45132 , n45133 );
xor ( n45135 , n45132 , n45133 );
xor ( n45136 , n43935 , n44220 );
nor ( n45137 , n20303 , n45049 );
and ( n45138 , n45136 , n45137 );
xor ( n45139 , n45136 , n45137 );
xor ( n45140 , n43939 , n44218 );
nor ( n45141 , n19365 , n45049 );
and ( n45142 , n45140 , n45141 );
xor ( n45143 , n45140 , n45141 );
xor ( n45144 , n43943 , n44216 );
nor ( n45145 , n18448 , n45049 );
and ( n45146 , n45144 , n45145 );
xor ( n45147 , n45144 , n45145 );
xor ( n45148 , n43947 , n44214 );
nor ( n45149 , n17548 , n45049 );
and ( n45150 , n45148 , n45149 );
xor ( n45151 , n45148 , n45149 );
xor ( n45152 , n43951 , n44212 );
nor ( n45153 , n16669 , n45049 );
and ( n45154 , n45152 , n45153 );
xor ( n45155 , n45152 , n45153 );
xor ( n45156 , n43955 , n44210 );
nor ( n45157 , n15809 , n45049 );
and ( n45158 , n45156 , n45157 );
xor ( n45159 , n45156 , n45157 );
xor ( n45160 , n43959 , n44208 );
nor ( n45161 , n14968 , n45049 );
and ( n45162 , n45160 , n45161 );
xor ( n45163 , n45160 , n45161 );
xor ( n45164 , n43963 , n44206 );
nor ( n45165 , n14147 , n45049 );
and ( n45166 , n45164 , n45165 );
xor ( n45167 , n45164 , n45165 );
xor ( n45168 , n43967 , n44204 );
nor ( n45169 , n13349 , n45049 );
and ( n45170 , n45168 , n45169 );
xor ( n45171 , n45168 , n45169 );
xor ( n45172 , n43971 , n44202 );
nor ( n45173 , n12564 , n45049 );
and ( n45174 , n45172 , n45173 );
xor ( n45175 , n45172 , n45173 );
xor ( n45176 , n43975 , n44200 );
nor ( n45177 , n11799 , n45049 );
and ( n45178 , n45176 , n45177 );
xor ( n45179 , n45176 , n45177 );
xor ( n45180 , n43979 , n44198 );
nor ( n45181 , n11050 , n45049 );
and ( n45182 , n45180 , n45181 );
xor ( n45183 , n45180 , n45181 );
xor ( n45184 , n43983 , n44196 );
nor ( n45185 , n10321 , n45049 );
and ( n45186 , n45184 , n45185 );
xor ( n45187 , n45184 , n45185 );
xor ( n45188 , n43987 , n44194 );
nor ( n45189 , n9429 , n45049 );
and ( n45190 , n45188 , n45189 );
xor ( n45191 , n45188 , n45189 );
xor ( n45192 , n43991 , n44192 );
nor ( n45193 , n8949 , n45049 );
and ( n45194 , n45192 , n45193 );
xor ( n45195 , n45192 , n45193 );
xor ( n45196 , n43995 , n44190 );
nor ( n45197 , n9437 , n45049 );
and ( n45198 , n45196 , n45197 );
xor ( n45199 , n45196 , n45197 );
xor ( n45200 , n43999 , n44188 );
nor ( n45201 , n9446 , n45049 );
and ( n45202 , n45200 , n45201 );
xor ( n45203 , n45200 , n45201 );
xor ( n45204 , n44003 , n44186 );
nor ( n45205 , n9455 , n45049 );
and ( n45206 , n45204 , n45205 );
xor ( n45207 , n45204 , n45205 );
xor ( n45208 , n44007 , n44184 );
nor ( n45209 , n9464 , n45049 );
and ( n45210 , n45208 , n45209 );
xor ( n45211 , n45208 , n45209 );
xor ( n45212 , n44011 , n44182 );
nor ( n45213 , n9473 , n45049 );
and ( n45214 , n45212 , n45213 );
xor ( n45215 , n45212 , n45213 );
xor ( n45216 , n44015 , n44180 );
nor ( n45217 , n9482 , n45049 );
and ( n45218 , n45216 , n45217 );
xor ( n45219 , n45216 , n45217 );
xor ( n45220 , n44019 , n44178 );
nor ( n45221 , n9491 , n45049 );
and ( n45222 , n45220 , n45221 );
xor ( n45223 , n45220 , n45221 );
xor ( n45224 , n44023 , n44176 );
nor ( n45225 , n9500 , n45049 );
and ( n45226 , n45224 , n45225 );
xor ( n45227 , n45224 , n45225 );
xor ( n45228 , n44027 , n44174 );
nor ( n45229 , n9509 , n45049 );
and ( n45230 , n45228 , n45229 );
xor ( n45231 , n45228 , n45229 );
xor ( n45232 , n44031 , n44172 );
nor ( n45233 , n9518 , n45049 );
and ( n45234 , n45232 , n45233 );
xor ( n45235 , n45232 , n45233 );
xor ( n45236 , n44035 , n44170 );
nor ( n45237 , n9527 , n45049 );
and ( n45238 , n45236 , n45237 );
xor ( n45239 , n45236 , n45237 );
xor ( n45240 , n44039 , n44168 );
nor ( n45241 , n9536 , n45049 );
and ( n45242 , n45240 , n45241 );
xor ( n45243 , n45240 , n45241 );
xor ( n45244 , n44043 , n44166 );
nor ( n45245 , n9545 , n45049 );
and ( n45246 , n45244 , n45245 );
xor ( n45247 , n45244 , n45245 );
xor ( n45248 , n44047 , n44164 );
nor ( n45249 , n9554 , n45049 );
and ( n45250 , n45248 , n45249 );
xor ( n45251 , n45248 , n45249 );
xor ( n45252 , n44051 , n44162 );
nor ( n45253 , n9563 , n45049 );
and ( n45254 , n45252 , n45253 );
xor ( n45255 , n45252 , n45253 );
xor ( n45256 , n44055 , n44160 );
nor ( n45257 , n9572 , n45049 );
and ( n45258 , n45256 , n45257 );
xor ( n45259 , n45256 , n45257 );
xor ( n45260 , n44059 , n44158 );
nor ( n45261 , n9581 , n45049 );
and ( n45262 , n45260 , n45261 );
xor ( n45263 , n45260 , n45261 );
xor ( n45264 , n44063 , n44156 );
nor ( n45265 , n9590 , n45049 );
and ( n45266 , n45264 , n45265 );
xor ( n45267 , n45264 , n45265 );
xor ( n45268 , n44067 , n44154 );
nor ( n45269 , n9599 , n45049 );
and ( n45270 , n45268 , n45269 );
xor ( n45271 , n45268 , n45269 );
xor ( n45272 , n44071 , n44152 );
nor ( n45273 , n9608 , n45049 );
and ( n45274 , n45272 , n45273 );
xor ( n45275 , n45272 , n45273 );
xor ( n45276 , n44075 , n44150 );
nor ( n45277 , n9617 , n45049 );
and ( n45278 , n45276 , n45277 );
xor ( n45279 , n45276 , n45277 );
xor ( n45280 , n44079 , n44148 );
nor ( n45281 , n9626 , n45049 );
and ( n45282 , n45280 , n45281 );
xor ( n45283 , n45280 , n45281 );
xor ( n45284 , n44083 , n44146 );
nor ( n45285 , n9635 , n45049 );
and ( n45286 , n45284 , n45285 );
xor ( n45287 , n45284 , n45285 );
xor ( n45288 , n44087 , n44144 );
nor ( n45289 , n9644 , n45049 );
and ( n45290 , n45288 , n45289 );
xor ( n45291 , n45288 , n45289 );
xor ( n45292 , n44091 , n44142 );
nor ( n45293 , n9653 , n45049 );
and ( n45294 , n45292 , n45293 );
xor ( n45295 , n45292 , n45293 );
xor ( n45296 , n44095 , n44140 );
nor ( n45297 , n9662 , n45049 );
and ( n45298 , n45296 , n45297 );
xor ( n45299 , n45296 , n45297 );
xor ( n45300 , n44099 , n44138 );
nor ( n45301 , n9671 , n45049 );
and ( n45302 , n45300 , n45301 );
xor ( n45303 , n45300 , n45301 );
xor ( n45304 , n44103 , n44136 );
nor ( n45305 , n9680 , n45049 );
and ( n45306 , n45304 , n45305 );
xor ( n45307 , n45304 , n45305 );
xor ( n45308 , n44107 , n44134 );
nor ( n45309 , n9689 , n45049 );
and ( n45310 , n45308 , n45309 );
xor ( n45311 , n45308 , n45309 );
xor ( n45312 , n44111 , n44132 );
nor ( n45313 , n9698 , n45049 );
and ( n45314 , n45312 , n45313 );
xor ( n45315 , n45312 , n45313 );
xor ( n45316 , n44115 , n44130 );
nor ( n45317 , n9707 , n45049 );
and ( n45318 , n45316 , n45317 );
xor ( n45319 , n45316 , n45317 );
xor ( n45320 , n44119 , n44128 );
nor ( n45321 , n9716 , n45049 );
and ( n45322 , n45320 , n45321 );
xor ( n45323 , n45320 , n45321 );
xor ( n45324 , n44123 , n44126 );
nor ( n45325 , n9725 , n45049 );
and ( n45326 , n45324 , n45325 );
xor ( n45327 , n45324 , n45325 );
xor ( n45328 , n44124 , n44125 );
nor ( n45329 , n9734 , n45049 );
and ( n45330 , n45328 , n45329 );
xor ( n45331 , n45328 , n45329 );
nor ( n45332 , n9752 , n43845 );
nor ( n45333 , n9743 , n45049 );
and ( n45334 , n45332 , n45333 );
and ( n45335 , n45331 , n45334 );
or ( n45336 , n45330 , n45335 );
and ( n45337 , n45327 , n45336 );
or ( n45338 , n45326 , n45337 );
and ( n45339 , n45323 , n45338 );
or ( n45340 , n45322 , n45339 );
and ( n45341 , n45319 , n45340 );
or ( n45342 , n45318 , n45341 );
and ( n45343 , n45315 , n45342 );
or ( n45344 , n45314 , n45343 );
and ( n45345 , n45311 , n45344 );
or ( n45346 , n45310 , n45345 );
and ( n45347 , n45307 , n45346 );
or ( n45348 , n45306 , n45347 );
and ( n45349 , n45303 , n45348 );
or ( n45350 , n45302 , n45349 );
and ( n45351 , n45299 , n45350 );
or ( n45352 , n45298 , n45351 );
and ( n45353 , n45295 , n45352 );
or ( n45354 , n45294 , n45353 );
and ( n45355 , n45291 , n45354 );
or ( n45356 , n45290 , n45355 );
and ( n45357 , n45287 , n45356 );
or ( n45358 , n45286 , n45357 );
and ( n45359 , n45283 , n45358 );
or ( n45360 , n45282 , n45359 );
and ( n45361 , n45279 , n45360 );
or ( n45362 , n45278 , n45361 );
and ( n45363 , n45275 , n45362 );
or ( n45364 , n45274 , n45363 );
and ( n45365 , n45271 , n45364 );
or ( n45366 , n45270 , n45365 );
and ( n45367 , n45267 , n45366 );
or ( n45368 , n45266 , n45367 );
and ( n45369 , n45263 , n45368 );
or ( n45370 , n45262 , n45369 );
and ( n45371 , n45259 , n45370 );
or ( n45372 , n45258 , n45371 );
and ( n45373 , n45255 , n45372 );
or ( n45374 , n45254 , n45373 );
and ( n45375 , n45251 , n45374 );
or ( n45376 , n45250 , n45375 );
and ( n45377 , n45247 , n45376 );
or ( n45378 , n45246 , n45377 );
and ( n45379 , n45243 , n45378 );
or ( n45380 , n45242 , n45379 );
and ( n45381 , n45239 , n45380 );
or ( n45382 , n45238 , n45381 );
and ( n45383 , n45235 , n45382 );
or ( n45384 , n45234 , n45383 );
and ( n45385 , n45231 , n45384 );
or ( n45386 , n45230 , n45385 );
and ( n45387 , n45227 , n45386 );
or ( n45388 , n45226 , n45387 );
and ( n45389 , n45223 , n45388 );
or ( n45390 , n45222 , n45389 );
and ( n45391 , n45219 , n45390 );
or ( n45392 , n45218 , n45391 );
and ( n45393 , n45215 , n45392 );
or ( n45394 , n45214 , n45393 );
and ( n45395 , n45211 , n45394 );
or ( n45396 , n45210 , n45395 );
and ( n45397 , n45207 , n45396 );
or ( n45398 , n45206 , n45397 );
and ( n45399 , n45203 , n45398 );
or ( n45400 , n45202 , n45399 );
and ( n45401 , n45199 , n45400 );
or ( n45402 , n45198 , n45401 );
and ( n45403 , n45195 , n45402 );
or ( n45404 , n45194 , n45403 );
and ( n45405 , n45191 , n45404 );
or ( n45406 , n45190 , n45405 );
and ( n45407 , n45187 , n45406 );
or ( n45408 , n45186 , n45407 );
and ( n45409 , n45183 , n45408 );
or ( n45410 , n45182 , n45409 );
and ( n45411 , n45179 , n45410 );
or ( n45412 , n45178 , n45411 );
and ( n45413 , n45175 , n45412 );
or ( n45414 , n45174 , n45413 );
and ( n45415 , n45171 , n45414 );
or ( n45416 , n45170 , n45415 );
and ( n45417 , n45167 , n45416 );
or ( n45418 , n45166 , n45417 );
and ( n45419 , n45163 , n45418 );
or ( n45420 , n45162 , n45419 );
and ( n45421 , n45159 , n45420 );
or ( n45422 , n45158 , n45421 );
and ( n45423 , n45155 , n45422 );
or ( n45424 , n45154 , n45423 );
and ( n45425 , n45151 , n45424 );
or ( n45426 , n45150 , n45425 );
and ( n45427 , n45147 , n45426 );
or ( n45428 , n45146 , n45427 );
and ( n45429 , n45143 , n45428 );
or ( n45430 , n45142 , n45429 );
and ( n45431 , n45139 , n45430 );
or ( n45432 , n45138 , n45431 );
and ( n45433 , n45135 , n45432 );
or ( n45434 , n45134 , n45433 );
and ( n45435 , n45131 , n45434 );
or ( n45436 , n45130 , n45435 );
and ( n45437 , n45127 , n45436 );
or ( n45438 , n45126 , n45437 );
and ( n45439 , n45123 , n45438 );
or ( n45440 , n45122 , n45439 );
and ( n45441 , n45119 , n45440 );
or ( n45442 , n45118 , n45441 );
and ( n45443 , n45115 , n45442 );
or ( n45444 , n45114 , n45443 );
and ( n45445 , n45111 , n45444 );
or ( n45446 , n45110 , n45445 );
and ( n45447 , n45107 , n45446 );
or ( n45448 , n45106 , n45447 );
and ( n45449 , n45103 , n45448 );
or ( n45450 , n45102 , n45449 );
and ( n45451 , n45099 , n45450 );
or ( n45452 , n45098 , n45451 );
and ( n45453 , n45095 , n45452 );
or ( n45454 , n45094 , n45453 );
and ( n45455 , n45091 , n45454 );
or ( n45456 , n45090 , n45455 );
and ( n45457 , n45087 , n45456 );
or ( n45458 , n45086 , n45457 );
and ( n45459 , n45083 , n45458 );
or ( n45460 , n45082 , n45459 );
and ( n45461 , n45079 , n45460 );
or ( n45462 , n45078 , n45461 );
and ( n45463 , n45075 , n45462 );
or ( n45464 , n45074 , n45463 );
and ( n45465 , n45071 , n45464 );
or ( n45466 , n45070 , n45465 );
and ( n45467 , n45067 , n45466 );
or ( n45468 , n45066 , n45467 );
and ( n45469 , n45063 , n45468 );
or ( n45470 , n45062 , n45469 );
and ( n45471 , n45059 , n45470 );
or ( n45472 , n45058 , n45471 );
and ( n45473 , n45055 , n45472 );
or ( n45474 , n45054 , n45473 );
xor ( n45475 , n45051 , n45474 );
and ( n45476 , n33403 , n1175 );
nor ( n45477 , n1176 , n45476 );
nor ( n45478 , n1303 , n32231 );
xor ( n45479 , n45477 , n45478 );
and ( n45480 , n44267 , n44268 );
and ( n45481 , n44269 , n44272 );
or ( n45482 , n45480 , n45481 );
xor ( n45483 , n45479 , n45482 );
nor ( n45484 , n1445 , n31083 );
xor ( n45485 , n45483 , n45484 );
and ( n45486 , n44273 , n44274 );
and ( n45487 , n44275 , n44278 );
or ( n45488 , n45486 , n45487 );
xor ( n45489 , n45485 , n45488 );
nor ( n45490 , n1598 , n29948 );
xor ( n45491 , n45489 , n45490 );
and ( n45492 , n44279 , n44280 );
and ( n45493 , n44281 , n44284 );
or ( n45494 , n45492 , n45493 );
xor ( n45495 , n45491 , n45494 );
nor ( n45496 , n1766 , n28833 );
xor ( n45497 , n45495 , n45496 );
and ( n45498 , n44285 , n44286 );
and ( n45499 , n44287 , n44290 );
or ( n45500 , n45498 , n45499 );
xor ( n45501 , n45497 , n45500 );
nor ( n45502 , n1945 , n27737 );
xor ( n45503 , n45501 , n45502 );
and ( n45504 , n44291 , n44292 );
and ( n45505 , n44293 , n44296 );
or ( n45506 , n45504 , n45505 );
xor ( n45507 , n45503 , n45506 );
nor ( n45508 , n2137 , n26660 );
xor ( n45509 , n45507 , n45508 );
and ( n45510 , n44297 , n44298 );
and ( n45511 , n44299 , n44302 );
or ( n45512 , n45510 , n45511 );
xor ( n45513 , n45509 , n45512 );
nor ( n45514 , n2343 , n25600 );
xor ( n45515 , n45513 , n45514 );
and ( n45516 , n44303 , n44304 );
and ( n45517 , n44305 , n44308 );
or ( n45518 , n45516 , n45517 );
xor ( n45519 , n45515 , n45518 );
nor ( n45520 , n2566 , n24564 );
xor ( n45521 , n45519 , n45520 );
and ( n45522 , n44309 , n44310 );
and ( n45523 , n44311 , n44314 );
or ( n45524 , n45522 , n45523 );
xor ( n45525 , n45521 , n45524 );
nor ( n45526 , n2797 , n23541 );
xor ( n45527 , n45525 , n45526 );
and ( n45528 , n44315 , n44316 );
and ( n45529 , n44317 , n44320 );
or ( n45530 , n45528 , n45529 );
xor ( n45531 , n45527 , n45530 );
nor ( n45532 , n3043 , n22541 );
xor ( n45533 , n45531 , n45532 );
and ( n45534 , n44321 , n44322 );
and ( n45535 , n44323 , n44326 );
or ( n45536 , n45534 , n45535 );
xor ( n45537 , n45533 , n45536 );
nor ( n45538 , n3300 , n21562 );
xor ( n45539 , n45537 , n45538 );
and ( n45540 , n44327 , n44328 );
and ( n45541 , n44329 , n44332 );
or ( n45542 , n45540 , n45541 );
xor ( n45543 , n45539 , n45542 );
nor ( n45544 , n3570 , n20601 );
xor ( n45545 , n45543 , n45544 );
and ( n45546 , n44333 , n44334 );
and ( n45547 , n44335 , n44338 );
or ( n45548 , n45546 , n45547 );
xor ( n45549 , n45545 , n45548 );
nor ( n45550 , n3853 , n19657 );
xor ( n45551 , n45549 , n45550 );
and ( n45552 , n44339 , n44340 );
and ( n45553 , n44341 , n44344 );
or ( n45554 , n45552 , n45553 );
xor ( n45555 , n45551 , n45554 );
nor ( n45556 , n4151 , n18734 );
xor ( n45557 , n45555 , n45556 );
and ( n45558 , n44345 , n44346 );
and ( n45559 , n44347 , n44350 );
or ( n45560 , n45558 , n45559 );
xor ( n45561 , n45557 , n45560 );
nor ( n45562 , n4458 , n17828 );
xor ( n45563 , n45561 , n45562 );
and ( n45564 , n44351 , n44352 );
and ( n45565 , n44353 , n44356 );
or ( n45566 , n45564 , n45565 );
xor ( n45567 , n45563 , n45566 );
nor ( n45568 , n4786 , n16943 );
xor ( n45569 , n45567 , n45568 );
and ( n45570 , n44357 , n44358 );
and ( n45571 , n44359 , n44362 );
or ( n45572 , n45570 , n45571 );
xor ( n45573 , n45569 , n45572 );
nor ( n45574 , n5126 , n16077 );
xor ( n45575 , n45573 , n45574 );
and ( n45576 , n44363 , n44364 );
and ( n45577 , n44365 , n44368 );
or ( n45578 , n45576 , n45577 );
xor ( n45579 , n45575 , n45578 );
nor ( n45580 , n5477 , n15230 );
xor ( n45581 , n45579 , n45580 );
and ( n45582 , n44369 , n44370 );
and ( n45583 , n44371 , n44374 );
or ( n45584 , n45582 , n45583 );
xor ( n45585 , n45581 , n45584 );
nor ( n45586 , n5838 , n14403 );
xor ( n45587 , n45585 , n45586 );
and ( n45588 , n44375 , n44376 );
and ( n45589 , n44377 , n44380 );
or ( n45590 , n45588 , n45589 );
xor ( n45591 , n45587 , n45590 );
nor ( n45592 , n6212 , n13599 );
xor ( n45593 , n45591 , n45592 );
and ( n45594 , n44381 , n44382 );
and ( n45595 , n44383 , n44386 );
or ( n45596 , n45594 , n45595 );
xor ( n45597 , n45593 , n45596 );
nor ( n45598 , n6596 , n12808 );
xor ( n45599 , n45597 , n45598 );
and ( n45600 , n44387 , n44388 );
and ( n45601 , n44389 , n44392 );
or ( n45602 , n45600 , n45601 );
xor ( n45603 , n45599 , n45602 );
nor ( n45604 , n6997 , n12037 );
xor ( n45605 , n45603 , n45604 );
and ( n45606 , n44393 , n44394 );
and ( n45607 , n44395 , n44398 );
or ( n45608 , n45606 , n45607 );
xor ( n45609 , n45605 , n45608 );
nor ( n45610 , n7413 , n11282 );
xor ( n45611 , n45609 , n45610 );
and ( n45612 , n44399 , n44400 );
and ( n45613 , n44401 , n44404 );
or ( n45614 , n45612 , n45613 );
xor ( n45615 , n45611 , n45614 );
nor ( n45616 , n7841 , n10547 );
xor ( n45617 , n45615 , n45616 );
and ( n45618 , n44405 , n44406 );
and ( n45619 , n44407 , n44410 );
or ( n45620 , n45618 , n45619 );
xor ( n45621 , n45617 , n45620 );
nor ( n45622 , n8281 , n9829 );
xor ( n45623 , n45621 , n45622 );
and ( n45624 , n44411 , n44412 );
and ( n45625 , n44413 , n44416 );
or ( n45626 , n45624 , n45625 );
xor ( n45627 , n45623 , n45626 );
nor ( n45628 , n8737 , n8955 );
xor ( n45629 , n45627 , n45628 );
and ( n45630 , n44417 , n44418 );
and ( n45631 , n44419 , n44422 );
or ( n45632 , n45630 , n45631 );
xor ( n45633 , n45629 , n45632 );
nor ( n45634 , n9420 , n603 );
xor ( n45635 , n45633 , n45634 );
and ( n45636 , n44423 , n44424 );
and ( n45637 , n44425 , n44428 );
or ( n45638 , n45636 , n45637 );
xor ( n45639 , n45635 , n45638 );
nor ( n45640 , n10312 , n652 );
xor ( n45641 , n45639 , n45640 );
and ( n45642 , n44429 , n44430 );
and ( n45643 , n44431 , n44434 );
or ( n45644 , n45642 , n45643 );
xor ( n45645 , n45641 , n45644 );
nor ( n45646 , n11041 , n624 );
xor ( n45647 , n45645 , n45646 );
and ( n45648 , n44435 , n44436 );
and ( n45649 , n44437 , n44440 );
or ( n45650 , n45648 , n45649 );
xor ( n45651 , n45647 , n45650 );
nor ( n45652 , n11790 , n648 );
xor ( n45653 , n45651 , n45652 );
and ( n45654 , n44441 , n44442 );
and ( n45655 , n44443 , n44446 );
or ( n45656 , n45654 , n45655 );
xor ( n45657 , n45653 , n45656 );
nor ( n45658 , n12555 , n686 );
xor ( n45659 , n45657 , n45658 );
and ( n45660 , n44447 , n44448 );
and ( n45661 , n44449 , n44452 );
or ( n45662 , n45660 , n45661 );
xor ( n45663 , n45659 , n45662 );
nor ( n45664 , n13340 , n735 );
xor ( n45665 , n45663 , n45664 );
and ( n45666 , n44453 , n44454 );
and ( n45667 , n44455 , n44458 );
or ( n45668 , n45666 , n45667 );
xor ( n45669 , n45665 , n45668 );
nor ( n45670 , n14138 , n798 );
xor ( n45671 , n45669 , n45670 );
and ( n45672 , n44459 , n44460 );
and ( n45673 , n44461 , n44464 );
or ( n45674 , n45672 , n45673 );
xor ( n45675 , n45671 , n45674 );
nor ( n45676 , n14959 , n870 );
xor ( n45677 , n45675 , n45676 );
and ( n45678 , n44465 , n44466 );
and ( n45679 , n44467 , n44470 );
or ( n45680 , n45678 , n45679 );
xor ( n45681 , n45677 , n45680 );
nor ( n45682 , n15800 , n960 );
xor ( n45683 , n45681 , n45682 );
and ( n45684 , n44471 , n44472 );
and ( n45685 , n44473 , n44476 );
or ( n45686 , n45684 , n45685 );
xor ( n45687 , n45683 , n45686 );
nor ( n45688 , n16660 , n1064 );
xor ( n45689 , n45687 , n45688 );
and ( n45690 , n44477 , n44478 );
and ( n45691 , n44479 , n44482 );
or ( n45692 , n45690 , n45691 );
xor ( n45693 , n45689 , n45692 );
nor ( n45694 , n17539 , n1178 );
xor ( n45695 , n45693 , n45694 );
and ( n45696 , n44483 , n44484 );
and ( n45697 , n44485 , n44488 );
or ( n45698 , n45696 , n45697 );
xor ( n45699 , n45695 , n45698 );
nor ( n45700 , n18439 , n1305 );
xor ( n45701 , n45699 , n45700 );
and ( n45702 , n44489 , n44490 );
and ( n45703 , n44491 , n44494 );
or ( n45704 , n45702 , n45703 );
xor ( n45705 , n45701 , n45704 );
nor ( n45706 , n19356 , n1447 );
xor ( n45707 , n45705 , n45706 );
and ( n45708 , n44495 , n44496 );
and ( n45709 , n44497 , n44500 );
or ( n45710 , n45708 , n45709 );
xor ( n45711 , n45707 , n45710 );
nor ( n45712 , n20294 , n1600 );
xor ( n45713 , n45711 , n45712 );
and ( n45714 , n44501 , n44502 );
and ( n45715 , n44503 , n44506 );
or ( n45716 , n45714 , n45715 );
xor ( n45717 , n45713 , n45716 );
nor ( n45718 , n21249 , n1768 );
xor ( n45719 , n45717 , n45718 );
and ( n45720 , n44507 , n44508 );
and ( n45721 , n44509 , n44512 );
or ( n45722 , n45720 , n45721 );
xor ( n45723 , n45719 , n45722 );
nor ( n45724 , n22222 , n1947 );
xor ( n45725 , n45723 , n45724 );
and ( n45726 , n44513 , n44514 );
and ( n45727 , n44515 , n44518 );
or ( n45728 , n45726 , n45727 );
xor ( n45729 , n45725 , n45728 );
nor ( n45730 , n23216 , n2139 );
xor ( n45731 , n45729 , n45730 );
and ( n45732 , n44519 , n44520 );
and ( n45733 , n44521 , n44524 );
or ( n45734 , n45732 , n45733 );
xor ( n45735 , n45731 , n45734 );
nor ( n45736 , n24233 , n2345 );
xor ( n45737 , n45735 , n45736 );
and ( n45738 , n44525 , n44526 );
and ( n45739 , n44527 , n44530 );
or ( n45740 , n45738 , n45739 );
xor ( n45741 , n45737 , n45740 );
nor ( n45742 , n25263 , n2568 );
xor ( n45743 , n45741 , n45742 );
and ( n45744 , n44531 , n44532 );
and ( n45745 , n44533 , n44536 );
or ( n45746 , n45744 , n45745 );
xor ( n45747 , n45743 , n45746 );
nor ( n45748 , n26317 , n2799 );
xor ( n45749 , n45747 , n45748 );
and ( n45750 , n44537 , n44538 );
and ( n45751 , n44539 , n44542 );
or ( n45752 , n45750 , n45751 );
xor ( n45753 , n45749 , n45752 );
nor ( n45754 , n27388 , n3045 );
xor ( n45755 , n45753 , n45754 );
and ( n45756 , n44543 , n44544 );
and ( n45757 , n44545 , n44548 );
or ( n45758 , n45756 , n45757 );
xor ( n45759 , n45755 , n45758 );
nor ( n45760 , n28478 , n3302 );
xor ( n45761 , n45759 , n45760 );
and ( n45762 , n44549 , n44550 );
and ( n45763 , n44551 , n44554 );
or ( n45764 , n45762 , n45763 );
xor ( n45765 , n45761 , n45764 );
nor ( n45766 , n29587 , n3572 );
xor ( n45767 , n45765 , n45766 );
and ( n45768 , n44555 , n44556 );
and ( n45769 , n44557 , n44560 );
or ( n45770 , n45768 , n45769 );
xor ( n45771 , n45767 , n45770 );
nor ( n45772 , n30716 , n3855 );
xor ( n45773 , n45771 , n45772 );
and ( n45774 , n44561 , n44562 );
and ( n45775 , n44563 , n44566 );
or ( n45776 , n45774 , n45775 );
xor ( n45777 , n45773 , n45776 );
nor ( n45778 , n31858 , n4153 );
xor ( n45779 , n45777 , n45778 );
and ( n45780 , n44567 , n44568 );
and ( n45781 , n44569 , n44572 );
or ( n45782 , n45780 , n45781 );
xor ( n45783 , n45779 , n45782 );
nor ( n45784 , n33024 , n4460 );
xor ( n45785 , n45783 , n45784 );
and ( n45786 , n44573 , n44574 );
and ( n45787 , n44575 , n44578 );
or ( n45788 , n45786 , n45787 );
xor ( n45789 , n45785 , n45788 );
nor ( n45790 , n34215 , n4788 );
xor ( n45791 , n45789 , n45790 );
and ( n45792 , n44579 , n44580 );
and ( n45793 , n44581 , n44584 );
or ( n45794 , n45792 , n45793 );
xor ( n45795 , n45791 , n45794 );
nor ( n45796 , n35410 , n5128 );
xor ( n45797 , n45795 , n45796 );
and ( n45798 , n44585 , n44586 );
and ( n45799 , n44587 , n44590 );
or ( n45800 , n45798 , n45799 );
xor ( n45801 , n45797 , n45800 );
nor ( n45802 , n36611 , n5479 );
xor ( n45803 , n45801 , n45802 );
and ( n45804 , n44591 , n44592 );
and ( n45805 , n44593 , n44596 );
or ( n45806 , n45804 , n45805 );
xor ( n45807 , n45803 , n45806 );
nor ( n45808 , n37816 , n5840 );
xor ( n45809 , n45807 , n45808 );
and ( n45810 , n44597 , n44598 );
and ( n45811 , n44599 , n44602 );
or ( n45812 , n45810 , n45811 );
xor ( n45813 , n45809 , n45812 );
nor ( n45814 , n39018 , n6214 );
xor ( n45815 , n45813 , n45814 );
and ( n45816 , n44603 , n44604 );
and ( n45817 , n44605 , n44608 );
or ( n45818 , n45816 , n45817 );
xor ( n45819 , n45815 , n45818 );
nor ( n45820 , n40223 , n6598 );
xor ( n45821 , n45819 , n45820 );
and ( n45822 , n44609 , n44610 );
and ( n45823 , n44611 , n44614 );
or ( n45824 , n45822 , n45823 );
xor ( n45825 , n45821 , n45824 );
nor ( n45826 , n41428 , n6999 );
xor ( n45827 , n45825 , n45826 );
and ( n45828 , n44615 , n44616 );
and ( n45829 , n44617 , n44620 );
or ( n45830 , n45828 , n45829 );
xor ( n45831 , n45827 , n45830 );
nor ( n45832 , n42632 , n7415 );
xor ( n45833 , n45831 , n45832 );
and ( n45834 , n44621 , n44622 );
and ( n45835 , n44623 , n44626 );
or ( n45836 , n45834 , n45835 );
xor ( n45837 , n45833 , n45836 );
nor ( n45838 , n43834 , n7843 );
xor ( n45839 , n45837 , n45838 );
and ( n45840 , n44627 , n44628 );
and ( n45841 , n44629 , n44632 );
or ( n45842 , n45840 , n45841 );
xor ( n45843 , n45839 , n45842 );
nor ( n45844 , n45038 , n8283 );
xor ( n45845 , n45843 , n45844 );
and ( n45846 , n44633 , n44634 );
and ( n45847 , n44635 , n44638 );
or ( n45848 , n45846 , n45847 );
xor ( n45849 , n45845 , n45848 );
and ( n45850 , n44651 , n44655 );
and ( n45851 , n44655 , n45024 );
and ( n45852 , n44651 , n45024 );
or ( n45853 , n45850 , n45851 , n45852 );
and ( n45854 , n33774 , n1134 );
not ( n45855 , n1134 );
nor ( n45856 , n45854 , n45855 );
xor ( n45857 , n45853 , n45856 );
and ( n45858 , n44664 , n44668 );
and ( n45859 , n44668 , n44736 );
and ( n45860 , n44664 , n44736 );
or ( n45861 , n45858 , n45859 , n45860 );
and ( n45862 , n44660 , n44737 );
and ( n45863 , n44737 , n45023 );
and ( n45864 , n44660 , n45023 );
or ( n45865 , n45862 , n45863 , n45864 );
xor ( n45866 , n45861 , n45865 );
and ( n45867 , n44742 , n44862 );
and ( n45868 , n44862 , n45022 );
and ( n45869 , n44742 , n45022 );
or ( n45870 , n45867 , n45868 , n45869 );
and ( n45871 , n44673 , n44677 );
and ( n45872 , n44677 , n44735 );
and ( n45873 , n44673 , n44735 );
or ( n45874 , n45871 , n45872 , n45873 );
and ( n45875 , n44746 , n44750 );
and ( n45876 , n44750 , n44861 );
and ( n45877 , n44746 , n44861 );
or ( n45878 , n45875 , n45876 , n45877 );
xor ( n45879 , n45874 , n45878 );
and ( n45880 , n44704 , n44708 );
and ( n45881 , n44708 , n44714 );
and ( n45882 , n44704 , n44714 );
or ( n45883 , n45880 , n45881 , n45882 );
and ( n45884 , n44682 , n44686 );
and ( n45885 , n44686 , n44734 );
and ( n45886 , n44682 , n44734 );
or ( n45887 , n45884 , n45885 , n45886 );
xor ( n45888 , n45883 , n45887 );
and ( n45889 , n44691 , n44695 );
and ( n45890 , n44695 , n44733 );
and ( n45891 , n44691 , n44733 );
or ( n45892 , n45889 , n45890 , n45891 );
and ( n45893 , n44759 , n44784 );
and ( n45894 , n44784 , n44822 );
and ( n45895 , n44759 , n44822 );
or ( n45896 , n45893 , n45894 , n45895 );
xor ( n45897 , n45892 , n45896 );
and ( n45898 , n44700 , n44715 );
and ( n45899 , n44715 , n44732 );
and ( n45900 , n44700 , n44732 );
or ( n45901 , n45898 , n45899 , n45900 );
and ( n45902 , n44763 , n44767 );
and ( n45903 , n44767 , n44783 );
and ( n45904 , n44763 , n44783 );
or ( n45905 , n45902 , n45903 , n45904 );
xor ( n45906 , n45901 , n45905 );
and ( n45907 , n44720 , n44725 );
and ( n45908 , n44725 , n44731 );
and ( n45909 , n44720 , n44731 );
or ( n45910 , n45907 , n45908 , n45909 );
and ( n45911 , n44710 , n44711 );
and ( n45912 , n44711 , n44713 );
and ( n45913 , n44710 , n44713 );
or ( n45914 , n45911 , n45912 , n45913 );
and ( n45915 , n44721 , n44722 );
and ( n45916 , n44722 , n44724 );
and ( n45917 , n44721 , n44724 );
or ( n45918 , n45915 , n45916 , n45917 );
xor ( n45919 , n45914 , n45918 );
and ( n45920 , n30695 , n1551 );
and ( n45921 , n31836 , n1424 );
xor ( n45922 , n45920 , n45921 );
and ( n45923 , n32649 , n1254 );
xor ( n45924 , n45922 , n45923 );
xor ( n45925 , n45919 , n45924 );
xor ( n45926 , n45910 , n45925 );
and ( n45927 , n44727 , n44728 );
and ( n45928 , n44728 , n44730 );
and ( n45929 , n44727 , n44730 );
or ( n45930 , n45927 , n45928 , n45929 );
and ( n45931 , n27361 , n2100 );
and ( n45932 , n28456 , n1882 );
xor ( n45933 , n45931 , n45932 );
and ( n45934 , n29559 , n1738 );
xor ( n45935 , n45933 , n45934 );
xor ( n45936 , n45930 , n45935 );
and ( n45937 , n24214 , n2739 );
and ( n45938 , n25243 , n2544 );
xor ( n45939 , n45937 , n45938 );
and ( n45940 , n26296 , n2298 );
xor ( n45941 , n45939 , n45940 );
xor ( n45942 , n45936 , n45941 );
xor ( n45943 , n45926 , n45942 );
xor ( n45944 , n45906 , n45943 );
xor ( n45945 , n45897 , n45944 );
xor ( n45946 , n45888 , n45945 );
xor ( n45947 , n45879 , n45946 );
xor ( n45948 , n45870 , n45947 );
and ( n45949 , n44867 , n44945 );
and ( n45950 , n44945 , n45021 );
and ( n45951 , n44867 , n45021 );
or ( n45952 , n45949 , n45950 , n45951 );
and ( n45953 , n44755 , n44823 );
and ( n45954 , n44823 , n44860 );
and ( n45955 , n44755 , n44860 );
or ( n45956 , n45953 , n45954 , n45955 );
and ( n45957 , n44871 , n44875 );
and ( n45958 , n44875 , n44944 );
and ( n45959 , n44871 , n44944 );
or ( n45960 , n45957 , n45958 , n45959 );
xor ( n45961 , n45956 , n45960 );
and ( n45962 , n44828 , n44832 );
and ( n45963 , n44832 , n44859 );
and ( n45964 , n44828 , n44859 );
or ( n45965 , n45962 , n45963 , n45964 );
and ( n45966 , n44789 , n44805 );
and ( n45967 , n44805 , n44821 );
and ( n45968 , n44789 , n44821 );
or ( n45969 , n45966 , n45967 , n45968 );
and ( n45970 , n44772 , n44776 );
and ( n45971 , n44776 , n44782 );
and ( n45972 , n44772 , n44782 );
or ( n45973 , n45970 , n45971 , n45972 );
and ( n45974 , n44793 , n44798 );
and ( n45975 , n44798 , n44804 );
and ( n45976 , n44793 , n44804 );
or ( n45977 , n45974 , n45975 , n45976 );
xor ( n45978 , n45973 , n45977 );
and ( n45979 , n44778 , n44779 );
and ( n45980 , n44779 , n44781 );
and ( n45981 , n44778 , n44781 );
or ( n45982 , n45979 , n45980 , n45981 );
and ( n45983 , n44794 , n44795 );
and ( n45984 , n44795 , n44797 );
and ( n45985 , n44794 , n44797 );
or ( n45986 , n45983 , n45984 , n45985 );
xor ( n45987 , n45982 , n45986 );
and ( n45988 , n21216 , n3495 );
and ( n45989 , n22186 , n3271 );
xor ( n45990 , n45988 , n45989 );
and ( n45991 , n22892 , n2981 );
xor ( n45992 , n45990 , n45991 );
xor ( n45993 , n45987 , n45992 );
xor ( n45994 , n45978 , n45993 );
xor ( n45995 , n45969 , n45994 );
and ( n45996 , n44810 , n44814 );
and ( n45997 , n44814 , n44820 );
and ( n45998 , n44810 , n44820 );
or ( n45999 , n45996 , n45997 , n45998 );
and ( n46000 , n44800 , n44801 );
and ( n46001 , n44801 , n44803 );
and ( n46002 , n44800 , n44803 );
or ( n46003 , n46000 , n46001 , n46002 );
and ( n46004 , n18144 , n4403 );
and ( n46005 , n19324 , n4102 );
xor ( n46006 , n46004 , n46005 );
and ( n46007 , n20233 , n3749 );
xor ( n46008 , n46006 , n46007 );
xor ( n46009 , n46003 , n46008 );
and ( n46010 , n15758 , n5408 );
and ( n46011 , n16637 , n5103 );
xor ( n46012 , n46010 , n46011 );
and ( n46013 , n17512 , n4730 );
xor ( n46014 , n46012 , n46013 );
xor ( n46015 , n46009 , n46014 );
xor ( n46016 , n45999 , n46015 );
and ( n46017 , n44816 , n44817 );
and ( n46018 , n44817 , n44819 );
and ( n46019 , n44816 , n44819 );
or ( n46020 , n46017 , n46018 , n46019 );
and ( n46021 , n44847 , n44848 );
and ( n46022 , n44848 , n44850 );
and ( n46023 , n44847 , n44850 );
or ( n46024 , n46021 , n46022 , n46023 );
xor ( n46025 , n46020 , n46024 );
and ( n46026 , n13322 , n6504 );
and ( n46027 , n14118 , n6132 );
xor ( n46028 , n46026 , n46027 );
and ( n46029 , n14938 , n5765 );
xor ( n46030 , n46028 , n46029 );
xor ( n46031 , n46025 , n46030 );
xor ( n46032 , n46016 , n46031 );
xor ( n46033 , n45995 , n46032 );
xor ( n46034 , n45965 , n46033 );
and ( n46035 , n44837 , n44841 );
and ( n46036 , n44841 , n44858 );
and ( n46037 , n44837 , n44858 );
or ( n46038 , n46035 , n46036 , n46037 );
and ( n46039 , n44884 , n44899 );
and ( n46040 , n44899 , n44916 );
and ( n46041 , n44884 , n44916 );
or ( n46042 , n46039 , n46040 , n46041 );
xor ( n46043 , n46038 , n46042 );
and ( n46044 , n44846 , n44851 );
and ( n46045 , n44851 , n44857 );
and ( n46046 , n44846 , n44857 );
or ( n46047 , n46044 , n46045 , n46046 );
and ( n46048 , n44888 , n44892 );
and ( n46049 , n44892 , n44898 );
and ( n46050 , n44888 , n44898 );
or ( n46051 , n46048 , n46049 , n46050 );
xor ( n46052 , n46047 , n46051 );
and ( n46053 , n44853 , n44854 );
and ( n46054 , n44854 , n44856 );
and ( n46055 , n44853 , n44856 );
or ( n46056 , n46053 , n46054 , n46055 );
and ( n46057 , n11015 , n7662 );
and ( n46058 , n11769 , n7310 );
xor ( n46059 , n46057 , n46058 );
and ( n46060 , n12320 , n6971 );
xor ( n46061 , n46059 , n46060 );
xor ( n46062 , n46056 , n46061 );
and ( n46063 , n10291 , n8243 );
buf ( n46064 , n46063 );
xor ( n46065 , n46062 , n46064 );
xor ( n46066 , n46052 , n46065 );
xor ( n46067 , n46043 , n46066 );
xor ( n46068 , n46034 , n46067 );
xor ( n46069 , n45961 , n46068 );
xor ( n46070 , n45952 , n46069 );
and ( n46071 , n44947 , n44972 );
and ( n46072 , n44972 , n45020 );
and ( n46073 , n44947 , n45020 );
or ( n46074 , n46071 , n46072 , n46073 );
and ( n46075 , n44880 , n44917 );
and ( n46076 , n44917 , n44943 );
and ( n46077 , n44880 , n44943 );
or ( n46078 , n46075 , n46076 , n46077 );
and ( n46079 , n44977 , n44981 );
and ( n46080 , n44981 , n45019 );
and ( n46081 , n44977 , n45019 );
or ( n46082 , n46079 , n46080 , n46081 );
xor ( n46083 , n46078 , n46082 );
and ( n46084 , n44922 , n44926 );
and ( n46085 , n44926 , n44942 );
and ( n46086 , n44922 , n44942 );
or ( n46087 , n46084 , n46085 , n46086 );
and ( n46088 , n44904 , n44909 );
and ( n46089 , n44909 , n44915 );
and ( n46090 , n44904 , n44915 );
or ( n46091 , n46088 , n46089 , n46090 );
and ( n46092 , n44894 , n44895 );
and ( n46093 , n44895 , n44897 );
and ( n46094 , n44894 , n44897 );
or ( n46095 , n46092 , n46093 , n46094 );
and ( n46096 , n44905 , n44906 );
and ( n46097 , n44906 , n44908 );
and ( n46098 , n44905 , n44908 );
or ( n46099 , n46096 , n46097 , n46098 );
xor ( n46100 , n46095 , n46099 );
and ( n46101 , n7385 , n11718 );
and ( n46102 , n7808 , n10977 );
xor ( n46103 , n46101 , n46102 );
and ( n46104 , n8079 , n10239 );
xor ( n46105 , n46103 , n46104 );
xor ( n46106 , n46100 , n46105 );
xor ( n46107 , n46091 , n46106 );
and ( n46108 , n44911 , n44912 );
and ( n46109 , n44912 , n44914 );
and ( n46110 , n44911 , n44914 );
or ( n46111 , n46108 , n46109 , n46110 );
and ( n46112 , n6187 , n14044 );
and ( n46113 , n6569 , n13256 );
xor ( n46114 , n46112 , n46113 );
and ( n46115 , n6816 , n12531 );
xor ( n46116 , n46114 , n46115 );
xor ( n46117 , n46111 , n46116 );
and ( n46118 , n4959 , n16550 );
and ( n46119 , n5459 , n15691 );
xor ( n46120 , n46118 , n46119 );
and ( n46121 , n5819 , n14838 );
xor ( n46122 , n46120 , n46121 );
xor ( n46123 , n46117 , n46122 );
xor ( n46124 , n46107 , n46123 );
xor ( n46125 , n46087 , n46124 );
and ( n46126 , n44931 , n44935 );
and ( n46127 , n44935 , n44941 );
and ( n46128 , n44931 , n44941 );
or ( n46129 , n46126 , n46127 , n46128 );
and ( n46130 , n44990 , n44995 );
and ( n46131 , n44995 , n45001 );
and ( n46132 , n44990 , n45001 );
or ( n46133 , n46130 , n46131 , n46132 );
xor ( n46134 , n46129 , n46133 );
and ( n46135 , n44937 , n44938 );
and ( n46136 , n44938 , n44940 );
and ( n46137 , n44937 , n44940 );
or ( n46138 , n46135 , n46136 , n46137 );
and ( n46139 , n44991 , n44992 );
and ( n46140 , n44992 , n44994 );
and ( n46141 , n44991 , n44994 );
or ( n46142 , n46139 , n46140 , n46141 );
xor ( n46143 , n46138 , n46142 );
and ( n46144 , n4132 , n19222 );
and ( n46145 , n4438 , n18407 );
xor ( n46146 , n46144 , n46145 );
and ( n46147 , n4766 , n17422 );
xor ( n46148 , n46146 , n46147 );
xor ( n46149 , n46143 , n46148 );
xor ( n46150 , n46134 , n46149 );
xor ( n46151 , n46125 , n46150 );
xor ( n46152 , n46083 , n46151 );
xor ( n46153 , n46074 , n46152 );
and ( n46154 , n44951 , n44952 );
and ( n46155 , n44952 , n44971 );
and ( n46156 , n44951 , n44971 );
or ( n46157 , n46154 , n46155 , n46156 );
and ( n46158 , n44986 , n45002 );
and ( n46159 , n45002 , n45018 );
and ( n46160 , n44986 , n45018 );
or ( n46161 , n46158 , n46159 , n46160 );
xor ( n46162 , n46157 , n46161 );
and ( n46163 , n45007 , n45011 );
and ( n46164 , n45011 , n45017 );
and ( n46165 , n45007 , n45017 );
or ( n46166 , n46163 , n46164 , n46165 );
and ( n46167 , n44997 , n44998 );
and ( n46168 , n44998 , n45000 );
and ( n46169 , n44997 , n45000 );
or ( n46170 , n46167 , n46168 , n46169 );
and ( n46171 , n3182 , n22065 );
and ( n46172 , n3545 , n20976 );
xor ( n46173 , n46171 , n46172 );
and ( n46174 , n3801 , n20156 );
xor ( n46175 , n46173 , n46174 );
xor ( n46176 , n46170 , n46175 );
and ( n46177 , n2462 , n25163 );
and ( n46178 , n2779 , n24137 );
xor ( n46179 , n46177 , n46178 );
and ( n46180 , n3024 , n23075 );
xor ( n46181 , n46179 , n46180 );
xor ( n46182 , n46176 , n46181 );
xor ( n46183 , n46166 , n46182 );
and ( n46184 , n45013 , n45014 );
and ( n46185 , n45014 , n45016 );
and ( n46186 , n45013 , n45016 );
or ( n46187 , n46184 , n46185 , n46186 );
and ( n46188 , n44958 , n44959 );
and ( n46189 , n44959 , n44961 );
and ( n46190 , n44958 , n44961 );
or ( n46191 , n46188 , n46189 , n46190 );
xor ( n46192 , n46187 , n46191 );
and ( n46193 , n1933 , n28406 );
and ( n46194 , n2120 , n27296 );
xor ( n46195 , n46193 , n46194 );
and ( n46196 , n2324 , n26216 );
xor ( n46197 , n46195 , n46196 );
xor ( n46198 , n46192 , n46197 );
xor ( n46199 , n46183 , n46198 );
xor ( n46200 , n46162 , n46199 );
and ( n46201 , n44957 , n44962 );
and ( n46202 , n44962 , n44970 );
and ( n46203 , n44957 , n44970 );
or ( n46204 , n46201 , n46202 , n46203 );
and ( n46205 , n44966 , n44967 );
and ( n46206 , n44967 , n44969 );
and ( n46207 , n44966 , n44969 );
or ( n46208 , n46205 , n46206 , n46207 );
and ( n46209 , n1383 , n31761 );
and ( n46210 , n1580 , n30629 );
xor ( n46211 , n46209 , n46210 );
and ( n46212 , n1694 , n29508 );
xor ( n46213 , n46211 , n46212 );
xor ( n46214 , n46208 , n46213 );
not ( n46215 , n1164 );
and ( n46216 , n34193 , n1164 );
nor ( n46217 , n46215 , n46216 );
and ( n46218 , n1287 , n32999 );
xor ( n46219 , n46217 , n46218 );
xor ( n46220 , n46214 , n46219 );
xor ( n46221 , n46204 , n46220 );
xor ( n46222 , n46200 , n46221 );
xor ( n46223 , n46153 , n46222 );
xor ( n46224 , n46070 , n46223 );
xor ( n46225 , n45948 , n46224 );
xor ( n46226 , n45866 , n46225 );
xor ( n46227 , n45857 , n46226 );
and ( n46228 , n44643 , n44646 );
and ( n46229 , n44646 , n45025 );
and ( n46230 , n44643 , n45025 );
or ( n46231 , n46228 , n46229 , n46230 );
xor ( n46232 , n46227 , n46231 );
and ( n46233 , n45026 , n45030 );
and ( n46234 , n45031 , n45034 );
or ( n46235 , n46233 , n46234 );
xor ( n46236 , n46232 , n46235 );
buf ( n46237 , n46236 );
buf ( n46238 , n46237 );
not ( n46239 , n46238 );
nor ( n46240 , n46239 , n8739 );
xor ( n46241 , n45849 , n46240 );
and ( n46242 , n44639 , n45039 );
and ( n46243 , n45040 , n45043 );
or ( n46244 , n46242 , n46243 );
xor ( n46245 , n46241 , n46244 );
buf ( n46246 , n46245 );
buf ( n46247 , n46246 );
not ( n46248 , n46247 );
buf ( n46249 , n572 );
not ( n46250 , n46249 );
nor ( n46251 , n46248 , n46250 );
xor ( n46252 , n45475 , n46251 );
xor ( n46253 , n45055 , n45472 );
nor ( n46254 , n45047 , n46250 );
and ( n46255 , n46253 , n46254 );
xor ( n46256 , n46253 , n46254 );
xor ( n46257 , n45059 , n45470 );
nor ( n46258 , n43843 , n46250 );
and ( n46259 , n46257 , n46258 );
xor ( n46260 , n46257 , n46258 );
xor ( n46261 , n45063 , n45468 );
nor ( n46262 , n42641 , n46250 );
and ( n46263 , n46261 , n46262 );
xor ( n46264 , n46261 , n46262 );
xor ( n46265 , n45067 , n45466 );
nor ( n46266 , n41437 , n46250 );
and ( n46267 , n46265 , n46266 );
xor ( n46268 , n46265 , n46266 );
xor ( n46269 , n45071 , n45464 );
nor ( n46270 , n40232 , n46250 );
and ( n46271 , n46269 , n46270 );
xor ( n46272 , n46269 , n46270 );
xor ( n46273 , n45075 , n45462 );
nor ( n46274 , n39027 , n46250 );
and ( n46275 , n46273 , n46274 );
xor ( n46276 , n46273 , n46274 );
xor ( n46277 , n45079 , n45460 );
nor ( n46278 , n37825 , n46250 );
and ( n46279 , n46277 , n46278 );
xor ( n46280 , n46277 , n46278 );
xor ( n46281 , n45083 , n45458 );
nor ( n46282 , n36620 , n46250 );
and ( n46283 , n46281 , n46282 );
xor ( n46284 , n46281 , n46282 );
xor ( n46285 , n45087 , n45456 );
nor ( n46286 , n35419 , n46250 );
and ( n46287 , n46285 , n46286 );
xor ( n46288 , n46285 , n46286 );
xor ( n46289 , n45091 , n45454 );
nor ( n46290 , n34224 , n46250 );
and ( n46291 , n46289 , n46290 );
xor ( n46292 , n46289 , n46290 );
xor ( n46293 , n45095 , n45452 );
nor ( n46294 , n33033 , n46250 );
and ( n46295 , n46293 , n46294 );
xor ( n46296 , n46293 , n46294 );
xor ( n46297 , n45099 , n45450 );
nor ( n46298 , n31867 , n46250 );
and ( n46299 , n46297 , n46298 );
xor ( n46300 , n46297 , n46298 );
xor ( n46301 , n45103 , n45448 );
nor ( n46302 , n30725 , n46250 );
and ( n46303 , n46301 , n46302 );
xor ( n46304 , n46301 , n46302 );
xor ( n46305 , n45107 , n45446 );
nor ( n46306 , n29596 , n46250 );
and ( n46307 , n46305 , n46306 );
xor ( n46308 , n46305 , n46306 );
xor ( n46309 , n45111 , n45444 );
nor ( n46310 , n28487 , n46250 );
and ( n46311 , n46309 , n46310 );
xor ( n46312 , n46309 , n46310 );
xor ( n46313 , n45115 , n45442 );
nor ( n46314 , n27397 , n46250 );
and ( n46315 , n46313 , n46314 );
xor ( n46316 , n46313 , n46314 );
xor ( n46317 , n45119 , n45440 );
nor ( n46318 , n26326 , n46250 );
and ( n46319 , n46317 , n46318 );
xor ( n46320 , n46317 , n46318 );
xor ( n46321 , n45123 , n45438 );
nor ( n46322 , n25272 , n46250 );
and ( n46323 , n46321 , n46322 );
xor ( n46324 , n46321 , n46322 );
xor ( n46325 , n45127 , n45436 );
nor ( n46326 , n24242 , n46250 );
and ( n46327 , n46325 , n46326 );
xor ( n46328 , n46325 , n46326 );
xor ( n46329 , n45131 , n45434 );
nor ( n46330 , n23225 , n46250 );
and ( n46331 , n46329 , n46330 );
xor ( n46332 , n46329 , n46330 );
xor ( n46333 , n45135 , n45432 );
nor ( n46334 , n22231 , n46250 );
and ( n46335 , n46333 , n46334 );
xor ( n46336 , n46333 , n46334 );
xor ( n46337 , n45139 , n45430 );
nor ( n46338 , n21258 , n46250 );
and ( n46339 , n46337 , n46338 );
xor ( n46340 , n46337 , n46338 );
xor ( n46341 , n45143 , n45428 );
nor ( n46342 , n20303 , n46250 );
and ( n46343 , n46341 , n46342 );
xor ( n46344 , n46341 , n46342 );
xor ( n46345 , n45147 , n45426 );
nor ( n46346 , n19365 , n46250 );
and ( n46347 , n46345 , n46346 );
xor ( n46348 , n46345 , n46346 );
xor ( n46349 , n45151 , n45424 );
nor ( n46350 , n18448 , n46250 );
and ( n46351 , n46349 , n46350 );
xor ( n46352 , n46349 , n46350 );
xor ( n46353 , n45155 , n45422 );
nor ( n46354 , n17548 , n46250 );
and ( n46355 , n46353 , n46354 );
xor ( n46356 , n46353 , n46354 );
xor ( n46357 , n45159 , n45420 );
nor ( n46358 , n16669 , n46250 );
and ( n46359 , n46357 , n46358 );
xor ( n46360 , n46357 , n46358 );
xor ( n46361 , n45163 , n45418 );
nor ( n46362 , n15809 , n46250 );
and ( n46363 , n46361 , n46362 );
xor ( n46364 , n46361 , n46362 );
xor ( n46365 , n45167 , n45416 );
nor ( n46366 , n14968 , n46250 );
and ( n46367 , n46365 , n46366 );
xor ( n46368 , n46365 , n46366 );
xor ( n46369 , n45171 , n45414 );
nor ( n46370 , n14147 , n46250 );
and ( n46371 , n46369 , n46370 );
xor ( n46372 , n46369 , n46370 );
xor ( n46373 , n45175 , n45412 );
nor ( n46374 , n13349 , n46250 );
and ( n46375 , n46373 , n46374 );
xor ( n46376 , n46373 , n46374 );
xor ( n46377 , n45179 , n45410 );
nor ( n46378 , n12564 , n46250 );
and ( n46379 , n46377 , n46378 );
xor ( n46380 , n46377 , n46378 );
xor ( n46381 , n45183 , n45408 );
nor ( n46382 , n11799 , n46250 );
and ( n46383 , n46381 , n46382 );
xor ( n46384 , n46381 , n46382 );
xor ( n46385 , n45187 , n45406 );
nor ( n46386 , n11050 , n46250 );
and ( n46387 , n46385 , n46386 );
xor ( n46388 , n46385 , n46386 );
xor ( n46389 , n45191 , n45404 );
nor ( n46390 , n10321 , n46250 );
and ( n46391 , n46389 , n46390 );
xor ( n46392 , n46389 , n46390 );
xor ( n46393 , n45195 , n45402 );
nor ( n46394 , n9429 , n46250 );
and ( n46395 , n46393 , n46394 );
xor ( n46396 , n46393 , n46394 );
xor ( n46397 , n45199 , n45400 );
nor ( n46398 , n8949 , n46250 );
and ( n46399 , n46397 , n46398 );
xor ( n46400 , n46397 , n46398 );
xor ( n46401 , n45203 , n45398 );
nor ( n46402 , n9437 , n46250 );
and ( n46403 , n46401 , n46402 );
xor ( n46404 , n46401 , n46402 );
xor ( n46405 , n45207 , n45396 );
nor ( n46406 , n9446 , n46250 );
and ( n46407 , n46405 , n46406 );
xor ( n46408 , n46405 , n46406 );
xor ( n46409 , n45211 , n45394 );
nor ( n46410 , n9455 , n46250 );
and ( n46411 , n46409 , n46410 );
xor ( n46412 , n46409 , n46410 );
xor ( n46413 , n45215 , n45392 );
nor ( n46414 , n9464 , n46250 );
and ( n46415 , n46413 , n46414 );
xor ( n46416 , n46413 , n46414 );
xor ( n46417 , n45219 , n45390 );
nor ( n46418 , n9473 , n46250 );
and ( n46419 , n46417 , n46418 );
xor ( n46420 , n46417 , n46418 );
xor ( n46421 , n45223 , n45388 );
nor ( n46422 , n9482 , n46250 );
and ( n46423 , n46421 , n46422 );
xor ( n46424 , n46421 , n46422 );
xor ( n46425 , n45227 , n45386 );
nor ( n46426 , n9491 , n46250 );
and ( n46427 , n46425 , n46426 );
xor ( n46428 , n46425 , n46426 );
xor ( n46429 , n45231 , n45384 );
nor ( n46430 , n9500 , n46250 );
and ( n46431 , n46429 , n46430 );
xor ( n46432 , n46429 , n46430 );
xor ( n46433 , n45235 , n45382 );
nor ( n46434 , n9509 , n46250 );
and ( n46435 , n46433 , n46434 );
xor ( n46436 , n46433 , n46434 );
xor ( n46437 , n45239 , n45380 );
nor ( n46438 , n9518 , n46250 );
and ( n46439 , n46437 , n46438 );
xor ( n46440 , n46437 , n46438 );
xor ( n46441 , n45243 , n45378 );
nor ( n46442 , n9527 , n46250 );
and ( n46443 , n46441 , n46442 );
xor ( n46444 , n46441 , n46442 );
xor ( n46445 , n45247 , n45376 );
nor ( n46446 , n9536 , n46250 );
and ( n46447 , n46445 , n46446 );
xor ( n46448 , n46445 , n46446 );
xor ( n46449 , n45251 , n45374 );
nor ( n46450 , n9545 , n46250 );
and ( n46451 , n46449 , n46450 );
xor ( n46452 , n46449 , n46450 );
xor ( n46453 , n45255 , n45372 );
nor ( n46454 , n9554 , n46250 );
and ( n46455 , n46453 , n46454 );
xor ( n46456 , n46453 , n46454 );
xor ( n46457 , n45259 , n45370 );
nor ( n46458 , n9563 , n46250 );
and ( n46459 , n46457 , n46458 );
xor ( n46460 , n46457 , n46458 );
xor ( n46461 , n45263 , n45368 );
nor ( n46462 , n9572 , n46250 );
and ( n46463 , n46461 , n46462 );
xor ( n46464 , n46461 , n46462 );
xor ( n46465 , n45267 , n45366 );
nor ( n46466 , n9581 , n46250 );
and ( n46467 , n46465 , n46466 );
xor ( n46468 , n46465 , n46466 );
xor ( n46469 , n45271 , n45364 );
nor ( n46470 , n9590 , n46250 );
and ( n46471 , n46469 , n46470 );
xor ( n46472 , n46469 , n46470 );
xor ( n46473 , n45275 , n45362 );
nor ( n46474 , n9599 , n46250 );
and ( n46475 , n46473 , n46474 );
xor ( n46476 , n46473 , n46474 );
xor ( n46477 , n45279 , n45360 );
nor ( n46478 , n9608 , n46250 );
and ( n46479 , n46477 , n46478 );
xor ( n46480 , n46477 , n46478 );
xor ( n46481 , n45283 , n45358 );
nor ( n46482 , n9617 , n46250 );
and ( n46483 , n46481 , n46482 );
xor ( n46484 , n46481 , n46482 );
xor ( n46485 , n45287 , n45356 );
nor ( n46486 , n9626 , n46250 );
and ( n46487 , n46485 , n46486 );
xor ( n46488 , n46485 , n46486 );
xor ( n46489 , n45291 , n45354 );
nor ( n46490 , n9635 , n46250 );
and ( n46491 , n46489 , n46490 );
xor ( n46492 , n46489 , n46490 );
xor ( n46493 , n45295 , n45352 );
nor ( n46494 , n9644 , n46250 );
and ( n46495 , n46493 , n46494 );
xor ( n46496 , n46493 , n46494 );
xor ( n46497 , n45299 , n45350 );
nor ( n46498 , n9653 , n46250 );
and ( n46499 , n46497 , n46498 );
xor ( n46500 , n46497 , n46498 );
xor ( n46501 , n45303 , n45348 );
nor ( n46502 , n9662 , n46250 );
and ( n46503 , n46501 , n46502 );
xor ( n46504 , n46501 , n46502 );
xor ( n46505 , n45307 , n45346 );
nor ( n46506 , n9671 , n46250 );
and ( n46507 , n46505 , n46506 );
xor ( n46508 , n46505 , n46506 );
xor ( n46509 , n45311 , n45344 );
nor ( n46510 , n9680 , n46250 );
and ( n46511 , n46509 , n46510 );
xor ( n46512 , n46509 , n46510 );
xor ( n46513 , n45315 , n45342 );
nor ( n46514 , n9689 , n46250 );
and ( n46515 , n46513 , n46514 );
xor ( n46516 , n46513 , n46514 );
xor ( n46517 , n45319 , n45340 );
nor ( n46518 , n9698 , n46250 );
and ( n46519 , n46517 , n46518 );
xor ( n46520 , n46517 , n46518 );
xor ( n46521 , n45323 , n45338 );
nor ( n46522 , n9707 , n46250 );
and ( n46523 , n46521 , n46522 );
xor ( n46524 , n46521 , n46522 );
xor ( n46525 , n45327 , n45336 );
nor ( n46526 , n9716 , n46250 );
and ( n46527 , n46525 , n46526 );
xor ( n46528 , n46525 , n46526 );
xor ( n46529 , n45331 , n45334 );
nor ( n46530 , n9725 , n46250 );
and ( n46531 , n46529 , n46530 );
xor ( n46532 , n46529 , n46530 );
xor ( n46533 , n45332 , n45333 );
nor ( n46534 , n9734 , n46250 );
and ( n46535 , n46533 , n46534 );
xor ( n46536 , n46533 , n46534 );
nor ( n46537 , n9752 , n45049 );
nor ( n46538 , n9743 , n46250 );
and ( n46539 , n46537 , n46538 );
and ( n46540 , n46536 , n46539 );
or ( n46541 , n46535 , n46540 );
and ( n46542 , n46532 , n46541 );
or ( n46543 , n46531 , n46542 );
and ( n46544 , n46528 , n46543 );
or ( n46545 , n46527 , n46544 );
and ( n46546 , n46524 , n46545 );
or ( n46547 , n46523 , n46546 );
and ( n46548 , n46520 , n46547 );
or ( n46549 , n46519 , n46548 );
and ( n46550 , n46516 , n46549 );
or ( n46551 , n46515 , n46550 );
and ( n46552 , n46512 , n46551 );
or ( n46553 , n46511 , n46552 );
and ( n46554 , n46508 , n46553 );
or ( n46555 , n46507 , n46554 );
and ( n46556 , n46504 , n46555 );
or ( n46557 , n46503 , n46556 );
and ( n46558 , n46500 , n46557 );
or ( n46559 , n46499 , n46558 );
and ( n46560 , n46496 , n46559 );
or ( n46561 , n46495 , n46560 );
and ( n46562 , n46492 , n46561 );
or ( n46563 , n46491 , n46562 );
and ( n46564 , n46488 , n46563 );
or ( n46565 , n46487 , n46564 );
and ( n46566 , n46484 , n46565 );
or ( n46567 , n46483 , n46566 );
and ( n46568 , n46480 , n46567 );
or ( n46569 , n46479 , n46568 );
and ( n46570 , n46476 , n46569 );
or ( n46571 , n46475 , n46570 );
and ( n46572 , n46472 , n46571 );
or ( n46573 , n46471 , n46572 );
and ( n46574 , n46468 , n46573 );
or ( n46575 , n46467 , n46574 );
and ( n46576 , n46464 , n46575 );
or ( n46577 , n46463 , n46576 );
and ( n46578 , n46460 , n46577 );
or ( n46579 , n46459 , n46578 );
and ( n46580 , n46456 , n46579 );
or ( n46581 , n46455 , n46580 );
and ( n46582 , n46452 , n46581 );
or ( n46583 , n46451 , n46582 );
and ( n46584 , n46448 , n46583 );
or ( n46585 , n46447 , n46584 );
and ( n46586 , n46444 , n46585 );
or ( n46587 , n46443 , n46586 );
and ( n46588 , n46440 , n46587 );
or ( n46589 , n46439 , n46588 );
and ( n46590 , n46436 , n46589 );
or ( n46591 , n46435 , n46590 );
and ( n46592 , n46432 , n46591 );
or ( n46593 , n46431 , n46592 );
and ( n46594 , n46428 , n46593 );
or ( n46595 , n46427 , n46594 );
and ( n46596 , n46424 , n46595 );
or ( n46597 , n46423 , n46596 );
and ( n46598 , n46420 , n46597 );
or ( n46599 , n46419 , n46598 );
and ( n46600 , n46416 , n46599 );
or ( n46601 , n46415 , n46600 );
and ( n46602 , n46412 , n46601 );
or ( n46603 , n46411 , n46602 );
and ( n46604 , n46408 , n46603 );
or ( n46605 , n46407 , n46604 );
and ( n46606 , n46404 , n46605 );
or ( n46607 , n46403 , n46606 );
and ( n46608 , n46400 , n46607 );
or ( n46609 , n46399 , n46608 );
and ( n46610 , n46396 , n46609 );
or ( n46611 , n46395 , n46610 );
and ( n46612 , n46392 , n46611 );
or ( n46613 , n46391 , n46612 );
and ( n46614 , n46388 , n46613 );
or ( n46615 , n46387 , n46614 );
and ( n46616 , n46384 , n46615 );
or ( n46617 , n46383 , n46616 );
and ( n46618 , n46380 , n46617 );
or ( n46619 , n46379 , n46618 );
and ( n46620 , n46376 , n46619 );
or ( n46621 , n46375 , n46620 );
and ( n46622 , n46372 , n46621 );
or ( n46623 , n46371 , n46622 );
and ( n46624 , n46368 , n46623 );
or ( n46625 , n46367 , n46624 );
and ( n46626 , n46364 , n46625 );
or ( n46627 , n46363 , n46626 );
and ( n46628 , n46360 , n46627 );
or ( n46629 , n46359 , n46628 );
and ( n46630 , n46356 , n46629 );
or ( n46631 , n46355 , n46630 );
and ( n46632 , n46352 , n46631 );
or ( n46633 , n46351 , n46632 );
and ( n46634 , n46348 , n46633 );
or ( n46635 , n46347 , n46634 );
and ( n46636 , n46344 , n46635 );
or ( n46637 , n46343 , n46636 );
and ( n46638 , n46340 , n46637 );
or ( n46639 , n46339 , n46638 );
and ( n46640 , n46336 , n46639 );
or ( n46641 , n46335 , n46640 );
and ( n46642 , n46332 , n46641 );
or ( n46643 , n46331 , n46642 );
and ( n46644 , n46328 , n46643 );
or ( n46645 , n46327 , n46644 );
and ( n46646 , n46324 , n46645 );
or ( n46647 , n46323 , n46646 );
and ( n46648 , n46320 , n46647 );
or ( n46649 , n46319 , n46648 );
and ( n46650 , n46316 , n46649 );
or ( n46651 , n46315 , n46650 );
and ( n46652 , n46312 , n46651 );
or ( n46653 , n46311 , n46652 );
and ( n46654 , n46308 , n46653 );
or ( n46655 , n46307 , n46654 );
and ( n46656 , n46304 , n46655 );
or ( n46657 , n46303 , n46656 );
and ( n46658 , n46300 , n46657 );
or ( n46659 , n46299 , n46658 );
and ( n46660 , n46296 , n46659 );
or ( n46661 , n46295 , n46660 );
and ( n46662 , n46292 , n46661 );
or ( n46663 , n46291 , n46662 );
and ( n46664 , n46288 , n46663 );
or ( n46665 , n46287 , n46664 );
and ( n46666 , n46284 , n46665 );
or ( n46667 , n46283 , n46666 );
and ( n46668 , n46280 , n46667 );
or ( n46669 , n46279 , n46668 );
and ( n46670 , n46276 , n46669 );
or ( n46671 , n46275 , n46670 );
and ( n46672 , n46272 , n46671 );
or ( n46673 , n46271 , n46672 );
and ( n46674 , n46268 , n46673 );
or ( n46675 , n46267 , n46674 );
and ( n46676 , n46264 , n46675 );
or ( n46677 , n46263 , n46676 );
and ( n46678 , n46260 , n46677 );
or ( n46679 , n46259 , n46678 );
and ( n46680 , n46256 , n46679 );
or ( n46681 , n46255 , n46680 );
xor ( n46682 , n46252 , n46681 );
and ( n46683 , n33403 , n1302 );
nor ( n46684 , n1303 , n46683 );
nor ( n46685 , n1445 , n32231 );
xor ( n46686 , n46684 , n46685 );
and ( n46687 , n45477 , n45478 );
and ( n46688 , n45479 , n45482 );
or ( n46689 , n46687 , n46688 );
xor ( n46690 , n46686 , n46689 );
nor ( n46691 , n1598 , n31083 );
xor ( n46692 , n46690 , n46691 );
and ( n46693 , n45483 , n45484 );
and ( n46694 , n45485 , n45488 );
or ( n46695 , n46693 , n46694 );
xor ( n46696 , n46692 , n46695 );
nor ( n46697 , n1766 , n29948 );
xor ( n46698 , n46696 , n46697 );
and ( n46699 , n45489 , n45490 );
and ( n46700 , n45491 , n45494 );
or ( n46701 , n46699 , n46700 );
xor ( n46702 , n46698 , n46701 );
nor ( n46703 , n1945 , n28833 );
xor ( n46704 , n46702 , n46703 );
and ( n46705 , n45495 , n45496 );
and ( n46706 , n45497 , n45500 );
or ( n46707 , n46705 , n46706 );
xor ( n46708 , n46704 , n46707 );
nor ( n46709 , n2137 , n27737 );
xor ( n46710 , n46708 , n46709 );
and ( n46711 , n45501 , n45502 );
and ( n46712 , n45503 , n45506 );
or ( n46713 , n46711 , n46712 );
xor ( n46714 , n46710 , n46713 );
nor ( n46715 , n2343 , n26660 );
xor ( n46716 , n46714 , n46715 );
and ( n46717 , n45507 , n45508 );
and ( n46718 , n45509 , n45512 );
or ( n46719 , n46717 , n46718 );
xor ( n46720 , n46716 , n46719 );
nor ( n46721 , n2566 , n25600 );
xor ( n46722 , n46720 , n46721 );
and ( n46723 , n45513 , n45514 );
and ( n46724 , n45515 , n45518 );
or ( n46725 , n46723 , n46724 );
xor ( n46726 , n46722 , n46725 );
nor ( n46727 , n2797 , n24564 );
xor ( n46728 , n46726 , n46727 );
and ( n46729 , n45519 , n45520 );
and ( n46730 , n45521 , n45524 );
or ( n46731 , n46729 , n46730 );
xor ( n46732 , n46728 , n46731 );
nor ( n46733 , n3043 , n23541 );
xor ( n46734 , n46732 , n46733 );
and ( n46735 , n45525 , n45526 );
and ( n46736 , n45527 , n45530 );
or ( n46737 , n46735 , n46736 );
xor ( n46738 , n46734 , n46737 );
nor ( n46739 , n3300 , n22541 );
xor ( n46740 , n46738 , n46739 );
and ( n46741 , n45531 , n45532 );
and ( n46742 , n45533 , n45536 );
or ( n46743 , n46741 , n46742 );
xor ( n46744 , n46740 , n46743 );
nor ( n46745 , n3570 , n21562 );
xor ( n46746 , n46744 , n46745 );
and ( n46747 , n45537 , n45538 );
and ( n46748 , n45539 , n45542 );
or ( n46749 , n46747 , n46748 );
xor ( n46750 , n46746 , n46749 );
nor ( n46751 , n3853 , n20601 );
xor ( n46752 , n46750 , n46751 );
and ( n46753 , n45543 , n45544 );
and ( n46754 , n45545 , n45548 );
or ( n46755 , n46753 , n46754 );
xor ( n46756 , n46752 , n46755 );
nor ( n46757 , n4151 , n19657 );
xor ( n46758 , n46756 , n46757 );
and ( n46759 , n45549 , n45550 );
and ( n46760 , n45551 , n45554 );
or ( n46761 , n46759 , n46760 );
xor ( n46762 , n46758 , n46761 );
nor ( n46763 , n4458 , n18734 );
xor ( n46764 , n46762 , n46763 );
and ( n46765 , n45555 , n45556 );
and ( n46766 , n45557 , n45560 );
or ( n46767 , n46765 , n46766 );
xor ( n46768 , n46764 , n46767 );
nor ( n46769 , n4786 , n17828 );
xor ( n46770 , n46768 , n46769 );
and ( n46771 , n45561 , n45562 );
and ( n46772 , n45563 , n45566 );
or ( n46773 , n46771 , n46772 );
xor ( n46774 , n46770 , n46773 );
nor ( n46775 , n5126 , n16943 );
xor ( n46776 , n46774 , n46775 );
and ( n46777 , n45567 , n45568 );
and ( n46778 , n45569 , n45572 );
or ( n46779 , n46777 , n46778 );
xor ( n46780 , n46776 , n46779 );
nor ( n46781 , n5477 , n16077 );
xor ( n46782 , n46780 , n46781 );
and ( n46783 , n45573 , n45574 );
and ( n46784 , n45575 , n45578 );
or ( n46785 , n46783 , n46784 );
xor ( n46786 , n46782 , n46785 );
nor ( n46787 , n5838 , n15230 );
xor ( n46788 , n46786 , n46787 );
and ( n46789 , n45579 , n45580 );
and ( n46790 , n45581 , n45584 );
or ( n46791 , n46789 , n46790 );
xor ( n46792 , n46788 , n46791 );
nor ( n46793 , n6212 , n14403 );
xor ( n46794 , n46792 , n46793 );
and ( n46795 , n45585 , n45586 );
and ( n46796 , n45587 , n45590 );
or ( n46797 , n46795 , n46796 );
xor ( n46798 , n46794 , n46797 );
nor ( n46799 , n6596 , n13599 );
xor ( n46800 , n46798 , n46799 );
and ( n46801 , n45591 , n45592 );
and ( n46802 , n45593 , n45596 );
or ( n46803 , n46801 , n46802 );
xor ( n46804 , n46800 , n46803 );
nor ( n46805 , n6997 , n12808 );
xor ( n46806 , n46804 , n46805 );
and ( n46807 , n45597 , n45598 );
and ( n46808 , n45599 , n45602 );
or ( n46809 , n46807 , n46808 );
xor ( n46810 , n46806 , n46809 );
nor ( n46811 , n7413 , n12037 );
xor ( n46812 , n46810 , n46811 );
and ( n46813 , n45603 , n45604 );
and ( n46814 , n45605 , n45608 );
or ( n46815 , n46813 , n46814 );
xor ( n46816 , n46812 , n46815 );
nor ( n46817 , n7841 , n11282 );
xor ( n46818 , n46816 , n46817 );
and ( n46819 , n45609 , n45610 );
and ( n46820 , n45611 , n45614 );
or ( n46821 , n46819 , n46820 );
xor ( n46822 , n46818 , n46821 );
nor ( n46823 , n8281 , n10547 );
xor ( n46824 , n46822 , n46823 );
and ( n46825 , n45615 , n45616 );
and ( n46826 , n45617 , n45620 );
or ( n46827 , n46825 , n46826 );
xor ( n46828 , n46824 , n46827 );
nor ( n46829 , n8737 , n9829 );
xor ( n46830 , n46828 , n46829 );
and ( n46831 , n45621 , n45622 );
and ( n46832 , n45623 , n45626 );
or ( n46833 , n46831 , n46832 );
xor ( n46834 , n46830 , n46833 );
nor ( n46835 , n9420 , n8955 );
xor ( n46836 , n46834 , n46835 );
and ( n46837 , n45627 , n45628 );
and ( n46838 , n45629 , n45632 );
or ( n46839 , n46837 , n46838 );
xor ( n46840 , n46836 , n46839 );
nor ( n46841 , n10312 , n603 );
xor ( n46842 , n46840 , n46841 );
and ( n46843 , n45633 , n45634 );
and ( n46844 , n45635 , n45638 );
or ( n46845 , n46843 , n46844 );
xor ( n46846 , n46842 , n46845 );
nor ( n46847 , n11041 , n652 );
xor ( n46848 , n46846 , n46847 );
and ( n46849 , n45639 , n45640 );
and ( n46850 , n45641 , n45644 );
or ( n46851 , n46849 , n46850 );
xor ( n46852 , n46848 , n46851 );
nor ( n46853 , n11790 , n624 );
xor ( n46854 , n46852 , n46853 );
and ( n46855 , n45645 , n45646 );
and ( n46856 , n45647 , n45650 );
or ( n46857 , n46855 , n46856 );
xor ( n46858 , n46854 , n46857 );
nor ( n46859 , n12555 , n648 );
xor ( n46860 , n46858 , n46859 );
and ( n46861 , n45651 , n45652 );
and ( n46862 , n45653 , n45656 );
or ( n46863 , n46861 , n46862 );
xor ( n46864 , n46860 , n46863 );
nor ( n46865 , n13340 , n686 );
xor ( n46866 , n46864 , n46865 );
and ( n46867 , n45657 , n45658 );
and ( n46868 , n45659 , n45662 );
or ( n46869 , n46867 , n46868 );
xor ( n46870 , n46866 , n46869 );
nor ( n46871 , n14138 , n735 );
xor ( n46872 , n46870 , n46871 );
and ( n46873 , n45663 , n45664 );
and ( n46874 , n45665 , n45668 );
or ( n46875 , n46873 , n46874 );
xor ( n46876 , n46872 , n46875 );
nor ( n46877 , n14959 , n798 );
xor ( n46878 , n46876 , n46877 );
and ( n46879 , n45669 , n45670 );
and ( n46880 , n45671 , n45674 );
or ( n46881 , n46879 , n46880 );
xor ( n46882 , n46878 , n46881 );
nor ( n46883 , n15800 , n870 );
xor ( n46884 , n46882 , n46883 );
and ( n46885 , n45675 , n45676 );
and ( n46886 , n45677 , n45680 );
or ( n46887 , n46885 , n46886 );
xor ( n46888 , n46884 , n46887 );
nor ( n46889 , n16660 , n960 );
xor ( n46890 , n46888 , n46889 );
and ( n46891 , n45681 , n45682 );
and ( n46892 , n45683 , n45686 );
or ( n46893 , n46891 , n46892 );
xor ( n46894 , n46890 , n46893 );
nor ( n46895 , n17539 , n1064 );
xor ( n46896 , n46894 , n46895 );
and ( n46897 , n45687 , n45688 );
and ( n46898 , n45689 , n45692 );
or ( n46899 , n46897 , n46898 );
xor ( n46900 , n46896 , n46899 );
nor ( n46901 , n18439 , n1178 );
xor ( n46902 , n46900 , n46901 );
and ( n46903 , n45693 , n45694 );
and ( n46904 , n45695 , n45698 );
or ( n46905 , n46903 , n46904 );
xor ( n46906 , n46902 , n46905 );
nor ( n46907 , n19356 , n1305 );
xor ( n46908 , n46906 , n46907 );
and ( n46909 , n45699 , n45700 );
and ( n46910 , n45701 , n45704 );
or ( n46911 , n46909 , n46910 );
xor ( n46912 , n46908 , n46911 );
nor ( n46913 , n20294 , n1447 );
xor ( n46914 , n46912 , n46913 );
and ( n46915 , n45705 , n45706 );
and ( n46916 , n45707 , n45710 );
or ( n46917 , n46915 , n46916 );
xor ( n46918 , n46914 , n46917 );
nor ( n46919 , n21249 , n1600 );
xor ( n46920 , n46918 , n46919 );
and ( n46921 , n45711 , n45712 );
and ( n46922 , n45713 , n45716 );
or ( n46923 , n46921 , n46922 );
xor ( n46924 , n46920 , n46923 );
nor ( n46925 , n22222 , n1768 );
xor ( n46926 , n46924 , n46925 );
and ( n46927 , n45717 , n45718 );
and ( n46928 , n45719 , n45722 );
or ( n46929 , n46927 , n46928 );
xor ( n46930 , n46926 , n46929 );
nor ( n46931 , n23216 , n1947 );
xor ( n46932 , n46930 , n46931 );
and ( n46933 , n45723 , n45724 );
and ( n46934 , n45725 , n45728 );
or ( n46935 , n46933 , n46934 );
xor ( n46936 , n46932 , n46935 );
nor ( n46937 , n24233 , n2139 );
xor ( n46938 , n46936 , n46937 );
and ( n46939 , n45729 , n45730 );
and ( n46940 , n45731 , n45734 );
or ( n46941 , n46939 , n46940 );
xor ( n46942 , n46938 , n46941 );
nor ( n46943 , n25263 , n2345 );
xor ( n46944 , n46942 , n46943 );
and ( n46945 , n45735 , n45736 );
and ( n46946 , n45737 , n45740 );
or ( n46947 , n46945 , n46946 );
xor ( n46948 , n46944 , n46947 );
nor ( n46949 , n26317 , n2568 );
xor ( n46950 , n46948 , n46949 );
and ( n46951 , n45741 , n45742 );
and ( n46952 , n45743 , n45746 );
or ( n46953 , n46951 , n46952 );
xor ( n46954 , n46950 , n46953 );
nor ( n46955 , n27388 , n2799 );
xor ( n46956 , n46954 , n46955 );
and ( n46957 , n45747 , n45748 );
and ( n46958 , n45749 , n45752 );
or ( n46959 , n46957 , n46958 );
xor ( n46960 , n46956 , n46959 );
nor ( n46961 , n28478 , n3045 );
xor ( n46962 , n46960 , n46961 );
and ( n46963 , n45753 , n45754 );
and ( n46964 , n45755 , n45758 );
or ( n46965 , n46963 , n46964 );
xor ( n46966 , n46962 , n46965 );
nor ( n46967 , n29587 , n3302 );
xor ( n46968 , n46966 , n46967 );
and ( n46969 , n45759 , n45760 );
and ( n46970 , n45761 , n45764 );
or ( n46971 , n46969 , n46970 );
xor ( n46972 , n46968 , n46971 );
nor ( n46973 , n30716 , n3572 );
xor ( n46974 , n46972 , n46973 );
and ( n46975 , n45765 , n45766 );
and ( n46976 , n45767 , n45770 );
or ( n46977 , n46975 , n46976 );
xor ( n46978 , n46974 , n46977 );
nor ( n46979 , n31858 , n3855 );
xor ( n46980 , n46978 , n46979 );
and ( n46981 , n45771 , n45772 );
and ( n46982 , n45773 , n45776 );
or ( n46983 , n46981 , n46982 );
xor ( n46984 , n46980 , n46983 );
nor ( n46985 , n33024 , n4153 );
xor ( n46986 , n46984 , n46985 );
and ( n46987 , n45777 , n45778 );
and ( n46988 , n45779 , n45782 );
or ( n46989 , n46987 , n46988 );
xor ( n46990 , n46986 , n46989 );
nor ( n46991 , n34215 , n4460 );
xor ( n46992 , n46990 , n46991 );
and ( n46993 , n45783 , n45784 );
and ( n46994 , n45785 , n45788 );
or ( n46995 , n46993 , n46994 );
xor ( n46996 , n46992 , n46995 );
nor ( n46997 , n35410 , n4788 );
xor ( n46998 , n46996 , n46997 );
and ( n46999 , n45789 , n45790 );
and ( n47000 , n45791 , n45794 );
or ( n47001 , n46999 , n47000 );
xor ( n47002 , n46998 , n47001 );
nor ( n47003 , n36611 , n5128 );
xor ( n47004 , n47002 , n47003 );
and ( n47005 , n45795 , n45796 );
and ( n47006 , n45797 , n45800 );
or ( n47007 , n47005 , n47006 );
xor ( n47008 , n47004 , n47007 );
nor ( n47009 , n37816 , n5479 );
xor ( n47010 , n47008 , n47009 );
and ( n47011 , n45801 , n45802 );
and ( n47012 , n45803 , n45806 );
or ( n47013 , n47011 , n47012 );
xor ( n47014 , n47010 , n47013 );
nor ( n47015 , n39018 , n5840 );
xor ( n47016 , n47014 , n47015 );
and ( n47017 , n45807 , n45808 );
and ( n47018 , n45809 , n45812 );
or ( n47019 , n47017 , n47018 );
xor ( n47020 , n47016 , n47019 );
nor ( n47021 , n40223 , n6214 );
xor ( n47022 , n47020 , n47021 );
and ( n47023 , n45813 , n45814 );
and ( n47024 , n45815 , n45818 );
or ( n47025 , n47023 , n47024 );
xor ( n47026 , n47022 , n47025 );
nor ( n47027 , n41428 , n6598 );
xor ( n47028 , n47026 , n47027 );
and ( n47029 , n45819 , n45820 );
and ( n47030 , n45821 , n45824 );
or ( n47031 , n47029 , n47030 );
xor ( n47032 , n47028 , n47031 );
nor ( n47033 , n42632 , n6999 );
xor ( n47034 , n47032 , n47033 );
and ( n47035 , n45825 , n45826 );
and ( n47036 , n45827 , n45830 );
or ( n47037 , n47035 , n47036 );
xor ( n47038 , n47034 , n47037 );
nor ( n47039 , n43834 , n7415 );
xor ( n47040 , n47038 , n47039 );
and ( n47041 , n45831 , n45832 );
and ( n47042 , n45833 , n45836 );
or ( n47043 , n47041 , n47042 );
xor ( n47044 , n47040 , n47043 );
nor ( n47045 , n45038 , n7843 );
xor ( n47046 , n47044 , n47045 );
and ( n47047 , n45837 , n45838 );
and ( n47048 , n45839 , n45842 );
or ( n47049 , n47047 , n47048 );
xor ( n47050 , n47046 , n47049 );
nor ( n47051 , n46239 , n8283 );
xor ( n47052 , n47050 , n47051 );
and ( n47053 , n45843 , n45844 );
and ( n47054 , n45845 , n45848 );
or ( n47055 , n47053 , n47054 );
xor ( n47056 , n47052 , n47055 );
and ( n47057 , n45861 , n45865 );
and ( n47058 , n45865 , n46225 );
and ( n47059 , n45861 , n46225 );
or ( n47060 , n47057 , n47058 , n47059 );
and ( n47061 , n33774 , n1254 );
not ( n47062 , n1254 );
nor ( n47063 , n47061 , n47062 );
xor ( n47064 , n47060 , n47063 );
and ( n47065 , n45874 , n45878 );
and ( n47066 , n45878 , n45946 );
and ( n47067 , n45874 , n45946 );
or ( n47068 , n47065 , n47066 , n47067 );
and ( n47069 , n45870 , n45947 );
and ( n47070 , n45947 , n46224 );
and ( n47071 , n45870 , n46224 );
or ( n47072 , n47069 , n47070 , n47071 );
xor ( n47073 , n47068 , n47072 );
and ( n47074 , n45952 , n46069 );
and ( n47075 , n46069 , n46223 );
and ( n47076 , n45952 , n46223 );
or ( n47077 , n47074 , n47075 , n47076 );
and ( n47078 , n45883 , n45887 );
and ( n47079 , n45887 , n45945 );
and ( n47080 , n45883 , n45945 );
or ( n47081 , n47078 , n47079 , n47080 );
and ( n47082 , n45956 , n45960 );
and ( n47083 , n45960 , n46068 );
and ( n47084 , n45956 , n46068 );
or ( n47085 , n47082 , n47083 , n47084 );
xor ( n47086 , n47081 , n47085 );
and ( n47087 , n45914 , n45918 );
and ( n47088 , n45918 , n45924 );
and ( n47089 , n45914 , n45924 );
or ( n47090 , n47087 , n47088 , n47089 );
and ( n47091 , n45892 , n45896 );
and ( n47092 , n45896 , n45944 );
and ( n47093 , n45892 , n45944 );
or ( n47094 , n47091 , n47092 , n47093 );
xor ( n47095 , n47090 , n47094 );
and ( n47096 , n45901 , n45905 );
and ( n47097 , n45905 , n45943 );
and ( n47098 , n45901 , n45943 );
or ( n47099 , n47096 , n47097 , n47098 );
and ( n47100 , n45969 , n45994 );
and ( n47101 , n45994 , n46032 );
and ( n47102 , n45969 , n46032 );
or ( n47103 , n47100 , n47101 , n47102 );
xor ( n47104 , n47099 , n47103 );
and ( n47105 , n45910 , n45925 );
and ( n47106 , n45925 , n45942 );
and ( n47107 , n45910 , n45942 );
or ( n47108 , n47105 , n47106 , n47107 );
and ( n47109 , n45973 , n45977 );
and ( n47110 , n45977 , n45993 );
and ( n47111 , n45973 , n45993 );
or ( n47112 , n47109 , n47110 , n47111 );
xor ( n47113 , n47108 , n47112 );
and ( n47114 , n45930 , n45935 );
and ( n47115 , n45935 , n45941 );
and ( n47116 , n45930 , n45941 );
or ( n47117 , n47114 , n47115 , n47116 );
and ( n47118 , n45920 , n45921 );
and ( n47119 , n45921 , n45923 );
and ( n47120 , n45920 , n45923 );
or ( n47121 , n47118 , n47119 , n47120 );
and ( n47122 , n45931 , n45932 );
and ( n47123 , n45932 , n45934 );
and ( n47124 , n45931 , n45934 );
or ( n47125 , n47122 , n47123 , n47124 );
xor ( n47126 , n47121 , n47125 );
and ( n47127 , n30695 , n1738 );
and ( n47128 , n31836 , n1551 );
xor ( n47129 , n47127 , n47128 );
and ( n47130 , n32649 , n1424 );
xor ( n47131 , n47129 , n47130 );
xor ( n47132 , n47126 , n47131 );
xor ( n47133 , n47117 , n47132 );
and ( n47134 , n45937 , n45938 );
and ( n47135 , n45938 , n45940 );
and ( n47136 , n45937 , n45940 );
or ( n47137 , n47134 , n47135 , n47136 );
and ( n47138 , n27361 , n2298 );
and ( n47139 , n28456 , n2100 );
xor ( n47140 , n47138 , n47139 );
and ( n47141 , n29559 , n1882 );
xor ( n47142 , n47140 , n47141 );
xor ( n47143 , n47137 , n47142 );
and ( n47144 , n24214 , n2981 );
and ( n47145 , n25243 , n2739 );
xor ( n47146 , n47144 , n47145 );
and ( n47147 , n26296 , n2544 );
xor ( n47148 , n47146 , n47147 );
xor ( n47149 , n47143 , n47148 );
xor ( n47150 , n47133 , n47149 );
xor ( n47151 , n47113 , n47150 );
xor ( n47152 , n47104 , n47151 );
xor ( n47153 , n47095 , n47152 );
xor ( n47154 , n47086 , n47153 );
xor ( n47155 , n47077 , n47154 );
and ( n47156 , n46074 , n46152 );
and ( n47157 , n46152 , n46222 );
and ( n47158 , n46074 , n46222 );
or ( n47159 , n47156 , n47157 , n47158 );
and ( n47160 , n45965 , n46033 );
and ( n47161 , n46033 , n46067 );
and ( n47162 , n45965 , n46067 );
or ( n47163 , n47160 , n47161 , n47162 );
and ( n47164 , n46078 , n46082 );
and ( n47165 , n46082 , n46151 );
and ( n47166 , n46078 , n46151 );
or ( n47167 , n47164 , n47165 , n47166 );
xor ( n47168 , n47163 , n47167 );
and ( n47169 , n46038 , n46042 );
and ( n47170 , n46042 , n46066 );
and ( n47171 , n46038 , n46066 );
or ( n47172 , n47169 , n47170 , n47171 );
and ( n47173 , n45999 , n46015 );
and ( n47174 , n46015 , n46031 );
and ( n47175 , n45999 , n46031 );
or ( n47176 , n47173 , n47174 , n47175 );
and ( n47177 , n45982 , n45986 );
and ( n47178 , n45986 , n45992 );
and ( n47179 , n45982 , n45992 );
or ( n47180 , n47177 , n47178 , n47179 );
and ( n47181 , n46003 , n46008 );
and ( n47182 , n46008 , n46014 );
and ( n47183 , n46003 , n46014 );
or ( n47184 , n47181 , n47182 , n47183 );
xor ( n47185 , n47180 , n47184 );
and ( n47186 , n45988 , n45989 );
and ( n47187 , n45989 , n45991 );
and ( n47188 , n45988 , n45991 );
or ( n47189 , n47186 , n47187 , n47188 );
and ( n47190 , n46004 , n46005 );
and ( n47191 , n46005 , n46007 );
and ( n47192 , n46004 , n46007 );
or ( n47193 , n47190 , n47191 , n47192 );
xor ( n47194 , n47189 , n47193 );
and ( n47195 , n21216 , n3749 );
and ( n47196 , n22186 , n3495 );
xor ( n47197 , n47195 , n47196 );
and ( n47198 , n22892 , n3271 );
xor ( n47199 , n47197 , n47198 );
xor ( n47200 , n47194 , n47199 );
xor ( n47201 , n47185 , n47200 );
xor ( n47202 , n47176 , n47201 );
and ( n47203 , n46020 , n46024 );
and ( n47204 , n46024 , n46030 );
and ( n47205 , n46020 , n46030 );
or ( n47206 , n47203 , n47204 , n47205 );
and ( n47207 , n46010 , n46011 );
and ( n47208 , n46011 , n46013 );
and ( n47209 , n46010 , n46013 );
or ( n47210 , n47207 , n47208 , n47209 );
and ( n47211 , n18144 , n4730 );
and ( n47212 , n19324 , n4403 );
xor ( n47213 , n47211 , n47212 );
and ( n47214 , n20233 , n4102 );
xor ( n47215 , n47213 , n47214 );
xor ( n47216 , n47210 , n47215 );
and ( n47217 , n15758 , n5765 );
and ( n47218 , n16637 , n5408 );
xor ( n47219 , n47217 , n47218 );
and ( n47220 , n17512 , n5103 );
xor ( n47221 , n47219 , n47220 );
xor ( n47222 , n47216 , n47221 );
xor ( n47223 , n47206 , n47222 );
and ( n47224 , n46026 , n46027 );
and ( n47225 , n46027 , n46029 );
and ( n47226 , n46026 , n46029 );
or ( n47227 , n47224 , n47225 , n47226 );
and ( n47228 , n46057 , n46058 );
and ( n47229 , n46058 , n46060 );
and ( n47230 , n46057 , n46060 );
or ( n47231 , n47228 , n47229 , n47230 );
xor ( n47232 , n47227 , n47231 );
and ( n47233 , n13322 , n6971 );
and ( n47234 , n14118 , n6504 );
xor ( n47235 , n47233 , n47234 );
and ( n47236 , n14938 , n6132 );
xor ( n47237 , n47235 , n47236 );
xor ( n47238 , n47232 , n47237 );
xor ( n47239 , n47223 , n47238 );
xor ( n47240 , n47202 , n47239 );
xor ( n47241 , n47172 , n47240 );
and ( n47242 , n46047 , n46051 );
and ( n47243 , n46051 , n46065 );
and ( n47244 , n46047 , n46065 );
or ( n47245 , n47242 , n47243 , n47244 );
and ( n47246 , n46091 , n46106 );
and ( n47247 , n46106 , n46123 );
and ( n47248 , n46091 , n46123 );
or ( n47249 , n47246 , n47247 , n47248 );
xor ( n47250 , n47245 , n47249 );
and ( n47251 , n46056 , n46061 );
and ( n47252 , n46061 , n46064 );
and ( n47253 , n46056 , n46064 );
or ( n47254 , n47251 , n47252 , n47253 );
and ( n47255 , n46095 , n46099 );
and ( n47256 , n46099 , n46105 );
and ( n47257 , n46095 , n46105 );
or ( n47258 , n47255 , n47256 , n47257 );
xor ( n47259 , n47254 , n47258 );
and ( n47260 , n8718 , n9348 );
and ( n47261 , n9400 , n8669 );
and ( n47262 , n47260 , n47261 );
and ( n47263 , n47261 , n46063 );
and ( n47264 , n47260 , n46063 );
or ( n47265 , n47262 , n47263 , n47264 );
and ( n47266 , n11015 , n8243 );
and ( n47267 , n11769 , n7662 );
xor ( n47268 , n47266 , n47267 );
and ( n47269 , n12320 , n7310 );
xor ( n47270 , n47268 , n47269 );
xor ( n47271 , n47265 , n47270 );
and ( n47272 , n8718 , n10239 );
buf ( n47273 , n9400 );
xor ( n47274 , n47272 , n47273 );
and ( n47275 , n10291 , n8669 );
xor ( n47276 , n47274 , n47275 );
xor ( n47277 , n47271 , n47276 );
xor ( n47278 , n47259 , n47277 );
xor ( n47279 , n47250 , n47278 );
xor ( n47280 , n47241 , n47279 );
xor ( n47281 , n47168 , n47280 );
xor ( n47282 , n47159 , n47281 );
and ( n47283 , n46200 , n46221 );
and ( n47284 , n46157 , n46161 );
and ( n47285 , n46161 , n46199 );
and ( n47286 , n46157 , n46199 );
or ( n47287 , n47284 , n47285 , n47286 );
and ( n47288 , n46087 , n46124 );
and ( n47289 , n46124 , n46150 );
and ( n47290 , n46087 , n46150 );
or ( n47291 , n47288 , n47289 , n47290 );
xor ( n47292 , n47287 , n47291 );
and ( n47293 , n46129 , n46133 );
and ( n47294 , n46133 , n46149 );
and ( n47295 , n46129 , n46149 );
or ( n47296 , n47293 , n47294 , n47295 );
and ( n47297 , n46111 , n46116 );
and ( n47298 , n46116 , n46122 );
and ( n47299 , n46111 , n46122 );
or ( n47300 , n47297 , n47298 , n47299 );
and ( n47301 , n46101 , n46102 );
and ( n47302 , n46102 , n46104 );
and ( n47303 , n46101 , n46104 );
or ( n47304 , n47301 , n47302 , n47303 );
and ( n47305 , n46112 , n46113 );
and ( n47306 , n46113 , n46115 );
and ( n47307 , n46112 , n46115 );
or ( n47308 , n47305 , n47306 , n47307 );
xor ( n47309 , n47304 , n47308 );
and ( n47310 , n7385 , n12531 );
and ( n47311 , n7808 , n11718 );
xor ( n47312 , n47310 , n47311 );
and ( n47313 , n8079 , n10977 );
xor ( n47314 , n47312 , n47313 );
xor ( n47315 , n47309 , n47314 );
xor ( n47316 , n47300 , n47315 );
and ( n47317 , n46118 , n46119 );
and ( n47318 , n46119 , n46121 );
and ( n47319 , n46118 , n46121 );
or ( n47320 , n47317 , n47318 , n47319 );
and ( n47321 , n6187 , n14838 );
and ( n47322 , n6569 , n14044 );
xor ( n47323 , n47321 , n47322 );
and ( n47324 , n6816 , n13256 );
xor ( n47325 , n47323 , n47324 );
xor ( n47326 , n47320 , n47325 );
and ( n47327 , n4959 , n17422 );
and ( n47328 , n5459 , n16550 );
xor ( n47329 , n47327 , n47328 );
and ( n47330 , n5819 , n15691 );
xor ( n47331 , n47329 , n47330 );
xor ( n47332 , n47326 , n47331 );
xor ( n47333 , n47316 , n47332 );
xor ( n47334 , n47296 , n47333 );
and ( n47335 , n46138 , n46142 );
and ( n47336 , n46142 , n46148 );
and ( n47337 , n46138 , n46148 );
or ( n47338 , n47335 , n47336 , n47337 );
and ( n47339 , n46170 , n46175 );
and ( n47340 , n46175 , n46181 );
and ( n47341 , n46170 , n46181 );
or ( n47342 , n47339 , n47340 , n47341 );
xor ( n47343 , n47338 , n47342 );
and ( n47344 , n46144 , n46145 );
and ( n47345 , n46145 , n46147 );
and ( n47346 , n46144 , n46147 );
or ( n47347 , n47344 , n47345 , n47346 );
and ( n47348 , n46171 , n46172 );
and ( n47349 , n46172 , n46174 );
and ( n47350 , n46171 , n46174 );
or ( n47351 , n47348 , n47349 , n47350 );
xor ( n47352 , n47347 , n47351 );
and ( n47353 , n4132 , n20156 );
and ( n47354 , n4438 , n19222 );
xor ( n47355 , n47353 , n47354 );
and ( n47356 , n4766 , n18407 );
xor ( n47357 , n47355 , n47356 );
xor ( n47358 , n47352 , n47357 );
xor ( n47359 , n47343 , n47358 );
xor ( n47360 , n47334 , n47359 );
xor ( n47361 , n47292 , n47360 );
xor ( n47362 , n47283 , n47361 );
and ( n47363 , n46166 , n46182 );
and ( n47364 , n46182 , n46198 );
and ( n47365 , n46166 , n46198 );
or ( n47366 , n47363 , n47364 , n47365 );
and ( n47367 , n46204 , n46220 );
xor ( n47368 , n47366 , n47367 );
and ( n47369 , n46187 , n46191 );
and ( n47370 , n46191 , n46197 );
and ( n47371 , n46187 , n46197 );
or ( n47372 , n47369 , n47370 , n47371 );
and ( n47373 , n46177 , n46178 );
and ( n47374 , n46178 , n46180 );
and ( n47375 , n46177 , n46180 );
or ( n47376 , n47373 , n47374 , n47375 );
and ( n47377 , n3182 , n23075 );
and ( n47378 , n3545 , n22065 );
xor ( n47379 , n47377 , n47378 );
and ( n47380 , n3801 , n20976 );
xor ( n47381 , n47379 , n47380 );
xor ( n47382 , n47376 , n47381 );
and ( n47383 , n2462 , n26216 );
and ( n47384 , n2779 , n25163 );
xor ( n47385 , n47383 , n47384 );
and ( n47386 , n3024 , n24137 );
xor ( n47387 , n47385 , n47386 );
xor ( n47388 , n47382 , n47387 );
xor ( n47389 , n47372 , n47388 );
and ( n47390 , n46193 , n46194 );
and ( n47391 , n46194 , n46196 );
and ( n47392 , n46193 , n46196 );
or ( n47393 , n47390 , n47391 , n47392 );
and ( n47394 , n46209 , n46210 );
and ( n47395 , n46210 , n46212 );
and ( n47396 , n46209 , n46212 );
or ( n47397 , n47394 , n47395 , n47396 );
xor ( n47398 , n47393 , n47397 );
and ( n47399 , n1933 , n29508 );
and ( n47400 , n2120 , n28406 );
xor ( n47401 , n47399 , n47400 );
and ( n47402 , n2324 , n27296 );
xor ( n47403 , n47401 , n47402 );
xor ( n47404 , n47398 , n47403 );
xor ( n47405 , n47389 , n47404 );
xor ( n47406 , n47368 , n47405 );
and ( n47407 , n46208 , n46213 );
and ( n47408 , n46213 , n46219 );
and ( n47409 , n46208 , n46219 );
or ( n47410 , n47407 , n47408 , n47409 );
and ( n47411 , n46217 , n46218 );
not ( n47412 , n1287 );
and ( n47413 , n34193 , n1287 );
nor ( n47414 , n47412 , n47413 );
xor ( n47415 , n47411 , n47414 );
and ( n47416 , n1383 , n32999 );
and ( n47417 , n1580 , n31761 );
xor ( n47418 , n47416 , n47417 );
and ( n47419 , n1694 , n30629 );
xor ( n47420 , n47418 , n47419 );
xor ( n47421 , n47415 , n47420 );
xor ( n47422 , n47410 , n47421 );
xor ( n47423 , n47406 , n47422 );
xor ( n47424 , n47362 , n47423 );
xor ( n47425 , n47282 , n47424 );
xor ( n47426 , n47155 , n47425 );
xor ( n47427 , n47073 , n47426 );
xor ( n47428 , n47064 , n47427 );
and ( n47429 , n45853 , n45856 );
and ( n47430 , n45856 , n46226 );
and ( n47431 , n45853 , n46226 );
or ( n47432 , n47429 , n47430 , n47431 );
xor ( n47433 , n47428 , n47432 );
and ( n47434 , n46227 , n46231 );
and ( n47435 , n46232 , n46235 );
or ( n47436 , n47434 , n47435 );
xor ( n47437 , n47433 , n47436 );
buf ( n47438 , n47437 );
buf ( n47439 , n47438 );
not ( n47440 , n47439 );
nor ( n47441 , n47440 , n8739 );
xor ( n47442 , n47056 , n47441 );
and ( n47443 , n45849 , n46240 );
and ( n47444 , n46241 , n46244 );
or ( n47445 , n47443 , n47444 );
xor ( n47446 , n47442 , n47445 );
buf ( n47447 , n47446 );
buf ( n47448 , n47447 );
not ( n47449 , n47448 );
buf ( n47450 , n573 );
not ( n47451 , n47450 );
nor ( n47452 , n47449 , n47451 );
xor ( n47453 , n46682 , n47452 );
xor ( n47454 , n46256 , n46679 );
nor ( n47455 , n46248 , n47451 );
and ( n47456 , n47454 , n47455 );
xor ( n47457 , n47454 , n47455 );
xor ( n47458 , n46260 , n46677 );
nor ( n47459 , n45047 , n47451 );
and ( n47460 , n47458 , n47459 );
xor ( n47461 , n47458 , n47459 );
xor ( n47462 , n46264 , n46675 );
nor ( n47463 , n43843 , n47451 );
and ( n47464 , n47462 , n47463 );
xor ( n47465 , n47462 , n47463 );
xor ( n47466 , n46268 , n46673 );
nor ( n47467 , n42641 , n47451 );
and ( n47468 , n47466 , n47467 );
xor ( n47469 , n47466 , n47467 );
xor ( n47470 , n46272 , n46671 );
nor ( n47471 , n41437 , n47451 );
and ( n47472 , n47470 , n47471 );
xor ( n47473 , n47470 , n47471 );
xor ( n47474 , n46276 , n46669 );
nor ( n47475 , n40232 , n47451 );
and ( n47476 , n47474 , n47475 );
xor ( n47477 , n47474 , n47475 );
xor ( n47478 , n46280 , n46667 );
nor ( n47479 , n39027 , n47451 );
and ( n47480 , n47478 , n47479 );
xor ( n47481 , n47478 , n47479 );
xor ( n47482 , n46284 , n46665 );
nor ( n47483 , n37825 , n47451 );
and ( n47484 , n47482 , n47483 );
xor ( n47485 , n47482 , n47483 );
xor ( n47486 , n46288 , n46663 );
nor ( n47487 , n36620 , n47451 );
and ( n47488 , n47486 , n47487 );
xor ( n47489 , n47486 , n47487 );
xor ( n47490 , n46292 , n46661 );
nor ( n47491 , n35419 , n47451 );
and ( n47492 , n47490 , n47491 );
xor ( n47493 , n47490 , n47491 );
xor ( n47494 , n46296 , n46659 );
nor ( n47495 , n34224 , n47451 );
and ( n47496 , n47494 , n47495 );
xor ( n47497 , n47494 , n47495 );
xor ( n47498 , n46300 , n46657 );
nor ( n47499 , n33033 , n47451 );
and ( n47500 , n47498 , n47499 );
xor ( n47501 , n47498 , n47499 );
xor ( n47502 , n46304 , n46655 );
nor ( n47503 , n31867 , n47451 );
and ( n47504 , n47502 , n47503 );
xor ( n47505 , n47502 , n47503 );
xor ( n47506 , n46308 , n46653 );
nor ( n47507 , n30725 , n47451 );
and ( n47508 , n47506 , n47507 );
xor ( n47509 , n47506 , n47507 );
xor ( n47510 , n46312 , n46651 );
nor ( n47511 , n29596 , n47451 );
and ( n47512 , n47510 , n47511 );
xor ( n47513 , n47510 , n47511 );
xor ( n47514 , n46316 , n46649 );
nor ( n47515 , n28487 , n47451 );
and ( n47516 , n47514 , n47515 );
xor ( n47517 , n47514 , n47515 );
xor ( n47518 , n46320 , n46647 );
nor ( n47519 , n27397 , n47451 );
and ( n47520 , n47518 , n47519 );
xor ( n47521 , n47518 , n47519 );
xor ( n47522 , n46324 , n46645 );
nor ( n47523 , n26326 , n47451 );
and ( n47524 , n47522 , n47523 );
xor ( n47525 , n47522 , n47523 );
xor ( n47526 , n46328 , n46643 );
nor ( n47527 , n25272 , n47451 );
and ( n47528 , n47526 , n47527 );
xor ( n47529 , n47526 , n47527 );
xor ( n47530 , n46332 , n46641 );
nor ( n47531 , n24242 , n47451 );
and ( n47532 , n47530 , n47531 );
xor ( n47533 , n47530 , n47531 );
xor ( n47534 , n46336 , n46639 );
nor ( n47535 , n23225 , n47451 );
and ( n47536 , n47534 , n47535 );
xor ( n47537 , n47534 , n47535 );
xor ( n47538 , n46340 , n46637 );
nor ( n47539 , n22231 , n47451 );
and ( n47540 , n47538 , n47539 );
xor ( n47541 , n47538 , n47539 );
xor ( n47542 , n46344 , n46635 );
nor ( n47543 , n21258 , n47451 );
and ( n47544 , n47542 , n47543 );
xor ( n47545 , n47542 , n47543 );
xor ( n47546 , n46348 , n46633 );
nor ( n47547 , n20303 , n47451 );
and ( n47548 , n47546 , n47547 );
xor ( n47549 , n47546 , n47547 );
xor ( n47550 , n46352 , n46631 );
nor ( n47551 , n19365 , n47451 );
and ( n47552 , n47550 , n47551 );
xor ( n47553 , n47550 , n47551 );
xor ( n47554 , n46356 , n46629 );
nor ( n47555 , n18448 , n47451 );
and ( n47556 , n47554 , n47555 );
xor ( n47557 , n47554 , n47555 );
xor ( n47558 , n46360 , n46627 );
nor ( n47559 , n17548 , n47451 );
and ( n47560 , n47558 , n47559 );
xor ( n47561 , n47558 , n47559 );
xor ( n47562 , n46364 , n46625 );
nor ( n47563 , n16669 , n47451 );
and ( n47564 , n47562 , n47563 );
xor ( n47565 , n47562 , n47563 );
xor ( n47566 , n46368 , n46623 );
nor ( n47567 , n15809 , n47451 );
and ( n47568 , n47566 , n47567 );
xor ( n47569 , n47566 , n47567 );
xor ( n47570 , n46372 , n46621 );
nor ( n47571 , n14968 , n47451 );
and ( n47572 , n47570 , n47571 );
xor ( n47573 , n47570 , n47571 );
xor ( n47574 , n46376 , n46619 );
nor ( n47575 , n14147 , n47451 );
and ( n47576 , n47574 , n47575 );
xor ( n47577 , n47574 , n47575 );
xor ( n47578 , n46380 , n46617 );
nor ( n47579 , n13349 , n47451 );
and ( n47580 , n47578 , n47579 );
xor ( n47581 , n47578 , n47579 );
xor ( n47582 , n46384 , n46615 );
nor ( n47583 , n12564 , n47451 );
and ( n47584 , n47582 , n47583 );
xor ( n47585 , n47582 , n47583 );
xor ( n47586 , n46388 , n46613 );
nor ( n47587 , n11799 , n47451 );
and ( n47588 , n47586 , n47587 );
xor ( n47589 , n47586 , n47587 );
xor ( n47590 , n46392 , n46611 );
nor ( n47591 , n11050 , n47451 );
and ( n47592 , n47590 , n47591 );
xor ( n47593 , n47590 , n47591 );
xor ( n47594 , n46396 , n46609 );
nor ( n47595 , n10321 , n47451 );
and ( n47596 , n47594 , n47595 );
xor ( n47597 , n47594 , n47595 );
xor ( n47598 , n46400 , n46607 );
nor ( n47599 , n9429 , n47451 );
and ( n47600 , n47598 , n47599 );
xor ( n47601 , n47598 , n47599 );
xor ( n47602 , n46404 , n46605 );
nor ( n47603 , n8949 , n47451 );
and ( n47604 , n47602 , n47603 );
xor ( n47605 , n47602 , n47603 );
xor ( n47606 , n46408 , n46603 );
nor ( n47607 , n9437 , n47451 );
and ( n47608 , n47606 , n47607 );
xor ( n47609 , n47606 , n47607 );
xor ( n47610 , n46412 , n46601 );
nor ( n47611 , n9446 , n47451 );
and ( n47612 , n47610 , n47611 );
xor ( n47613 , n47610 , n47611 );
xor ( n47614 , n46416 , n46599 );
nor ( n47615 , n9455 , n47451 );
and ( n47616 , n47614 , n47615 );
xor ( n47617 , n47614 , n47615 );
xor ( n47618 , n46420 , n46597 );
nor ( n47619 , n9464 , n47451 );
and ( n47620 , n47618 , n47619 );
xor ( n47621 , n47618 , n47619 );
xor ( n47622 , n46424 , n46595 );
nor ( n47623 , n9473 , n47451 );
and ( n47624 , n47622 , n47623 );
xor ( n47625 , n47622 , n47623 );
xor ( n47626 , n46428 , n46593 );
nor ( n47627 , n9482 , n47451 );
and ( n47628 , n47626 , n47627 );
xor ( n47629 , n47626 , n47627 );
xor ( n47630 , n46432 , n46591 );
nor ( n47631 , n9491 , n47451 );
and ( n47632 , n47630 , n47631 );
xor ( n47633 , n47630 , n47631 );
xor ( n47634 , n46436 , n46589 );
nor ( n47635 , n9500 , n47451 );
and ( n47636 , n47634 , n47635 );
xor ( n47637 , n47634 , n47635 );
xor ( n47638 , n46440 , n46587 );
nor ( n47639 , n9509 , n47451 );
and ( n47640 , n47638 , n47639 );
xor ( n47641 , n47638 , n47639 );
xor ( n47642 , n46444 , n46585 );
nor ( n47643 , n9518 , n47451 );
and ( n47644 , n47642 , n47643 );
xor ( n47645 , n47642 , n47643 );
xor ( n47646 , n46448 , n46583 );
nor ( n47647 , n9527 , n47451 );
and ( n47648 , n47646 , n47647 );
xor ( n47649 , n47646 , n47647 );
xor ( n47650 , n46452 , n46581 );
nor ( n47651 , n9536 , n47451 );
and ( n47652 , n47650 , n47651 );
xor ( n47653 , n47650 , n47651 );
xor ( n47654 , n46456 , n46579 );
nor ( n47655 , n9545 , n47451 );
and ( n47656 , n47654 , n47655 );
xor ( n47657 , n47654 , n47655 );
xor ( n47658 , n46460 , n46577 );
nor ( n47659 , n9554 , n47451 );
and ( n47660 , n47658 , n47659 );
xor ( n47661 , n47658 , n47659 );
xor ( n47662 , n46464 , n46575 );
nor ( n47663 , n9563 , n47451 );
and ( n47664 , n47662 , n47663 );
xor ( n47665 , n47662 , n47663 );
xor ( n47666 , n46468 , n46573 );
nor ( n47667 , n9572 , n47451 );
and ( n47668 , n47666 , n47667 );
xor ( n47669 , n47666 , n47667 );
xor ( n47670 , n46472 , n46571 );
nor ( n47671 , n9581 , n47451 );
and ( n47672 , n47670 , n47671 );
xor ( n47673 , n47670 , n47671 );
xor ( n47674 , n46476 , n46569 );
nor ( n47675 , n9590 , n47451 );
and ( n47676 , n47674 , n47675 );
xor ( n47677 , n47674 , n47675 );
xor ( n47678 , n46480 , n46567 );
nor ( n47679 , n9599 , n47451 );
and ( n47680 , n47678 , n47679 );
xor ( n47681 , n47678 , n47679 );
xor ( n47682 , n46484 , n46565 );
nor ( n47683 , n9608 , n47451 );
and ( n47684 , n47682 , n47683 );
xor ( n47685 , n47682 , n47683 );
xor ( n47686 , n46488 , n46563 );
nor ( n47687 , n9617 , n47451 );
and ( n47688 , n47686 , n47687 );
xor ( n47689 , n47686 , n47687 );
xor ( n47690 , n46492 , n46561 );
nor ( n47691 , n9626 , n47451 );
and ( n47692 , n47690 , n47691 );
xor ( n47693 , n47690 , n47691 );
xor ( n47694 , n46496 , n46559 );
nor ( n47695 , n9635 , n47451 );
and ( n47696 , n47694 , n47695 );
xor ( n47697 , n47694 , n47695 );
xor ( n47698 , n46500 , n46557 );
nor ( n47699 , n9644 , n47451 );
and ( n47700 , n47698 , n47699 );
xor ( n47701 , n47698 , n47699 );
xor ( n47702 , n46504 , n46555 );
nor ( n47703 , n9653 , n47451 );
and ( n47704 , n47702 , n47703 );
xor ( n47705 , n47702 , n47703 );
xor ( n47706 , n46508 , n46553 );
nor ( n47707 , n9662 , n47451 );
and ( n47708 , n47706 , n47707 );
xor ( n47709 , n47706 , n47707 );
xor ( n47710 , n46512 , n46551 );
nor ( n47711 , n9671 , n47451 );
and ( n47712 , n47710 , n47711 );
xor ( n47713 , n47710 , n47711 );
xor ( n47714 , n46516 , n46549 );
nor ( n47715 , n9680 , n47451 );
and ( n47716 , n47714 , n47715 );
xor ( n47717 , n47714 , n47715 );
xor ( n47718 , n46520 , n46547 );
nor ( n47719 , n9689 , n47451 );
and ( n47720 , n47718 , n47719 );
xor ( n47721 , n47718 , n47719 );
xor ( n47722 , n46524 , n46545 );
nor ( n47723 , n9698 , n47451 );
and ( n47724 , n47722 , n47723 );
xor ( n47725 , n47722 , n47723 );
xor ( n47726 , n46528 , n46543 );
nor ( n47727 , n9707 , n47451 );
and ( n47728 , n47726 , n47727 );
xor ( n47729 , n47726 , n47727 );
xor ( n47730 , n46532 , n46541 );
nor ( n47731 , n9716 , n47451 );
and ( n47732 , n47730 , n47731 );
xor ( n47733 , n47730 , n47731 );
xor ( n47734 , n46536 , n46539 );
nor ( n47735 , n9725 , n47451 );
and ( n47736 , n47734 , n47735 );
xor ( n47737 , n47734 , n47735 );
xor ( n47738 , n46537 , n46538 );
nor ( n47739 , n9734 , n47451 );
and ( n47740 , n47738 , n47739 );
xor ( n47741 , n47738 , n47739 );
nor ( n47742 , n9752 , n46250 );
nor ( n47743 , n9743 , n47451 );
and ( n47744 , n47742 , n47743 );
and ( n47745 , n47741 , n47744 );
or ( n47746 , n47740 , n47745 );
and ( n47747 , n47737 , n47746 );
or ( n47748 , n47736 , n47747 );
and ( n47749 , n47733 , n47748 );
or ( n47750 , n47732 , n47749 );
and ( n47751 , n47729 , n47750 );
or ( n47752 , n47728 , n47751 );
and ( n47753 , n47725 , n47752 );
or ( n47754 , n47724 , n47753 );
and ( n47755 , n47721 , n47754 );
or ( n47756 , n47720 , n47755 );
and ( n47757 , n47717 , n47756 );
or ( n47758 , n47716 , n47757 );
and ( n47759 , n47713 , n47758 );
or ( n47760 , n47712 , n47759 );
and ( n47761 , n47709 , n47760 );
or ( n47762 , n47708 , n47761 );
and ( n47763 , n47705 , n47762 );
or ( n47764 , n47704 , n47763 );
and ( n47765 , n47701 , n47764 );
or ( n47766 , n47700 , n47765 );
and ( n47767 , n47697 , n47766 );
or ( n47768 , n47696 , n47767 );
and ( n47769 , n47693 , n47768 );
or ( n47770 , n47692 , n47769 );
and ( n47771 , n47689 , n47770 );
or ( n47772 , n47688 , n47771 );
and ( n47773 , n47685 , n47772 );
or ( n47774 , n47684 , n47773 );
and ( n47775 , n47681 , n47774 );
or ( n47776 , n47680 , n47775 );
and ( n47777 , n47677 , n47776 );
or ( n47778 , n47676 , n47777 );
and ( n47779 , n47673 , n47778 );
or ( n47780 , n47672 , n47779 );
and ( n47781 , n47669 , n47780 );
or ( n47782 , n47668 , n47781 );
and ( n47783 , n47665 , n47782 );
or ( n47784 , n47664 , n47783 );
and ( n47785 , n47661 , n47784 );
or ( n47786 , n47660 , n47785 );
and ( n47787 , n47657 , n47786 );
or ( n47788 , n47656 , n47787 );
and ( n47789 , n47653 , n47788 );
or ( n47790 , n47652 , n47789 );
and ( n47791 , n47649 , n47790 );
or ( n47792 , n47648 , n47791 );
and ( n47793 , n47645 , n47792 );
or ( n47794 , n47644 , n47793 );
and ( n47795 , n47641 , n47794 );
or ( n47796 , n47640 , n47795 );
and ( n47797 , n47637 , n47796 );
or ( n47798 , n47636 , n47797 );
and ( n47799 , n47633 , n47798 );
or ( n47800 , n47632 , n47799 );
and ( n47801 , n47629 , n47800 );
or ( n47802 , n47628 , n47801 );
and ( n47803 , n47625 , n47802 );
or ( n47804 , n47624 , n47803 );
and ( n47805 , n47621 , n47804 );
or ( n47806 , n47620 , n47805 );
and ( n47807 , n47617 , n47806 );
or ( n47808 , n47616 , n47807 );
and ( n47809 , n47613 , n47808 );
or ( n47810 , n47612 , n47809 );
and ( n47811 , n47609 , n47810 );
or ( n47812 , n47608 , n47811 );
and ( n47813 , n47605 , n47812 );
or ( n47814 , n47604 , n47813 );
and ( n47815 , n47601 , n47814 );
or ( n47816 , n47600 , n47815 );
and ( n47817 , n47597 , n47816 );
or ( n47818 , n47596 , n47817 );
and ( n47819 , n47593 , n47818 );
or ( n47820 , n47592 , n47819 );
and ( n47821 , n47589 , n47820 );
or ( n47822 , n47588 , n47821 );
and ( n47823 , n47585 , n47822 );
or ( n47824 , n47584 , n47823 );
and ( n47825 , n47581 , n47824 );
or ( n47826 , n47580 , n47825 );
and ( n47827 , n47577 , n47826 );
or ( n47828 , n47576 , n47827 );
and ( n47829 , n47573 , n47828 );
or ( n47830 , n47572 , n47829 );
and ( n47831 , n47569 , n47830 );
or ( n47832 , n47568 , n47831 );
and ( n47833 , n47565 , n47832 );
or ( n47834 , n47564 , n47833 );
and ( n47835 , n47561 , n47834 );
or ( n47836 , n47560 , n47835 );
and ( n47837 , n47557 , n47836 );
or ( n47838 , n47556 , n47837 );
and ( n47839 , n47553 , n47838 );
or ( n47840 , n47552 , n47839 );
and ( n47841 , n47549 , n47840 );
or ( n47842 , n47548 , n47841 );
and ( n47843 , n47545 , n47842 );
or ( n47844 , n47544 , n47843 );
and ( n47845 , n47541 , n47844 );
or ( n47846 , n47540 , n47845 );
and ( n47847 , n47537 , n47846 );
or ( n47848 , n47536 , n47847 );
and ( n47849 , n47533 , n47848 );
or ( n47850 , n47532 , n47849 );
and ( n47851 , n47529 , n47850 );
or ( n47852 , n47528 , n47851 );
and ( n47853 , n47525 , n47852 );
or ( n47854 , n47524 , n47853 );
and ( n47855 , n47521 , n47854 );
or ( n47856 , n47520 , n47855 );
and ( n47857 , n47517 , n47856 );
or ( n47858 , n47516 , n47857 );
and ( n47859 , n47513 , n47858 );
or ( n47860 , n47512 , n47859 );
and ( n47861 , n47509 , n47860 );
or ( n47862 , n47508 , n47861 );
and ( n47863 , n47505 , n47862 );
or ( n47864 , n47504 , n47863 );
and ( n47865 , n47501 , n47864 );
or ( n47866 , n47500 , n47865 );
and ( n47867 , n47497 , n47866 );
or ( n47868 , n47496 , n47867 );
and ( n47869 , n47493 , n47868 );
or ( n47870 , n47492 , n47869 );
and ( n47871 , n47489 , n47870 );
or ( n47872 , n47488 , n47871 );
and ( n47873 , n47485 , n47872 );
or ( n47874 , n47484 , n47873 );
and ( n47875 , n47481 , n47874 );
or ( n47876 , n47480 , n47875 );
and ( n47877 , n47477 , n47876 );
or ( n47878 , n47476 , n47877 );
and ( n47879 , n47473 , n47878 );
or ( n47880 , n47472 , n47879 );
and ( n47881 , n47469 , n47880 );
or ( n47882 , n47468 , n47881 );
and ( n47883 , n47465 , n47882 );
or ( n47884 , n47464 , n47883 );
and ( n47885 , n47461 , n47884 );
or ( n47886 , n47460 , n47885 );
and ( n47887 , n47457 , n47886 );
or ( n47888 , n47456 , n47887 );
xor ( n47889 , n47453 , n47888 );
and ( n47890 , n33403 , n1444 );
nor ( n47891 , n1445 , n47890 );
nor ( n47892 , n1598 , n32231 );
xor ( n47893 , n47891 , n47892 );
and ( n47894 , n46684 , n46685 );
and ( n47895 , n46686 , n46689 );
or ( n47896 , n47894 , n47895 );
xor ( n47897 , n47893 , n47896 );
nor ( n47898 , n1766 , n31083 );
xor ( n47899 , n47897 , n47898 );
and ( n47900 , n46690 , n46691 );
and ( n47901 , n46692 , n46695 );
or ( n47902 , n47900 , n47901 );
xor ( n47903 , n47899 , n47902 );
nor ( n47904 , n1945 , n29948 );
xor ( n47905 , n47903 , n47904 );
and ( n47906 , n46696 , n46697 );
and ( n47907 , n46698 , n46701 );
or ( n47908 , n47906 , n47907 );
xor ( n47909 , n47905 , n47908 );
nor ( n47910 , n2137 , n28833 );
xor ( n47911 , n47909 , n47910 );
and ( n47912 , n46702 , n46703 );
and ( n47913 , n46704 , n46707 );
or ( n47914 , n47912 , n47913 );
xor ( n47915 , n47911 , n47914 );
nor ( n47916 , n2343 , n27737 );
xor ( n47917 , n47915 , n47916 );
and ( n47918 , n46708 , n46709 );
and ( n47919 , n46710 , n46713 );
or ( n47920 , n47918 , n47919 );
xor ( n47921 , n47917 , n47920 );
nor ( n47922 , n2566 , n26660 );
xor ( n47923 , n47921 , n47922 );
and ( n47924 , n46714 , n46715 );
and ( n47925 , n46716 , n46719 );
or ( n47926 , n47924 , n47925 );
xor ( n47927 , n47923 , n47926 );
nor ( n47928 , n2797 , n25600 );
xor ( n47929 , n47927 , n47928 );
and ( n47930 , n46720 , n46721 );
and ( n47931 , n46722 , n46725 );
or ( n47932 , n47930 , n47931 );
xor ( n47933 , n47929 , n47932 );
nor ( n47934 , n3043 , n24564 );
xor ( n47935 , n47933 , n47934 );
and ( n47936 , n46726 , n46727 );
and ( n47937 , n46728 , n46731 );
or ( n47938 , n47936 , n47937 );
xor ( n47939 , n47935 , n47938 );
nor ( n47940 , n3300 , n23541 );
xor ( n47941 , n47939 , n47940 );
and ( n47942 , n46732 , n46733 );
and ( n47943 , n46734 , n46737 );
or ( n47944 , n47942 , n47943 );
xor ( n47945 , n47941 , n47944 );
nor ( n47946 , n3570 , n22541 );
xor ( n47947 , n47945 , n47946 );
and ( n47948 , n46738 , n46739 );
and ( n47949 , n46740 , n46743 );
or ( n47950 , n47948 , n47949 );
xor ( n47951 , n47947 , n47950 );
nor ( n47952 , n3853 , n21562 );
xor ( n47953 , n47951 , n47952 );
and ( n47954 , n46744 , n46745 );
and ( n47955 , n46746 , n46749 );
or ( n47956 , n47954 , n47955 );
xor ( n47957 , n47953 , n47956 );
nor ( n47958 , n4151 , n20601 );
xor ( n47959 , n47957 , n47958 );
and ( n47960 , n46750 , n46751 );
and ( n47961 , n46752 , n46755 );
or ( n47962 , n47960 , n47961 );
xor ( n47963 , n47959 , n47962 );
nor ( n47964 , n4458 , n19657 );
xor ( n47965 , n47963 , n47964 );
and ( n47966 , n46756 , n46757 );
and ( n47967 , n46758 , n46761 );
or ( n47968 , n47966 , n47967 );
xor ( n47969 , n47965 , n47968 );
nor ( n47970 , n4786 , n18734 );
xor ( n47971 , n47969 , n47970 );
and ( n47972 , n46762 , n46763 );
and ( n47973 , n46764 , n46767 );
or ( n47974 , n47972 , n47973 );
xor ( n47975 , n47971 , n47974 );
nor ( n47976 , n5126 , n17828 );
xor ( n47977 , n47975 , n47976 );
and ( n47978 , n46768 , n46769 );
and ( n47979 , n46770 , n46773 );
or ( n47980 , n47978 , n47979 );
xor ( n47981 , n47977 , n47980 );
nor ( n47982 , n5477 , n16943 );
xor ( n47983 , n47981 , n47982 );
and ( n47984 , n46774 , n46775 );
and ( n47985 , n46776 , n46779 );
or ( n47986 , n47984 , n47985 );
xor ( n47987 , n47983 , n47986 );
nor ( n47988 , n5838 , n16077 );
xor ( n47989 , n47987 , n47988 );
and ( n47990 , n46780 , n46781 );
and ( n47991 , n46782 , n46785 );
or ( n47992 , n47990 , n47991 );
xor ( n47993 , n47989 , n47992 );
nor ( n47994 , n6212 , n15230 );
xor ( n47995 , n47993 , n47994 );
and ( n47996 , n46786 , n46787 );
and ( n47997 , n46788 , n46791 );
or ( n47998 , n47996 , n47997 );
xor ( n47999 , n47995 , n47998 );
nor ( n48000 , n6596 , n14403 );
xor ( n48001 , n47999 , n48000 );
and ( n48002 , n46792 , n46793 );
and ( n48003 , n46794 , n46797 );
or ( n48004 , n48002 , n48003 );
xor ( n48005 , n48001 , n48004 );
nor ( n48006 , n6997 , n13599 );
xor ( n48007 , n48005 , n48006 );
and ( n48008 , n46798 , n46799 );
and ( n48009 , n46800 , n46803 );
or ( n48010 , n48008 , n48009 );
xor ( n48011 , n48007 , n48010 );
nor ( n48012 , n7413 , n12808 );
xor ( n48013 , n48011 , n48012 );
and ( n48014 , n46804 , n46805 );
and ( n48015 , n46806 , n46809 );
or ( n48016 , n48014 , n48015 );
xor ( n48017 , n48013 , n48016 );
nor ( n48018 , n7841 , n12037 );
xor ( n48019 , n48017 , n48018 );
and ( n48020 , n46810 , n46811 );
and ( n48021 , n46812 , n46815 );
or ( n48022 , n48020 , n48021 );
xor ( n48023 , n48019 , n48022 );
nor ( n48024 , n8281 , n11282 );
xor ( n48025 , n48023 , n48024 );
and ( n48026 , n46816 , n46817 );
and ( n48027 , n46818 , n46821 );
or ( n48028 , n48026 , n48027 );
xor ( n48029 , n48025 , n48028 );
nor ( n48030 , n8737 , n10547 );
xor ( n48031 , n48029 , n48030 );
and ( n48032 , n46822 , n46823 );
and ( n48033 , n46824 , n46827 );
or ( n48034 , n48032 , n48033 );
xor ( n48035 , n48031 , n48034 );
nor ( n48036 , n9420 , n9829 );
xor ( n48037 , n48035 , n48036 );
and ( n48038 , n46828 , n46829 );
and ( n48039 , n46830 , n46833 );
or ( n48040 , n48038 , n48039 );
xor ( n48041 , n48037 , n48040 );
nor ( n48042 , n10312 , n8955 );
xor ( n48043 , n48041 , n48042 );
and ( n48044 , n46834 , n46835 );
and ( n48045 , n46836 , n46839 );
or ( n48046 , n48044 , n48045 );
xor ( n48047 , n48043 , n48046 );
nor ( n48048 , n11041 , n603 );
xor ( n48049 , n48047 , n48048 );
and ( n48050 , n46840 , n46841 );
and ( n48051 , n46842 , n46845 );
or ( n48052 , n48050 , n48051 );
xor ( n48053 , n48049 , n48052 );
nor ( n48054 , n11790 , n652 );
xor ( n48055 , n48053 , n48054 );
and ( n48056 , n46846 , n46847 );
and ( n48057 , n46848 , n46851 );
or ( n48058 , n48056 , n48057 );
xor ( n48059 , n48055 , n48058 );
nor ( n48060 , n12555 , n624 );
xor ( n48061 , n48059 , n48060 );
and ( n48062 , n46852 , n46853 );
and ( n48063 , n46854 , n46857 );
or ( n48064 , n48062 , n48063 );
xor ( n48065 , n48061 , n48064 );
nor ( n48066 , n13340 , n648 );
xor ( n48067 , n48065 , n48066 );
and ( n48068 , n46858 , n46859 );
and ( n48069 , n46860 , n46863 );
or ( n48070 , n48068 , n48069 );
xor ( n48071 , n48067 , n48070 );
nor ( n48072 , n14138 , n686 );
xor ( n48073 , n48071 , n48072 );
and ( n48074 , n46864 , n46865 );
and ( n48075 , n46866 , n46869 );
or ( n48076 , n48074 , n48075 );
xor ( n48077 , n48073 , n48076 );
nor ( n48078 , n14959 , n735 );
xor ( n48079 , n48077 , n48078 );
and ( n48080 , n46870 , n46871 );
and ( n48081 , n46872 , n46875 );
or ( n48082 , n48080 , n48081 );
xor ( n48083 , n48079 , n48082 );
nor ( n48084 , n15800 , n798 );
xor ( n48085 , n48083 , n48084 );
and ( n48086 , n46876 , n46877 );
and ( n48087 , n46878 , n46881 );
or ( n48088 , n48086 , n48087 );
xor ( n48089 , n48085 , n48088 );
nor ( n48090 , n16660 , n870 );
xor ( n48091 , n48089 , n48090 );
and ( n48092 , n46882 , n46883 );
and ( n48093 , n46884 , n46887 );
or ( n48094 , n48092 , n48093 );
xor ( n48095 , n48091 , n48094 );
nor ( n48096 , n17539 , n960 );
xor ( n48097 , n48095 , n48096 );
and ( n48098 , n46888 , n46889 );
and ( n48099 , n46890 , n46893 );
or ( n48100 , n48098 , n48099 );
xor ( n48101 , n48097 , n48100 );
nor ( n48102 , n18439 , n1064 );
xor ( n48103 , n48101 , n48102 );
and ( n48104 , n46894 , n46895 );
and ( n48105 , n46896 , n46899 );
or ( n48106 , n48104 , n48105 );
xor ( n48107 , n48103 , n48106 );
nor ( n48108 , n19356 , n1178 );
xor ( n48109 , n48107 , n48108 );
and ( n48110 , n46900 , n46901 );
and ( n48111 , n46902 , n46905 );
or ( n48112 , n48110 , n48111 );
xor ( n48113 , n48109 , n48112 );
nor ( n48114 , n20294 , n1305 );
xor ( n48115 , n48113 , n48114 );
and ( n48116 , n46906 , n46907 );
and ( n48117 , n46908 , n46911 );
or ( n48118 , n48116 , n48117 );
xor ( n48119 , n48115 , n48118 );
nor ( n48120 , n21249 , n1447 );
xor ( n48121 , n48119 , n48120 );
and ( n48122 , n46912 , n46913 );
and ( n48123 , n46914 , n46917 );
or ( n48124 , n48122 , n48123 );
xor ( n48125 , n48121 , n48124 );
nor ( n48126 , n22222 , n1600 );
xor ( n48127 , n48125 , n48126 );
and ( n48128 , n46918 , n46919 );
and ( n48129 , n46920 , n46923 );
or ( n48130 , n48128 , n48129 );
xor ( n48131 , n48127 , n48130 );
nor ( n48132 , n23216 , n1768 );
xor ( n48133 , n48131 , n48132 );
and ( n48134 , n46924 , n46925 );
and ( n48135 , n46926 , n46929 );
or ( n48136 , n48134 , n48135 );
xor ( n48137 , n48133 , n48136 );
nor ( n48138 , n24233 , n1947 );
xor ( n48139 , n48137 , n48138 );
and ( n48140 , n46930 , n46931 );
and ( n48141 , n46932 , n46935 );
or ( n48142 , n48140 , n48141 );
xor ( n48143 , n48139 , n48142 );
nor ( n48144 , n25263 , n2139 );
xor ( n48145 , n48143 , n48144 );
and ( n48146 , n46936 , n46937 );
and ( n48147 , n46938 , n46941 );
or ( n48148 , n48146 , n48147 );
xor ( n48149 , n48145 , n48148 );
nor ( n48150 , n26317 , n2345 );
xor ( n48151 , n48149 , n48150 );
and ( n48152 , n46942 , n46943 );
and ( n48153 , n46944 , n46947 );
or ( n48154 , n48152 , n48153 );
xor ( n48155 , n48151 , n48154 );
nor ( n48156 , n27388 , n2568 );
xor ( n48157 , n48155 , n48156 );
and ( n48158 , n46948 , n46949 );
and ( n48159 , n46950 , n46953 );
or ( n48160 , n48158 , n48159 );
xor ( n48161 , n48157 , n48160 );
nor ( n48162 , n28478 , n2799 );
xor ( n48163 , n48161 , n48162 );
and ( n48164 , n46954 , n46955 );
and ( n48165 , n46956 , n46959 );
or ( n48166 , n48164 , n48165 );
xor ( n48167 , n48163 , n48166 );
nor ( n48168 , n29587 , n3045 );
xor ( n48169 , n48167 , n48168 );
and ( n48170 , n46960 , n46961 );
and ( n48171 , n46962 , n46965 );
or ( n48172 , n48170 , n48171 );
xor ( n48173 , n48169 , n48172 );
nor ( n48174 , n30716 , n3302 );
xor ( n48175 , n48173 , n48174 );
and ( n48176 , n46966 , n46967 );
and ( n48177 , n46968 , n46971 );
or ( n48178 , n48176 , n48177 );
xor ( n48179 , n48175 , n48178 );
nor ( n48180 , n31858 , n3572 );
xor ( n48181 , n48179 , n48180 );
and ( n48182 , n46972 , n46973 );
and ( n48183 , n46974 , n46977 );
or ( n48184 , n48182 , n48183 );
xor ( n48185 , n48181 , n48184 );
nor ( n48186 , n33024 , n3855 );
xor ( n48187 , n48185 , n48186 );
and ( n48188 , n46978 , n46979 );
and ( n48189 , n46980 , n46983 );
or ( n48190 , n48188 , n48189 );
xor ( n48191 , n48187 , n48190 );
nor ( n48192 , n34215 , n4153 );
xor ( n48193 , n48191 , n48192 );
and ( n48194 , n46984 , n46985 );
and ( n48195 , n46986 , n46989 );
or ( n48196 , n48194 , n48195 );
xor ( n48197 , n48193 , n48196 );
nor ( n48198 , n35410 , n4460 );
xor ( n48199 , n48197 , n48198 );
and ( n48200 , n46990 , n46991 );
and ( n48201 , n46992 , n46995 );
or ( n48202 , n48200 , n48201 );
xor ( n48203 , n48199 , n48202 );
nor ( n48204 , n36611 , n4788 );
xor ( n48205 , n48203 , n48204 );
and ( n48206 , n46996 , n46997 );
and ( n48207 , n46998 , n47001 );
or ( n48208 , n48206 , n48207 );
xor ( n48209 , n48205 , n48208 );
nor ( n48210 , n37816 , n5128 );
xor ( n48211 , n48209 , n48210 );
and ( n48212 , n47002 , n47003 );
and ( n48213 , n47004 , n47007 );
or ( n48214 , n48212 , n48213 );
xor ( n48215 , n48211 , n48214 );
nor ( n48216 , n39018 , n5479 );
xor ( n48217 , n48215 , n48216 );
and ( n48218 , n47008 , n47009 );
and ( n48219 , n47010 , n47013 );
or ( n48220 , n48218 , n48219 );
xor ( n48221 , n48217 , n48220 );
nor ( n48222 , n40223 , n5840 );
xor ( n48223 , n48221 , n48222 );
and ( n48224 , n47014 , n47015 );
and ( n48225 , n47016 , n47019 );
or ( n48226 , n48224 , n48225 );
xor ( n48227 , n48223 , n48226 );
nor ( n48228 , n41428 , n6214 );
xor ( n48229 , n48227 , n48228 );
and ( n48230 , n47020 , n47021 );
and ( n48231 , n47022 , n47025 );
or ( n48232 , n48230 , n48231 );
xor ( n48233 , n48229 , n48232 );
nor ( n48234 , n42632 , n6598 );
xor ( n48235 , n48233 , n48234 );
and ( n48236 , n47026 , n47027 );
and ( n48237 , n47028 , n47031 );
or ( n48238 , n48236 , n48237 );
xor ( n48239 , n48235 , n48238 );
nor ( n48240 , n43834 , n6999 );
xor ( n48241 , n48239 , n48240 );
and ( n48242 , n47032 , n47033 );
and ( n48243 , n47034 , n47037 );
or ( n48244 , n48242 , n48243 );
xor ( n48245 , n48241 , n48244 );
nor ( n48246 , n45038 , n7415 );
xor ( n48247 , n48245 , n48246 );
and ( n48248 , n47038 , n47039 );
and ( n48249 , n47040 , n47043 );
or ( n48250 , n48248 , n48249 );
xor ( n48251 , n48247 , n48250 );
nor ( n48252 , n46239 , n7843 );
xor ( n48253 , n48251 , n48252 );
and ( n48254 , n47044 , n47045 );
and ( n48255 , n47046 , n47049 );
or ( n48256 , n48254 , n48255 );
xor ( n48257 , n48253 , n48256 );
nor ( n48258 , n47440 , n8283 );
xor ( n48259 , n48257 , n48258 );
and ( n48260 , n47050 , n47051 );
and ( n48261 , n47052 , n47055 );
or ( n48262 , n48260 , n48261 );
xor ( n48263 , n48259 , n48262 );
and ( n48264 , n47068 , n47072 );
and ( n48265 , n47072 , n47426 );
and ( n48266 , n47068 , n47426 );
or ( n48267 , n48264 , n48265 , n48266 );
and ( n48268 , n33774 , n1424 );
not ( n48269 , n1424 );
nor ( n48270 , n48268 , n48269 );
xor ( n48271 , n48267 , n48270 );
and ( n48272 , n47081 , n47085 );
and ( n48273 , n47085 , n47153 );
and ( n48274 , n47081 , n47153 );
or ( n48275 , n48272 , n48273 , n48274 );
and ( n48276 , n47077 , n47154 );
and ( n48277 , n47154 , n47425 );
and ( n48278 , n47077 , n47425 );
or ( n48279 , n48276 , n48277 , n48278 );
xor ( n48280 , n48275 , n48279 );
and ( n48281 , n47159 , n47281 );
and ( n48282 , n47281 , n47424 );
and ( n48283 , n47159 , n47424 );
or ( n48284 , n48281 , n48282 , n48283 );
and ( n48285 , n47090 , n47094 );
and ( n48286 , n47094 , n47152 );
and ( n48287 , n47090 , n47152 );
or ( n48288 , n48285 , n48286 , n48287 );
and ( n48289 , n47163 , n47167 );
and ( n48290 , n47167 , n47280 );
and ( n48291 , n47163 , n47280 );
or ( n48292 , n48289 , n48290 , n48291 );
xor ( n48293 , n48288 , n48292 );
and ( n48294 , n47121 , n47125 );
and ( n48295 , n47125 , n47131 );
and ( n48296 , n47121 , n47131 );
or ( n48297 , n48294 , n48295 , n48296 );
and ( n48298 , n47099 , n47103 );
and ( n48299 , n47103 , n47151 );
and ( n48300 , n47099 , n47151 );
or ( n48301 , n48298 , n48299 , n48300 );
xor ( n48302 , n48297 , n48301 );
and ( n48303 , n47108 , n47112 );
and ( n48304 , n47112 , n47150 );
and ( n48305 , n47108 , n47150 );
or ( n48306 , n48303 , n48304 , n48305 );
and ( n48307 , n47176 , n47201 );
and ( n48308 , n47201 , n47239 );
and ( n48309 , n47176 , n47239 );
or ( n48310 , n48307 , n48308 , n48309 );
xor ( n48311 , n48306 , n48310 );
and ( n48312 , n47117 , n47132 );
and ( n48313 , n47132 , n47149 );
and ( n48314 , n47117 , n47149 );
or ( n48315 , n48312 , n48313 , n48314 );
and ( n48316 , n47180 , n47184 );
and ( n48317 , n47184 , n47200 );
and ( n48318 , n47180 , n47200 );
or ( n48319 , n48316 , n48317 , n48318 );
xor ( n48320 , n48315 , n48319 );
and ( n48321 , n47137 , n47142 );
and ( n48322 , n47142 , n47148 );
and ( n48323 , n47137 , n47148 );
or ( n48324 , n48321 , n48322 , n48323 );
and ( n48325 , n47127 , n47128 );
and ( n48326 , n47128 , n47130 );
and ( n48327 , n47127 , n47130 );
or ( n48328 , n48325 , n48326 , n48327 );
and ( n48329 , n47138 , n47139 );
and ( n48330 , n47139 , n47141 );
and ( n48331 , n47138 , n47141 );
or ( n48332 , n48329 , n48330 , n48331 );
xor ( n48333 , n48328 , n48332 );
and ( n48334 , n30695 , n1882 );
and ( n48335 , n31836 , n1738 );
xor ( n48336 , n48334 , n48335 );
and ( n48337 , n32649 , n1551 );
xor ( n48338 , n48336 , n48337 );
xor ( n48339 , n48333 , n48338 );
xor ( n48340 , n48324 , n48339 );
and ( n48341 , n47144 , n47145 );
and ( n48342 , n47145 , n47147 );
and ( n48343 , n47144 , n47147 );
or ( n48344 , n48341 , n48342 , n48343 );
and ( n48345 , n27361 , n2544 );
and ( n48346 , n28456 , n2298 );
xor ( n48347 , n48345 , n48346 );
and ( n48348 , n29559 , n2100 );
xor ( n48349 , n48347 , n48348 );
xor ( n48350 , n48344 , n48349 );
and ( n48351 , n24214 , n3271 );
and ( n48352 , n25243 , n2981 );
xor ( n48353 , n48351 , n48352 );
and ( n48354 , n26296 , n2739 );
xor ( n48355 , n48353 , n48354 );
xor ( n48356 , n48350 , n48355 );
xor ( n48357 , n48340 , n48356 );
xor ( n48358 , n48320 , n48357 );
xor ( n48359 , n48311 , n48358 );
xor ( n48360 , n48302 , n48359 );
xor ( n48361 , n48293 , n48360 );
xor ( n48362 , n48284 , n48361 );
and ( n48363 , n47283 , n47361 );
and ( n48364 , n47361 , n47423 );
and ( n48365 , n47283 , n47423 );
or ( n48366 , n48363 , n48364 , n48365 );
and ( n48367 , n47172 , n47240 );
and ( n48368 , n47240 , n47279 );
and ( n48369 , n47172 , n47279 );
or ( n48370 , n48367 , n48368 , n48369 );
and ( n48371 , n47287 , n47291 );
and ( n48372 , n47291 , n47360 );
and ( n48373 , n47287 , n47360 );
or ( n48374 , n48371 , n48372 , n48373 );
xor ( n48375 , n48370 , n48374 );
and ( n48376 , n47245 , n47249 );
and ( n48377 , n47249 , n47278 );
and ( n48378 , n47245 , n47278 );
or ( n48379 , n48376 , n48377 , n48378 );
and ( n48380 , n47206 , n47222 );
and ( n48381 , n47222 , n47238 );
and ( n48382 , n47206 , n47238 );
or ( n48383 , n48380 , n48381 , n48382 );
and ( n48384 , n47189 , n47193 );
and ( n48385 , n47193 , n47199 );
and ( n48386 , n47189 , n47199 );
or ( n48387 , n48384 , n48385 , n48386 );
and ( n48388 , n47210 , n47215 );
and ( n48389 , n47215 , n47221 );
and ( n48390 , n47210 , n47221 );
or ( n48391 , n48388 , n48389 , n48390 );
xor ( n48392 , n48387 , n48391 );
and ( n48393 , n47195 , n47196 );
and ( n48394 , n47196 , n47198 );
and ( n48395 , n47195 , n47198 );
or ( n48396 , n48393 , n48394 , n48395 );
and ( n48397 , n47211 , n47212 );
and ( n48398 , n47212 , n47214 );
and ( n48399 , n47211 , n47214 );
or ( n48400 , n48397 , n48398 , n48399 );
xor ( n48401 , n48396 , n48400 );
and ( n48402 , n21216 , n4102 );
and ( n48403 , n22186 , n3749 );
xor ( n48404 , n48402 , n48403 );
and ( n48405 , n22892 , n3495 );
xor ( n48406 , n48404 , n48405 );
xor ( n48407 , n48401 , n48406 );
xor ( n48408 , n48392 , n48407 );
xor ( n48409 , n48383 , n48408 );
and ( n48410 , n47227 , n47231 );
and ( n48411 , n47231 , n47237 );
and ( n48412 , n47227 , n47237 );
or ( n48413 , n48410 , n48411 , n48412 );
and ( n48414 , n47217 , n47218 );
and ( n48415 , n47218 , n47220 );
and ( n48416 , n47217 , n47220 );
or ( n48417 , n48414 , n48415 , n48416 );
and ( n48418 , n18144 , n5103 );
and ( n48419 , n19324 , n4730 );
xor ( n48420 , n48418 , n48419 );
and ( n48421 , n20233 , n4403 );
xor ( n48422 , n48420 , n48421 );
xor ( n48423 , n48417 , n48422 );
and ( n48424 , n15758 , n6132 );
and ( n48425 , n16637 , n5765 );
xor ( n48426 , n48424 , n48425 );
and ( n48427 , n17512 , n5408 );
xor ( n48428 , n48426 , n48427 );
xor ( n48429 , n48423 , n48428 );
xor ( n48430 , n48413 , n48429 );
and ( n48431 , n47233 , n47234 );
and ( n48432 , n47234 , n47236 );
and ( n48433 , n47233 , n47236 );
or ( n48434 , n48431 , n48432 , n48433 );
and ( n48435 , n47266 , n47267 );
and ( n48436 , n47267 , n47269 );
and ( n48437 , n47266 , n47269 );
or ( n48438 , n48435 , n48436 , n48437 );
xor ( n48439 , n48434 , n48438 );
and ( n48440 , n13322 , n7310 );
and ( n48441 , n14118 , n6971 );
xor ( n48442 , n48440 , n48441 );
and ( n48443 , n14938 , n6504 );
xor ( n48444 , n48442 , n48443 );
xor ( n48445 , n48439 , n48444 );
xor ( n48446 , n48430 , n48445 );
xor ( n48447 , n48409 , n48446 );
xor ( n48448 , n48379 , n48447 );
and ( n48449 , n47254 , n47258 );
and ( n48450 , n47258 , n47277 );
and ( n48451 , n47254 , n47277 );
or ( n48452 , n48449 , n48450 , n48451 );
and ( n48453 , n47300 , n47315 );
and ( n48454 , n47315 , n47332 );
and ( n48455 , n47300 , n47332 );
or ( n48456 , n48453 , n48454 , n48455 );
xor ( n48457 , n48452 , n48456 );
and ( n48458 , n47265 , n47270 );
and ( n48459 , n47270 , n47276 );
and ( n48460 , n47265 , n47276 );
or ( n48461 , n48458 , n48459 , n48460 );
and ( n48462 , n47304 , n47308 );
and ( n48463 , n47308 , n47314 );
and ( n48464 , n47304 , n47314 );
or ( n48465 , n48462 , n48463 , n48464 );
xor ( n48466 , n48461 , n48465 );
and ( n48467 , n47272 , n47273 );
and ( n48468 , n47273 , n47275 );
and ( n48469 , n47272 , n47275 );
or ( n48470 , n48467 , n48468 , n48469 );
and ( n48471 , n11015 , n8669 );
and ( n48472 , n11769 , n8243 );
xor ( n48473 , n48471 , n48472 );
and ( n48474 , n12320 , n7662 );
xor ( n48475 , n48473 , n48474 );
xor ( n48476 , n48470 , n48475 );
and ( n48477 , n8718 , n10977 );
and ( n48478 , n9400 , n10239 );
xor ( n48479 , n48477 , n48478 );
and ( n48480 , n10291 , n9348 );
xor ( n48481 , n48479 , n48480 );
xor ( n48482 , n48476 , n48481 );
xor ( n48483 , n48466 , n48482 );
xor ( n48484 , n48457 , n48483 );
xor ( n48485 , n48448 , n48484 );
xor ( n48486 , n48375 , n48485 );
xor ( n48487 , n48366 , n48486 );
and ( n48488 , n47406 , n47422 );
and ( n48489 , n47366 , n47367 );
and ( n48490 , n47367 , n47405 );
and ( n48491 , n47366 , n47405 );
or ( n48492 , n48489 , n48490 , n48491 );
and ( n48493 , n47296 , n47333 );
and ( n48494 , n47333 , n47359 );
and ( n48495 , n47296 , n47359 );
or ( n48496 , n48493 , n48494 , n48495 );
xor ( n48497 , n48492 , n48496 );
and ( n48498 , n47338 , n47342 );
and ( n48499 , n47342 , n47358 );
and ( n48500 , n47338 , n47358 );
or ( n48501 , n48498 , n48499 , n48500 );
and ( n48502 , n47320 , n47325 );
and ( n48503 , n47325 , n47331 );
and ( n48504 , n47320 , n47331 );
or ( n48505 , n48502 , n48503 , n48504 );
and ( n48506 , n47310 , n47311 );
and ( n48507 , n47311 , n47313 );
and ( n48508 , n47310 , n47313 );
or ( n48509 , n48506 , n48507 , n48508 );
and ( n48510 , n47321 , n47322 );
and ( n48511 , n47322 , n47324 );
and ( n48512 , n47321 , n47324 );
or ( n48513 , n48510 , n48511 , n48512 );
xor ( n48514 , n48509 , n48513 );
and ( n48515 , n7385 , n13256 );
and ( n48516 , n7808 , n12531 );
xor ( n48517 , n48515 , n48516 );
and ( n48518 , n8079 , n11718 );
xor ( n48519 , n48517 , n48518 );
xor ( n48520 , n48514 , n48519 );
xor ( n48521 , n48505 , n48520 );
and ( n48522 , n47327 , n47328 );
and ( n48523 , n47328 , n47330 );
and ( n48524 , n47327 , n47330 );
or ( n48525 , n48522 , n48523 , n48524 );
and ( n48526 , n6187 , n15691 );
and ( n48527 , n6569 , n14838 );
xor ( n48528 , n48526 , n48527 );
and ( n48529 , n6816 , n14044 );
xor ( n48530 , n48528 , n48529 );
xor ( n48531 , n48525 , n48530 );
and ( n48532 , n4959 , n18407 );
and ( n48533 , n5459 , n17422 );
xor ( n48534 , n48532 , n48533 );
and ( n48535 , n5819 , n16550 );
xor ( n48536 , n48534 , n48535 );
xor ( n48537 , n48531 , n48536 );
xor ( n48538 , n48521 , n48537 );
xor ( n48539 , n48501 , n48538 );
and ( n48540 , n47347 , n47351 );
and ( n48541 , n47351 , n47357 );
and ( n48542 , n47347 , n47357 );
or ( n48543 , n48540 , n48541 , n48542 );
and ( n48544 , n47376 , n47381 );
and ( n48545 , n47381 , n47387 );
and ( n48546 , n47376 , n47387 );
or ( n48547 , n48544 , n48545 , n48546 );
xor ( n48548 , n48543 , n48547 );
and ( n48549 , n47353 , n47354 );
and ( n48550 , n47354 , n47356 );
and ( n48551 , n47353 , n47356 );
or ( n48552 , n48549 , n48550 , n48551 );
and ( n48553 , n47377 , n47378 );
and ( n48554 , n47378 , n47380 );
and ( n48555 , n47377 , n47380 );
or ( n48556 , n48553 , n48554 , n48555 );
xor ( n48557 , n48552 , n48556 );
and ( n48558 , n4132 , n20976 );
and ( n48559 , n4438 , n20156 );
xor ( n48560 , n48558 , n48559 );
and ( n48561 , n4766 , n19222 );
xor ( n48562 , n48560 , n48561 );
xor ( n48563 , n48557 , n48562 );
xor ( n48564 , n48548 , n48563 );
xor ( n48565 , n48539 , n48564 );
xor ( n48566 , n48497 , n48565 );
xor ( n48567 , n48488 , n48566 );
and ( n48568 , n47372 , n47388 );
and ( n48569 , n47388 , n47404 );
and ( n48570 , n47372 , n47404 );
or ( n48571 , n48568 , n48569 , n48570 );
and ( n48572 , n47410 , n47421 );
xor ( n48573 , n48571 , n48572 );
and ( n48574 , n47393 , n47397 );
and ( n48575 , n47397 , n47403 );
and ( n48576 , n47393 , n47403 );
or ( n48577 , n48574 , n48575 , n48576 );
and ( n48578 , n47383 , n47384 );
and ( n48579 , n47384 , n47386 );
and ( n48580 , n47383 , n47386 );
or ( n48581 , n48578 , n48579 , n48580 );
and ( n48582 , n3182 , n24137 );
and ( n48583 , n3545 , n23075 );
xor ( n48584 , n48582 , n48583 );
and ( n48585 , n3801 , n22065 );
xor ( n48586 , n48584 , n48585 );
xor ( n48587 , n48581 , n48586 );
and ( n48588 , n2462 , n27296 );
and ( n48589 , n2779 , n26216 );
xor ( n48590 , n48588 , n48589 );
and ( n48591 , n3024 , n25163 );
xor ( n48592 , n48590 , n48591 );
xor ( n48593 , n48587 , n48592 );
xor ( n48594 , n48577 , n48593 );
and ( n48595 , n47399 , n47400 );
and ( n48596 , n47400 , n47402 );
and ( n48597 , n47399 , n47402 );
or ( n48598 , n48595 , n48596 , n48597 );
and ( n48599 , n47416 , n47417 );
and ( n48600 , n47417 , n47419 );
and ( n48601 , n47416 , n47419 );
or ( n48602 , n48599 , n48600 , n48601 );
xor ( n48603 , n48598 , n48602 );
and ( n48604 , n1933 , n30629 );
and ( n48605 , n2120 , n29508 );
xor ( n48606 , n48604 , n48605 );
and ( n48607 , n2324 , n28406 );
xor ( n48608 , n48606 , n48607 );
xor ( n48609 , n48603 , n48608 );
xor ( n48610 , n48594 , n48609 );
xor ( n48611 , n48573 , n48610 );
and ( n48612 , n47411 , n47414 );
and ( n48613 , n47414 , n47420 );
and ( n48614 , n47411 , n47420 );
or ( n48615 , n48612 , n48613 , n48614 );
not ( n48616 , n1383 );
and ( n48617 , n34193 , n1383 );
nor ( n48618 , n48616 , n48617 );
and ( n48619 , n1580 , n32999 );
xor ( n48620 , n48618 , n48619 );
and ( n48621 , n1694 , n31761 );
xor ( n48622 , n48620 , n48621 );
xor ( n48623 , n48615 , n48622 );
xor ( n48624 , n48611 , n48623 );
xor ( n48625 , n48567 , n48624 );
xor ( n48626 , n48487 , n48625 );
xor ( n48627 , n48362 , n48626 );
xor ( n48628 , n48280 , n48627 );
xor ( n48629 , n48271 , n48628 );
and ( n48630 , n47060 , n47063 );
and ( n48631 , n47063 , n47427 );
and ( n48632 , n47060 , n47427 );
or ( n48633 , n48630 , n48631 , n48632 );
xor ( n48634 , n48629 , n48633 );
and ( n48635 , n47428 , n47432 );
and ( n48636 , n47433 , n47436 );
or ( n48637 , n48635 , n48636 );
xor ( n48638 , n48634 , n48637 );
buf ( n48639 , n48638 );
buf ( n48640 , n48639 );
not ( n48641 , n48640 );
nor ( n48642 , n48641 , n8739 );
xor ( n48643 , n48263 , n48642 );
and ( n48644 , n47056 , n47441 );
and ( n48645 , n47442 , n47445 );
or ( n48646 , n48644 , n48645 );
xor ( n48647 , n48643 , n48646 );
buf ( n48648 , n48647 );
buf ( n48649 , n48648 );
not ( n48650 , n48649 );
buf ( n48651 , n574 );
not ( n48652 , n48651 );
nor ( n48653 , n48650 , n48652 );
xor ( n48654 , n47889 , n48653 );
xor ( n48655 , n47457 , n47886 );
nor ( n48656 , n47449 , n48652 );
and ( n48657 , n48655 , n48656 );
xor ( n48658 , n48655 , n48656 );
xor ( n48659 , n47461 , n47884 );
nor ( n48660 , n46248 , n48652 );
and ( n48661 , n48659 , n48660 );
xor ( n48662 , n48659 , n48660 );
xor ( n48663 , n47465 , n47882 );
nor ( n48664 , n45047 , n48652 );
and ( n48665 , n48663 , n48664 );
xor ( n48666 , n48663 , n48664 );
xor ( n48667 , n47469 , n47880 );
nor ( n48668 , n43843 , n48652 );
and ( n48669 , n48667 , n48668 );
xor ( n48670 , n48667 , n48668 );
xor ( n48671 , n47473 , n47878 );
nor ( n48672 , n42641 , n48652 );
and ( n48673 , n48671 , n48672 );
xor ( n48674 , n48671 , n48672 );
xor ( n48675 , n47477 , n47876 );
nor ( n48676 , n41437 , n48652 );
and ( n48677 , n48675 , n48676 );
xor ( n48678 , n48675 , n48676 );
xor ( n48679 , n47481 , n47874 );
nor ( n48680 , n40232 , n48652 );
and ( n48681 , n48679 , n48680 );
xor ( n48682 , n48679 , n48680 );
xor ( n48683 , n47485 , n47872 );
nor ( n48684 , n39027 , n48652 );
and ( n48685 , n48683 , n48684 );
xor ( n48686 , n48683 , n48684 );
xor ( n48687 , n47489 , n47870 );
nor ( n48688 , n37825 , n48652 );
and ( n48689 , n48687 , n48688 );
xor ( n48690 , n48687 , n48688 );
xor ( n48691 , n47493 , n47868 );
nor ( n48692 , n36620 , n48652 );
and ( n48693 , n48691 , n48692 );
xor ( n48694 , n48691 , n48692 );
xor ( n48695 , n47497 , n47866 );
nor ( n48696 , n35419 , n48652 );
and ( n48697 , n48695 , n48696 );
xor ( n48698 , n48695 , n48696 );
xor ( n48699 , n47501 , n47864 );
nor ( n48700 , n34224 , n48652 );
and ( n48701 , n48699 , n48700 );
xor ( n48702 , n48699 , n48700 );
xor ( n48703 , n47505 , n47862 );
nor ( n48704 , n33033 , n48652 );
and ( n48705 , n48703 , n48704 );
xor ( n48706 , n48703 , n48704 );
xor ( n48707 , n47509 , n47860 );
nor ( n48708 , n31867 , n48652 );
and ( n48709 , n48707 , n48708 );
xor ( n48710 , n48707 , n48708 );
xor ( n48711 , n47513 , n47858 );
nor ( n48712 , n30725 , n48652 );
and ( n48713 , n48711 , n48712 );
xor ( n48714 , n48711 , n48712 );
xor ( n48715 , n47517 , n47856 );
nor ( n48716 , n29596 , n48652 );
and ( n48717 , n48715 , n48716 );
xor ( n48718 , n48715 , n48716 );
xor ( n48719 , n47521 , n47854 );
nor ( n48720 , n28487 , n48652 );
and ( n48721 , n48719 , n48720 );
xor ( n48722 , n48719 , n48720 );
xor ( n48723 , n47525 , n47852 );
nor ( n48724 , n27397 , n48652 );
and ( n48725 , n48723 , n48724 );
xor ( n48726 , n48723 , n48724 );
xor ( n48727 , n47529 , n47850 );
nor ( n48728 , n26326 , n48652 );
and ( n48729 , n48727 , n48728 );
xor ( n48730 , n48727 , n48728 );
xor ( n48731 , n47533 , n47848 );
nor ( n48732 , n25272 , n48652 );
and ( n48733 , n48731 , n48732 );
xor ( n48734 , n48731 , n48732 );
xor ( n48735 , n47537 , n47846 );
nor ( n48736 , n24242 , n48652 );
and ( n48737 , n48735 , n48736 );
xor ( n48738 , n48735 , n48736 );
xor ( n48739 , n47541 , n47844 );
nor ( n48740 , n23225 , n48652 );
and ( n48741 , n48739 , n48740 );
xor ( n48742 , n48739 , n48740 );
xor ( n48743 , n47545 , n47842 );
nor ( n48744 , n22231 , n48652 );
and ( n48745 , n48743 , n48744 );
xor ( n48746 , n48743 , n48744 );
xor ( n48747 , n47549 , n47840 );
nor ( n48748 , n21258 , n48652 );
and ( n48749 , n48747 , n48748 );
xor ( n48750 , n48747 , n48748 );
xor ( n48751 , n47553 , n47838 );
nor ( n48752 , n20303 , n48652 );
and ( n48753 , n48751 , n48752 );
xor ( n48754 , n48751 , n48752 );
xor ( n48755 , n47557 , n47836 );
nor ( n48756 , n19365 , n48652 );
and ( n48757 , n48755 , n48756 );
xor ( n48758 , n48755 , n48756 );
xor ( n48759 , n47561 , n47834 );
nor ( n48760 , n18448 , n48652 );
and ( n48761 , n48759 , n48760 );
xor ( n48762 , n48759 , n48760 );
xor ( n48763 , n47565 , n47832 );
nor ( n48764 , n17548 , n48652 );
and ( n48765 , n48763 , n48764 );
xor ( n48766 , n48763 , n48764 );
xor ( n48767 , n47569 , n47830 );
nor ( n48768 , n16669 , n48652 );
and ( n48769 , n48767 , n48768 );
xor ( n48770 , n48767 , n48768 );
xor ( n48771 , n47573 , n47828 );
nor ( n48772 , n15809 , n48652 );
and ( n48773 , n48771 , n48772 );
xor ( n48774 , n48771 , n48772 );
xor ( n48775 , n47577 , n47826 );
nor ( n48776 , n14968 , n48652 );
and ( n48777 , n48775 , n48776 );
xor ( n48778 , n48775 , n48776 );
xor ( n48779 , n47581 , n47824 );
nor ( n48780 , n14147 , n48652 );
and ( n48781 , n48779 , n48780 );
xor ( n48782 , n48779 , n48780 );
xor ( n48783 , n47585 , n47822 );
nor ( n48784 , n13349 , n48652 );
and ( n48785 , n48783 , n48784 );
xor ( n48786 , n48783 , n48784 );
xor ( n48787 , n47589 , n47820 );
nor ( n48788 , n12564 , n48652 );
and ( n48789 , n48787 , n48788 );
xor ( n48790 , n48787 , n48788 );
xor ( n48791 , n47593 , n47818 );
nor ( n48792 , n11799 , n48652 );
and ( n48793 , n48791 , n48792 );
xor ( n48794 , n48791 , n48792 );
xor ( n48795 , n47597 , n47816 );
nor ( n48796 , n11050 , n48652 );
and ( n48797 , n48795 , n48796 );
xor ( n48798 , n48795 , n48796 );
xor ( n48799 , n47601 , n47814 );
nor ( n48800 , n10321 , n48652 );
and ( n48801 , n48799 , n48800 );
xor ( n48802 , n48799 , n48800 );
xor ( n48803 , n47605 , n47812 );
nor ( n48804 , n9429 , n48652 );
and ( n48805 , n48803 , n48804 );
xor ( n48806 , n48803 , n48804 );
xor ( n48807 , n47609 , n47810 );
nor ( n48808 , n8949 , n48652 );
and ( n48809 , n48807 , n48808 );
xor ( n48810 , n48807 , n48808 );
xor ( n48811 , n47613 , n47808 );
nor ( n48812 , n9437 , n48652 );
and ( n48813 , n48811 , n48812 );
xor ( n48814 , n48811 , n48812 );
xor ( n48815 , n47617 , n47806 );
nor ( n48816 , n9446 , n48652 );
and ( n48817 , n48815 , n48816 );
xor ( n48818 , n48815 , n48816 );
xor ( n48819 , n47621 , n47804 );
nor ( n48820 , n9455 , n48652 );
and ( n48821 , n48819 , n48820 );
xor ( n48822 , n48819 , n48820 );
xor ( n48823 , n47625 , n47802 );
nor ( n48824 , n9464 , n48652 );
and ( n48825 , n48823 , n48824 );
xor ( n48826 , n48823 , n48824 );
xor ( n48827 , n47629 , n47800 );
nor ( n48828 , n9473 , n48652 );
and ( n48829 , n48827 , n48828 );
xor ( n48830 , n48827 , n48828 );
xor ( n48831 , n47633 , n47798 );
nor ( n48832 , n9482 , n48652 );
and ( n48833 , n48831 , n48832 );
xor ( n48834 , n48831 , n48832 );
xor ( n48835 , n47637 , n47796 );
nor ( n48836 , n9491 , n48652 );
and ( n48837 , n48835 , n48836 );
xor ( n48838 , n48835 , n48836 );
xor ( n48839 , n47641 , n47794 );
nor ( n48840 , n9500 , n48652 );
and ( n48841 , n48839 , n48840 );
xor ( n48842 , n48839 , n48840 );
xor ( n48843 , n47645 , n47792 );
nor ( n48844 , n9509 , n48652 );
and ( n48845 , n48843 , n48844 );
xor ( n48846 , n48843 , n48844 );
xor ( n48847 , n47649 , n47790 );
nor ( n48848 , n9518 , n48652 );
and ( n48849 , n48847 , n48848 );
xor ( n48850 , n48847 , n48848 );
xor ( n48851 , n47653 , n47788 );
nor ( n48852 , n9527 , n48652 );
and ( n48853 , n48851 , n48852 );
xor ( n48854 , n48851 , n48852 );
xor ( n48855 , n47657 , n47786 );
nor ( n48856 , n9536 , n48652 );
and ( n48857 , n48855 , n48856 );
xor ( n48858 , n48855 , n48856 );
xor ( n48859 , n47661 , n47784 );
nor ( n48860 , n9545 , n48652 );
and ( n48861 , n48859 , n48860 );
xor ( n48862 , n48859 , n48860 );
xor ( n48863 , n47665 , n47782 );
nor ( n48864 , n9554 , n48652 );
and ( n48865 , n48863 , n48864 );
xor ( n48866 , n48863 , n48864 );
xor ( n48867 , n47669 , n47780 );
nor ( n48868 , n9563 , n48652 );
and ( n48869 , n48867 , n48868 );
xor ( n48870 , n48867 , n48868 );
xor ( n48871 , n47673 , n47778 );
nor ( n48872 , n9572 , n48652 );
and ( n48873 , n48871 , n48872 );
xor ( n48874 , n48871 , n48872 );
xor ( n48875 , n47677 , n47776 );
nor ( n48876 , n9581 , n48652 );
and ( n48877 , n48875 , n48876 );
xor ( n48878 , n48875 , n48876 );
xor ( n48879 , n47681 , n47774 );
nor ( n48880 , n9590 , n48652 );
and ( n48881 , n48879 , n48880 );
xor ( n48882 , n48879 , n48880 );
xor ( n48883 , n47685 , n47772 );
nor ( n48884 , n9599 , n48652 );
and ( n48885 , n48883 , n48884 );
xor ( n48886 , n48883 , n48884 );
xor ( n48887 , n47689 , n47770 );
nor ( n48888 , n9608 , n48652 );
and ( n48889 , n48887 , n48888 );
xor ( n48890 , n48887 , n48888 );
xor ( n48891 , n47693 , n47768 );
nor ( n48892 , n9617 , n48652 );
and ( n48893 , n48891 , n48892 );
xor ( n48894 , n48891 , n48892 );
xor ( n48895 , n47697 , n47766 );
nor ( n48896 , n9626 , n48652 );
and ( n48897 , n48895 , n48896 );
xor ( n48898 , n48895 , n48896 );
xor ( n48899 , n47701 , n47764 );
nor ( n48900 , n9635 , n48652 );
and ( n48901 , n48899 , n48900 );
xor ( n48902 , n48899 , n48900 );
xor ( n48903 , n47705 , n47762 );
nor ( n48904 , n9644 , n48652 );
and ( n48905 , n48903 , n48904 );
xor ( n48906 , n48903 , n48904 );
xor ( n48907 , n47709 , n47760 );
nor ( n48908 , n9653 , n48652 );
and ( n48909 , n48907 , n48908 );
xor ( n48910 , n48907 , n48908 );
xor ( n48911 , n47713 , n47758 );
nor ( n48912 , n9662 , n48652 );
and ( n48913 , n48911 , n48912 );
xor ( n48914 , n48911 , n48912 );
xor ( n48915 , n47717 , n47756 );
nor ( n48916 , n9671 , n48652 );
and ( n48917 , n48915 , n48916 );
xor ( n48918 , n48915 , n48916 );
xor ( n48919 , n47721 , n47754 );
nor ( n48920 , n9680 , n48652 );
and ( n48921 , n48919 , n48920 );
xor ( n48922 , n48919 , n48920 );
xor ( n48923 , n47725 , n47752 );
nor ( n48924 , n9689 , n48652 );
and ( n48925 , n48923 , n48924 );
xor ( n48926 , n48923 , n48924 );
xor ( n48927 , n47729 , n47750 );
nor ( n48928 , n9698 , n48652 );
and ( n48929 , n48927 , n48928 );
xor ( n48930 , n48927 , n48928 );
xor ( n48931 , n47733 , n47748 );
nor ( n48932 , n9707 , n48652 );
and ( n48933 , n48931 , n48932 );
xor ( n48934 , n48931 , n48932 );
xor ( n48935 , n47737 , n47746 );
nor ( n48936 , n9716 , n48652 );
and ( n48937 , n48935 , n48936 );
xor ( n48938 , n48935 , n48936 );
xor ( n48939 , n47741 , n47744 );
nor ( n48940 , n9725 , n48652 );
and ( n48941 , n48939 , n48940 );
xor ( n48942 , n48939 , n48940 );
xor ( n48943 , n47742 , n47743 );
nor ( n48944 , n9734 , n48652 );
and ( n48945 , n48943 , n48944 );
xor ( n48946 , n48943 , n48944 );
nor ( n48947 , n9752 , n47451 );
nor ( n48948 , n9743 , n48652 );
and ( n48949 , n48947 , n48948 );
and ( n48950 , n48946 , n48949 );
or ( n48951 , n48945 , n48950 );
and ( n48952 , n48942 , n48951 );
or ( n48953 , n48941 , n48952 );
and ( n48954 , n48938 , n48953 );
or ( n48955 , n48937 , n48954 );
and ( n48956 , n48934 , n48955 );
or ( n48957 , n48933 , n48956 );
and ( n48958 , n48930 , n48957 );
or ( n48959 , n48929 , n48958 );
and ( n48960 , n48926 , n48959 );
or ( n48961 , n48925 , n48960 );
and ( n48962 , n48922 , n48961 );
or ( n48963 , n48921 , n48962 );
and ( n48964 , n48918 , n48963 );
or ( n48965 , n48917 , n48964 );
and ( n48966 , n48914 , n48965 );
or ( n48967 , n48913 , n48966 );
and ( n48968 , n48910 , n48967 );
or ( n48969 , n48909 , n48968 );
and ( n48970 , n48906 , n48969 );
or ( n48971 , n48905 , n48970 );
and ( n48972 , n48902 , n48971 );
or ( n48973 , n48901 , n48972 );
and ( n48974 , n48898 , n48973 );
or ( n48975 , n48897 , n48974 );
and ( n48976 , n48894 , n48975 );
or ( n48977 , n48893 , n48976 );
and ( n48978 , n48890 , n48977 );
or ( n48979 , n48889 , n48978 );
and ( n48980 , n48886 , n48979 );
or ( n48981 , n48885 , n48980 );
and ( n48982 , n48882 , n48981 );
or ( n48983 , n48881 , n48982 );
and ( n48984 , n48878 , n48983 );
or ( n48985 , n48877 , n48984 );
and ( n48986 , n48874 , n48985 );
or ( n48987 , n48873 , n48986 );
and ( n48988 , n48870 , n48987 );
or ( n48989 , n48869 , n48988 );
and ( n48990 , n48866 , n48989 );
or ( n48991 , n48865 , n48990 );
and ( n48992 , n48862 , n48991 );
or ( n48993 , n48861 , n48992 );
and ( n48994 , n48858 , n48993 );
or ( n48995 , n48857 , n48994 );
and ( n48996 , n48854 , n48995 );
or ( n48997 , n48853 , n48996 );
and ( n48998 , n48850 , n48997 );
or ( n48999 , n48849 , n48998 );
and ( n49000 , n48846 , n48999 );
or ( n49001 , n48845 , n49000 );
and ( n49002 , n48842 , n49001 );
or ( n49003 , n48841 , n49002 );
and ( n49004 , n48838 , n49003 );
or ( n49005 , n48837 , n49004 );
and ( n49006 , n48834 , n49005 );
or ( n49007 , n48833 , n49006 );
and ( n49008 , n48830 , n49007 );
or ( n49009 , n48829 , n49008 );
and ( n49010 , n48826 , n49009 );
or ( n49011 , n48825 , n49010 );
and ( n49012 , n48822 , n49011 );
or ( n49013 , n48821 , n49012 );
and ( n49014 , n48818 , n49013 );
or ( n49015 , n48817 , n49014 );
and ( n49016 , n48814 , n49015 );
or ( n49017 , n48813 , n49016 );
and ( n49018 , n48810 , n49017 );
or ( n49019 , n48809 , n49018 );
and ( n49020 , n48806 , n49019 );
or ( n49021 , n48805 , n49020 );
and ( n49022 , n48802 , n49021 );
or ( n49023 , n48801 , n49022 );
and ( n49024 , n48798 , n49023 );
or ( n49025 , n48797 , n49024 );
and ( n49026 , n48794 , n49025 );
or ( n49027 , n48793 , n49026 );
and ( n49028 , n48790 , n49027 );
or ( n49029 , n48789 , n49028 );
and ( n49030 , n48786 , n49029 );
or ( n49031 , n48785 , n49030 );
and ( n49032 , n48782 , n49031 );
or ( n49033 , n48781 , n49032 );
and ( n49034 , n48778 , n49033 );
or ( n49035 , n48777 , n49034 );
and ( n49036 , n48774 , n49035 );
or ( n49037 , n48773 , n49036 );
and ( n49038 , n48770 , n49037 );
or ( n49039 , n48769 , n49038 );
and ( n49040 , n48766 , n49039 );
or ( n49041 , n48765 , n49040 );
and ( n49042 , n48762 , n49041 );
or ( n49043 , n48761 , n49042 );
and ( n49044 , n48758 , n49043 );
or ( n49045 , n48757 , n49044 );
and ( n49046 , n48754 , n49045 );
or ( n49047 , n48753 , n49046 );
and ( n49048 , n48750 , n49047 );
or ( n49049 , n48749 , n49048 );
and ( n49050 , n48746 , n49049 );
or ( n49051 , n48745 , n49050 );
and ( n49052 , n48742 , n49051 );
or ( n49053 , n48741 , n49052 );
and ( n49054 , n48738 , n49053 );
or ( n49055 , n48737 , n49054 );
and ( n49056 , n48734 , n49055 );
or ( n49057 , n48733 , n49056 );
and ( n49058 , n48730 , n49057 );
or ( n49059 , n48729 , n49058 );
and ( n49060 , n48726 , n49059 );
or ( n49061 , n48725 , n49060 );
and ( n49062 , n48722 , n49061 );
or ( n49063 , n48721 , n49062 );
and ( n49064 , n48718 , n49063 );
or ( n49065 , n48717 , n49064 );
and ( n49066 , n48714 , n49065 );
or ( n49067 , n48713 , n49066 );
and ( n49068 , n48710 , n49067 );
or ( n49069 , n48709 , n49068 );
and ( n49070 , n48706 , n49069 );
or ( n49071 , n48705 , n49070 );
and ( n49072 , n48702 , n49071 );
or ( n49073 , n48701 , n49072 );
and ( n49074 , n48698 , n49073 );
or ( n49075 , n48697 , n49074 );
and ( n49076 , n48694 , n49075 );
or ( n49077 , n48693 , n49076 );
and ( n49078 , n48690 , n49077 );
or ( n49079 , n48689 , n49078 );
and ( n49080 , n48686 , n49079 );
or ( n49081 , n48685 , n49080 );
and ( n49082 , n48682 , n49081 );
or ( n49083 , n48681 , n49082 );
and ( n49084 , n48678 , n49083 );
or ( n49085 , n48677 , n49084 );
and ( n49086 , n48674 , n49085 );
or ( n49087 , n48673 , n49086 );
and ( n49088 , n48670 , n49087 );
or ( n49089 , n48669 , n49088 );
and ( n49090 , n48666 , n49089 );
or ( n49091 , n48665 , n49090 );
and ( n49092 , n48662 , n49091 );
or ( n49093 , n48661 , n49092 );
and ( n49094 , n48658 , n49093 );
or ( n49095 , n48657 , n49094 );
xor ( n49096 , n48654 , n49095 );
and ( n49097 , n33403 , n1597 );
nor ( n49098 , n1598 , n49097 );
nor ( n49099 , n1766 , n32231 );
xor ( n49100 , n49098 , n49099 );
and ( n49101 , n47891 , n47892 );
and ( n49102 , n47893 , n47896 );
or ( n49103 , n49101 , n49102 );
xor ( n49104 , n49100 , n49103 );
nor ( n49105 , n1945 , n31083 );
xor ( n49106 , n49104 , n49105 );
and ( n49107 , n47897 , n47898 );
and ( n49108 , n47899 , n47902 );
or ( n49109 , n49107 , n49108 );
xor ( n49110 , n49106 , n49109 );
nor ( n49111 , n2137 , n29948 );
xor ( n49112 , n49110 , n49111 );
and ( n49113 , n47903 , n47904 );
and ( n49114 , n47905 , n47908 );
or ( n49115 , n49113 , n49114 );
xor ( n49116 , n49112 , n49115 );
nor ( n49117 , n2343 , n28833 );
xor ( n49118 , n49116 , n49117 );
and ( n49119 , n47909 , n47910 );
and ( n49120 , n47911 , n47914 );
or ( n49121 , n49119 , n49120 );
xor ( n49122 , n49118 , n49121 );
nor ( n49123 , n2566 , n27737 );
xor ( n49124 , n49122 , n49123 );
and ( n49125 , n47915 , n47916 );
and ( n49126 , n47917 , n47920 );
or ( n49127 , n49125 , n49126 );
xor ( n49128 , n49124 , n49127 );
nor ( n49129 , n2797 , n26660 );
xor ( n49130 , n49128 , n49129 );
and ( n49131 , n47921 , n47922 );
and ( n49132 , n47923 , n47926 );
or ( n49133 , n49131 , n49132 );
xor ( n49134 , n49130 , n49133 );
nor ( n49135 , n3043 , n25600 );
xor ( n49136 , n49134 , n49135 );
and ( n49137 , n47927 , n47928 );
and ( n49138 , n47929 , n47932 );
or ( n49139 , n49137 , n49138 );
xor ( n49140 , n49136 , n49139 );
nor ( n49141 , n3300 , n24564 );
xor ( n49142 , n49140 , n49141 );
and ( n49143 , n47933 , n47934 );
and ( n49144 , n47935 , n47938 );
or ( n49145 , n49143 , n49144 );
xor ( n49146 , n49142 , n49145 );
nor ( n49147 , n3570 , n23541 );
xor ( n49148 , n49146 , n49147 );
and ( n49149 , n47939 , n47940 );
and ( n49150 , n47941 , n47944 );
or ( n49151 , n49149 , n49150 );
xor ( n49152 , n49148 , n49151 );
nor ( n49153 , n3853 , n22541 );
xor ( n49154 , n49152 , n49153 );
and ( n49155 , n47945 , n47946 );
and ( n49156 , n47947 , n47950 );
or ( n49157 , n49155 , n49156 );
xor ( n49158 , n49154 , n49157 );
nor ( n49159 , n4151 , n21562 );
xor ( n49160 , n49158 , n49159 );
and ( n49161 , n47951 , n47952 );
and ( n49162 , n47953 , n47956 );
or ( n49163 , n49161 , n49162 );
xor ( n49164 , n49160 , n49163 );
nor ( n49165 , n4458 , n20601 );
xor ( n49166 , n49164 , n49165 );
and ( n49167 , n47957 , n47958 );
and ( n49168 , n47959 , n47962 );
or ( n49169 , n49167 , n49168 );
xor ( n49170 , n49166 , n49169 );
nor ( n49171 , n4786 , n19657 );
xor ( n49172 , n49170 , n49171 );
and ( n49173 , n47963 , n47964 );
and ( n49174 , n47965 , n47968 );
or ( n49175 , n49173 , n49174 );
xor ( n49176 , n49172 , n49175 );
nor ( n49177 , n5126 , n18734 );
xor ( n49178 , n49176 , n49177 );
and ( n49179 , n47969 , n47970 );
and ( n49180 , n47971 , n47974 );
or ( n49181 , n49179 , n49180 );
xor ( n49182 , n49178 , n49181 );
nor ( n49183 , n5477 , n17828 );
xor ( n49184 , n49182 , n49183 );
and ( n49185 , n47975 , n47976 );
and ( n49186 , n47977 , n47980 );
or ( n49187 , n49185 , n49186 );
xor ( n49188 , n49184 , n49187 );
nor ( n49189 , n5838 , n16943 );
xor ( n49190 , n49188 , n49189 );
and ( n49191 , n47981 , n47982 );
and ( n49192 , n47983 , n47986 );
or ( n49193 , n49191 , n49192 );
xor ( n49194 , n49190 , n49193 );
nor ( n49195 , n6212 , n16077 );
xor ( n49196 , n49194 , n49195 );
and ( n49197 , n47987 , n47988 );
and ( n49198 , n47989 , n47992 );
or ( n49199 , n49197 , n49198 );
xor ( n49200 , n49196 , n49199 );
nor ( n49201 , n6596 , n15230 );
xor ( n49202 , n49200 , n49201 );
and ( n49203 , n47993 , n47994 );
and ( n49204 , n47995 , n47998 );
or ( n49205 , n49203 , n49204 );
xor ( n49206 , n49202 , n49205 );
nor ( n49207 , n6997 , n14403 );
xor ( n49208 , n49206 , n49207 );
and ( n49209 , n47999 , n48000 );
and ( n49210 , n48001 , n48004 );
or ( n49211 , n49209 , n49210 );
xor ( n49212 , n49208 , n49211 );
nor ( n49213 , n7413 , n13599 );
xor ( n49214 , n49212 , n49213 );
and ( n49215 , n48005 , n48006 );
and ( n49216 , n48007 , n48010 );
or ( n49217 , n49215 , n49216 );
xor ( n49218 , n49214 , n49217 );
nor ( n49219 , n7841 , n12808 );
xor ( n49220 , n49218 , n49219 );
and ( n49221 , n48011 , n48012 );
and ( n49222 , n48013 , n48016 );
or ( n49223 , n49221 , n49222 );
xor ( n49224 , n49220 , n49223 );
nor ( n49225 , n8281 , n12037 );
xor ( n49226 , n49224 , n49225 );
and ( n49227 , n48017 , n48018 );
and ( n49228 , n48019 , n48022 );
or ( n49229 , n49227 , n49228 );
xor ( n49230 , n49226 , n49229 );
nor ( n49231 , n8737 , n11282 );
xor ( n49232 , n49230 , n49231 );
and ( n49233 , n48023 , n48024 );
and ( n49234 , n48025 , n48028 );
or ( n49235 , n49233 , n49234 );
xor ( n49236 , n49232 , n49235 );
nor ( n49237 , n9420 , n10547 );
xor ( n49238 , n49236 , n49237 );
and ( n49239 , n48029 , n48030 );
and ( n49240 , n48031 , n48034 );
or ( n49241 , n49239 , n49240 );
xor ( n49242 , n49238 , n49241 );
nor ( n49243 , n10312 , n9829 );
xor ( n49244 , n49242 , n49243 );
and ( n49245 , n48035 , n48036 );
and ( n49246 , n48037 , n48040 );
or ( n49247 , n49245 , n49246 );
xor ( n49248 , n49244 , n49247 );
nor ( n49249 , n11041 , n8955 );
xor ( n49250 , n49248 , n49249 );
and ( n49251 , n48041 , n48042 );
and ( n49252 , n48043 , n48046 );
or ( n49253 , n49251 , n49252 );
xor ( n49254 , n49250 , n49253 );
nor ( n49255 , n11790 , n603 );
xor ( n49256 , n49254 , n49255 );
and ( n49257 , n48047 , n48048 );
and ( n49258 , n48049 , n48052 );
or ( n49259 , n49257 , n49258 );
xor ( n49260 , n49256 , n49259 );
nor ( n49261 , n12555 , n652 );
xor ( n49262 , n49260 , n49261 );
and ( n49263 , n48053 , n48054 );
and ( n49264 , n48055 , n48058 );
or ( n49265 , n49263 , n49264 );
xor ( n49266 , n49262 , n49265 );
nor ( n49267 , n13340 , n624 );
xor ( n49268 , n49266 , n49267 );
and ( n49269 , n48059 , n48060 );
and ( n49270 , n48061 , n48064 );
or ( n49271 , n49269 , n49270 );
xor ( n49272 , n49268 , n49271 );
nor ( n49273 , n14138 , n648 );
xor ( n49274 , n49272 , n49273 );
and ( n49275 , n48065 , n48066 );
and ( n49276 , n48067 , n48070 );
or ( n49277 , n49275 , n49276 );
xor ( n49278 , n49274 , n49277 );
nor ( n49279 , n14959 , n686 );
xor ( n49280 , n49278 , n49279 );
and ( n49281 , n48071 , n48072 );
and ( n49282 , n48073 , n48076 );
or ( n49283 , n49281 , n49282 );
xor ( n49284 , n49280 , n49283 );
nor ( n49285 , n15800 , n735 );
xor ( n49286 , n49284 , n49285 );
and ( n49287 , n48077 , n48078 );
and ( n49288 , n48079 , n48082 );
or ( n49289 , n49287 , n49288 );
xor ( n49290 , n49286 , n49289 );
nor ( n49291 , n16660 , n798 );
xor ( n49292 , n49290 , n49291 );
and ( n49293 , n48083 , n48084 );
and ( n49294 , n48085 , n48088 );
or ( n49295 , n49293 , n49294 );
xor ( n49296 , n49292 , n49295 );
nor ( n49297 , n17539 , n870 );
xor ( n49298 , n49296 , n49297 );
and ( n49299 , n48089 , n48090 );
and ( n49300 , n48091 , n48094 );
or ( n49301 , n49299 , n49300 );
xor ( n49302 , n49298 , n49301 );
nor ( n49303 , n18439 , n960 );
xor ( n49304 , n49302 , n49303 );
and ( n49305 , n48095 , n48096 );
and ( n49306 , n48097 , n48100 );
or ( n49307 , n49305 , n49306 );
xor ( n49308 , n49304 , n49307 );
nor ( n49309 , n19356 , n1064 );
xor ( n49310 , n49308 , n49309 );
and ( n49311 , n48101 , n48102 );
and ( n49312 , n48103 , n48106 );
or ( n49313 , n49311 , n49312 );
xor ( n49314 , n49310 , n49313 );
nor ( n49315 , n20294 , n1178 );
xor ( n49316 , n49314 , n49315 );
and ( n49317 , n48107 , n48108 );
and ( n49318 , n48109 , n48112 );
or ( n49319 , n49317 , n49318 );
xor ( n49320 , n49316 , n49319 );
nor ( n49321 , n21249 , n1305 );
xor ( n49322 , n49320 , n49321 );
and ( n49323 , n48113 , n48114 );
and ( n49324 , n48115 , n48118 );
or ( n49325 , n49323 , n49324 );
xor ( n49326 , n49322 , n49325 );
nor ( n49327 , n22222 , n1447 );
xor ( n49328 , n49326 , n49327 );
and ( n49329 , n48119 , n48120 );
and ( n49330 , n48121 , n48124 );
or ( n49331 , n49329 , n49330 );
xor ( n49332 , n49328 , n49331 );
nor ( n49333 , n23216 , n1600 );
xor ( n49334 , n49332 , n49333 );
and ( n49335 , n48125 , n48126 );
and ( n49336 , n48127 , n48130 );
or ( n49337 , n49335 , n49336 );
xor ( n49338 , n49334 , n49337 );
nor ( n49339 , n24233 , n1768 );
xor ( n49340 , n49338 , n49339 );
and ( n49341 , n48131 , n48132 );
and ( n49342 , n48133 , n48136 );
or ( n49343 , n49341 , n49342 );
xor ( n49344 , n49340 , n49343 );
nor ( n49345 , n25263 , n1947 );
xor ( n49346 , n49344 , n49345 );
and ( n49347 , n48137 , n48138 );
and ( n49348 , n48139 , n48142 );
or ( n49349 , n49347 , n49348 );
xor ( n49350 , n49346 , n49349 );
nor ( n49351 , n26317 , n2139 );
xor ( n49352 , n49350 , n49351 );
and ( n49353 , n48143 , n48144 );
and ( n49354 , n48145 , n48148 );
or ( n49355 , n49353 , n49354 );
xor ( n49356 , n49352 , n49355 );
nor ( n49357 , n27388 , n2345 );
xor ( n49358 , n49356 , n49357 );
and ( n49359 , n48149 , n48150 );
and ( n49360 , n48151 , n48154 );
or ( n49361 , n49359 , n49360 );
xor ( n49362 , n49358 , n49361 );
nor ( n49363 , n28478 , n2568 );
xor ( n49364 , n49362 , n49363 );
and ( n49365 , n48155 , n48156 );
and ( n49366 , n48157 , n48160 );
or ( n49367 , n49365 , n49366 );
xor ( n49368 , n49364 , n49367 );
nor ( n49369 , n29587 , n2799 );
xor ( n49370 , n49368 , n49369 );
and ( n49371 , n48161 , n48162 );
and ( n49372 , n48163 , n48166 );
or ( n49373 , n49371 , n49372 );
xor ( n49374 , n49370 , n49373 );
nor ( n49375 , n30716 , n3045 );
xor ( n49376 , n49374 , n49375 );
and ( n49377 , n48167 , n48168 );
and ( n49378 , n48169 , n48172 );
or ( n49379 , n49377 , n49378 );
xor ( n49380 , n49376 , n49379 );
nor ( n49381 , n31858 , n3302 );
xor ( n49382 , n49380 , n49381 );
and ( n49383 , n48173 , n48174 );
and ( n49384 , n48175 , n48178 );
or ( n49385 , n49383 , n49384 );
xor ( n49386 , n49382 , n49385 );
nor ( n49387 , n33024 , n3572 );
xor ( n49388 , n49386 , n49387 );
and ( n49389 , n48179 , n48180 );
and ( n49390 , n48181 , n48184 );
or ( n49391 , n49389 , n49390 );
xor ( n49392 , n49388 , n49391 );
nor ( n49393 , n34215 , n3855 );
xor ( n49394 , n49392 , n49393 );
and ( n49395 , n48185 , n48186 );
and ( n49396 , n48187 , n48190 );
or ( n49397 , n49395 , n49396 );
xor ( n49398 , n49394 , n49397 );
nor ( n49399 , n35410 , n4153 );
xor ( n49400 , n49398 , n49399 );
and ( n49401 , n48191 , n48192 );
and ( n49402 , n48193 , n48196 );
or ( n49403 , n49401 , n49402 );
xor ( n49404 , n49400 , n49403 );
nor ( n49405 , n36611 , n4460 );
xor ( n49406 , n49404 , n49405 );
and ( n49407 , n48197 , n48198 );
and ( n49408 , n48199 , n48202 );
or ( n49409 , n49407 , n49408 );
xor ( n49410 , n49406 , n49409 );
nor ( n49411 , n37816 , n4788 );
xor ( n49412 , n49410 , n49411 );
and ( n49413 , n48203 , n48204 );
and ( n49414 , n48205 , n48208 );
or ( n49415 , n49413 , n49414 );
xor ( n49416 , n49412 , n49415 );
nor ( n49417 , n39018 , n5128 );
xor ( n49418 , n49416 , n49417 );
and ( n49419 , n48209 , n48210 );
and ( n49420 , n48211 , n48214 );
or ( n49421 , n49419 , n49420 );
xor ( n49422 , n49418 , n49421 );
nor ( n49423 , n40223 , n5479 );
xor ( n49424 , n49422 , n49423 );
and ( n49425 , n48215 , n48216 );
and ( n49426 , n48217 , n48220 );
or ( n49427 , n49425 , n49426 );
xor ( n49428 , n49424 , n49427 );
nor ( n49429 , n41428 , n5840 );
xor ( n49430 , n49428 , n49429 );
and ( n49431 , n48221 , n48222 );
and ( n49432 , n48223 , n48226 );
or ( n49433 , n49431 , n49432 );
xor ( n49434 , n49430 , n49433 );
nor ( n49435 , n42632 , n6214 );
xor ( n49436 , n49434 , n49435 );
and ( n49437 , n48227 , n48228 );
and ( n49438 , n48229 , n48232 );
or ( n49439 , n49437 , n49438 );
xor ( n49440 , n49436 , n49439 );
nor ( n49441 , n43834 , n6598 );
xor ( n49442 , n49440 , n49441 );
and ( n49443 , n48233 , n48234 );
and ( n49444 , n48235 , n48238 );
or ( n49445 , n49443 , n49444 );
xor ( n49446 , n49442 , n49445 );
nor ( n49447 , n45038 , n6999 );
xor ( n49448 , n49446 , n49447 );
and ( n49449 , n48239 , n48240 );
and ( n49450 , n48241 , n48244 );
or ( n49451 , n49449 , n49450 );
xor ( n49452 , n49448 , n49451 );
nor ( n49453 , n46239 , n7415 );
xor ( n49454 , n49452 , n49453 );
and ( n49455 , n48245 , n48246 );
and ( n49456 , n48247 , n48250 );
or ( n49457 , n49455 , n49456 );
xor ( n49458 , n49454 , n49457 );
nor ( n49459 , n47440 , n7843 );
xor ( n49460 , n49458 , n49459 );
and ( n49461 , n48251 , n48252 );
and ( n49462 , n48253 , n48256 );
or ( n49463 , n49461 , n49462 );
xor ( n49464 , n49460 , n49463 );
nor ( n49465 , n48641 , n8283 );
xor ( n49466 , n49464 , n49465 );
and ( n49467 , n48257 , n48258 );
and ( n49468 , n48259 , n48262 );
or ( n49469 , n49467 , n49468 );
xor ( n49470 , n49466 , n49469 );
and ( n49471 , n48275 , n48279 );
and ( n49472 , n48279 , n48627 );
and ( n49473 , n48275 , n48627 );
or ( n49474 , n49471 , n49472 , n49473 );
and ( n49475 , n33774 , n1551 );
not ( n49476 , n1551 );
nor ( n49477 , n49475 , n49476 );
xor ( n49478 , n49474 , n49477 );
and ( n49479 , n48288 , n48292 );
and ( n49480 , n48292 , n48360 );
and ( n49481 , n48288 , n48360 );
or ( n49482 , n49479 , n49480 , n49481 );
and ( n49483 , n48284 , n48361 );
and ( n49484 , n48361 , n48626 );
and ( n49485 , n48284 , n48626 );
or ( n49486 , n49483 , n49484 , n49485 );
xor ( n49487 , n49482 , n49486 );
and ( n49488 , n48366 , n48486 );
and ( n49489 , n48486 , n48625 );
and ( n49490 , n48366 , n48625 );
or ( n49491 , n49488 , n49489 , n49490 );
and ( n49492 , n48297 , n48301 );
and ( n49493 , n48301 , n48359 );
and ( n49494 , n48297 , n48359 );
or ( n49495 , n49492 , n49493 , n49494 );
and ( n49496 , n48370 , n48374 );
and ( n49497 , n48374 , n48485 );
and ( n49498 , n48370 , n48485 );
or ( n49499 , n49496 , n49497 , n49498 );
xor ( n49500 , n49495 , n49499 );
and ( n49501 , n48328 , n48332 );
and ( n49502 , n48332 , n48338 );
and ( n49503 , n48328 , n48338 );
or ( n49504 , n49501 , n49502 , n49503 );
and ( n49505 , n48306 , n48310 );
and ( n49506 , n48310 , n48358 );
and ( n49507 , n48306 , n48358 );
or ( n49508 , n49505 , n49506 , n49507 );
xor ( n49509 , n49504 , n49508 );
and ( n49510 , n48315 , n48319 );
and ( n49511 , n48319 , n48357 );
and ( n49512 , n48315 , n48357 );
or ( n49513 , n49510 , n49511 , n49512 );
and ( n49514 , n48383 , n48408 );
and ( n49515 , n48408 , n48446 );
and ( n49516 , n48383 , n48446 );
or ( n49517 , n49514 , n49515 , n49516 );
xor ( n49518 , n49513 , n49517 );
and ( n49519 , n48324 , n48339 );
and ( n49520 , n48339 , n48356 );
and ( n49521 , n48324 , n48356 );
or ( n49522 , n49519 , n49520 , n49521 );
and ( n49523 , n48387 , n48391 );
and ( n49524 , n48391 , n48407 );
and ( n49525 , n48387 , n48407 );
or ( n49526 , n49523 , n49524 , n49525 );
xor ( n49527 , n49522 , n49526 );
and ( n49528 , n48344 , n48349 );
and ( n49529 , n48349 , n48355 );
and ( n49530 , n48344 , n48355 );
or ( n49531 , n49528 , n49529 , n49530 );
and ( n49532 , n48334 , n48335 );
and ( n49533 , n48335 , n48337 );
and ( n49534 , n48334 , n48337 );
or ( n49535 , n49532 , n49533 , n49534 );
and ( n49536 , n48345 , n48346 );
and ( n49537 , n48346 , n48348 );
and ( n49538 , n48345 , n48348 );
or ( n49539 , n49536 , n49537 , n49538 );
xor ( n49540 , n49535 , n49539 );
and ( n49541 , n30695 , n2100 );
and ( n49542 , n31836 , n1882 );
xor ( n49543 , n49541 , n49542 );
and ( n49544 , n32649 , n1738 );
xor ( n49545 , n49543 , n49544 );
xor ( n49546 , n49540 , n49545 );
xor ( n49547 , n49531 , n49546 );
and ( n49548 , n48351 , n48352 );
and ( n49549 , n48352 , n48354 );
and ( n49550 , n48351 , n48354 );
or ( n49551 , n49548 , n49549 , n49550 );
and ( n49552 , n27361 , n2739 );
and ( n49553 , n28456 , n2544 );
xor ( n49554 , n49552 , n49553 );
and ( n49555 , n29559 , n2298 );
xor ( n49556 , n49554 , n49555 );
xor ( n49557 , n49551 , n49556 );
and ( n49558 , n24214 , n3495 );
and ( n49559 , n25243 , n3271 );
xor ( n49560 , n49558 , n49559 );
and ( n49561 , n26296 , n2981 );
xor ( n49562 , n49560 , n49561 );
xor ( n49563 , n49557 , n49562 );
xor ( n49564 , n49547 , n49563 );
xor ( n49565 , n49527 , n49564 );
xor ( n49566 , n49518 , n49565 );
xor ( n49567 , n49509 , n49566 );
xor ( n49568 , n49500 , n49567 );
xor ( n49569 , n49491 , n49568 );
and ( n49570 , n48488 , n48566 );
and ( n49571 , n48566 , n48624 );
and ( n49572 , n48488 , n48624 );
or ( n49573 , n49570 , n49571 , n49572 );
and ( n49574 , n48379 , n48447 );
and ( n49575 , n48447 , n48484 );
and ( n49576 , n48379 , n48484 );
or ( n49577 , n49574 , n49575 , n49576 );
and ( n49578 , n48492 , n48496 );
and ( n49579 , n48496 , n48565 );
and ( n49580 , n48492 , n48565 );
or ( n49581 , n49578 , n49579 , n49580 );
xor ( n49582 , n49577 , n49581 );
and ( n49583 , n48452 , n48456 );
and ( n49584 , n48456 , n48483 );
and ( n49585 , n48452 , n48483 );
or ( n49586 , n49583 , n49584 , n49585 );
and ( n49587 , n48413 , n48429 );
and ( n49588 , n48429 , n48445 );
and ( n49589 , n48413 , n48445 );
or ( n49590 , n49587 , n49588 , n49589 );
and ( n49591 , n48396 , n48400 );
and ( n49592 , n48400 , n48406 );
and ( n49593 , n48396 , n48406 );
or ( n49594 , n49591 , n49592 , n49593 );
and ( n49595 , n48417 , n48422 );
and ( n49596 , n48422 , n48428 );
and ( n49597 , n48417 , n48428 );
or ( n49598 , n49595 , n49596 , n49597 );
xor ( n49599 , n49594 , n49598 );
and ( n49600 , n48402 , n48403 );
and ( n49601 , n48403 , n48405 );
and ( n49602 , n48402 , n48405 );
or ( n49603 , n49600 , n49601 , n49602 );
and ( n49604 , n48418 , n48419 );
and ( n49605 , n48419 , n48421 );
and ( n49606 , n48418 , n48421 );
or ( n49607 , n49604 , n49605 , n49606 );
xor ( n49608 , n49603 , n49607 );
and ( n49609 , n21216 , n4403 );
and ( n49610 , n22186 , n4102 );
xor ( n49611 , n49609 , n49610 );
and ( n49612 , n22892 , n3749 );
xor ( n49613 , n49611 , n49612 );
xor ( n49614 , n49608 , n49613 );
xor ( n49615 , n49599 , n49614 );
xor ( n49616 , n49590 , n49615 );
and ( n49617 , n48434 , n48438 );
and ( n49618 , n48438 , n48444 );
and ( n49619 , n48434 , n48444 );
or ( n49620 , n49617 , n49618 , n49619 );
and ( n49621 , n48424 , n48425 );
and ( n49622 , n48425 , n48427 );
and ( n49623 , n48424 , n48427 );
or ( n49624 , n49621 , n49622 , n49623 );
and ( n49625 , n18144 , n5408 );
and ( n49626 , n19324 , n5103 );
xor ( n49627 , n49625 , n49626 );
and ( n49628 , n20233 , n4730 );
xor ( n49629 , n49627 , n49628 );
xor ( n49630 , n49624 , n49629 );
and ( n49631 , n15758 , n6504 );
and ( n49632 , n16637 , n6132 );
xor ( n49633 , n49631 , n49632 );
and ( n49634 , n17512 , n5765 );
xor ( n49635 , n49633 , n49634 );
xor ( n49636 , n49630 , n49635 );
xor ( n49637 , n49620 , n49636 );
and ( n49638 , n48440 , n48441 );
and ( n49639 , n48441 , n48443 );
and ( n49640 , n48440 , n48443 );
or ( n49641 , n49638 , n49639 , n49640 );
and ( n49642 , n48471 , n48472 );
and ( n49643 , n48472 , n48474 );
and ( n49644 , n48471 , n48474 );
or ( n49645 , n49642 , n49643 , n49644 );
xor ( n49646 , n49641 , n49645 );
and ( n49647 , n13322 , n7662 );
and ( n49648 , n14118 , n7310 );
xor ( n49649 , n49647 , n49648 );
and ( n49650 , n14938 , n6971 );
xor ( n49651 , n49649 , n49650 );
xor ( n49652 , n49646 , n49651 );
xor ( n49653 , n49637 , n49652 );
xor ( n49654 , n49616 , n49653 );
xor ( n49655 , n49586 , n49654 );
and ( n49656 , n48461 , n48465 );
and ( n49657 , n48465 , n48482 );
and ( n49658 , n48461 , n48482 );
or ( n49659 , n49656 , n49657 , n49658 );
and ( n49660 , n48505 , n48520 );
and ( n49661 , n48520 , n48537 );
and ( n49662 , n48505 , n48537 );
or ( n49663 , n49660 , n49661 , n49662 );
xor ( n49664 , n49659 , n49663 );
and ( n49665 , n48470 , n48475 );
and ( n49666 , n48475 , n48481 );
and ( n49667 , n48470 , n48481 );
or ( n49668 , n49665 , n49666 , n49667 );
and ( n49669 , n48509 , n48513 );
and ( n49670 , n48513 , n48519 );
and ( n49671 , n48509 , n48519 );
or ( n49672 , n49669 , n49670 , n49671 );
xor ( n49673 , n49668 , n49672 );
and ( n49674 , n48477 , n48478 );
and ( n49675 , n48478 , n48480 );
and ( n49676 , n48477 , n48480 );
or ( n49677 , n49674 , n49675 , n49676 );
and ( n49678 , n11015 , n9348 );
and ( n49679 , n11769 , n8669 );
xor ( n49680 , n49678 , n49679 );
and ( n49681 , n12320 , n8243 );
xor ( n49682 , n49680 , n49681 );
xor ( n49683 , n49677 , n49682 );
and ( n49684 , n8718 , n11718 );
and ( n49685 , n9400 , n10977 );
xor ( n49686 , n49684 , n49685 );
buf ( n49687 , n10291 );
xor ( n49688 , n49686 , n49687 );
xor ( n49689 , n49683 , n49688 );
xor ( n49690 , n49673 , n49689 );
xor ( n49691 , n49664 , n49690 );
xor ( n49692 , n49655 , n49691 );
xor ( n49693 , n49582 , n49692 );
xor ( n49694 , n49573 , n49693 );
and ( n49695 , n48611 , n48623 );
and ( n49696 , n48571 , n48572 );
and ( n49697 , n48572 , n48610 );
and ( n49698 , n48571 , n48610 );
or ( n49699 , n49696 , n49697 , n49698 );
and ( n49700 , n48501 , n48538 );
and ( n49701 , n48538 , n48564 );
and ( n49702 , n48501 , n48564 );
or ( n49703 , n49700 , n49701 , n49702 );
xor ( n49704 , n49699 , n49703 );
and ( n49705 , n48543 , n48547 );
and ( n49706 , n48547 , n48563 );
and ( n49707 , n48543 , n48563 );
or ( n49708 , n49705 , n49706 , n49707 );
and ( n49709 , n48525 , n48530 );
and ( n49710 , n48530 , n48536 );
and ( n49711 , n48525 , n48536 );
or ( n49712 , n49709 , n49710 , n49711 );
and ( n49713 , n48515 , n48516 );
and ( n49714 , n48516 , n48518 );
and ( n49715 , n48515 , n48518 );
or ( n49716 , n49713 , n49714 , n49715 );
and ( n49717 , n48526 , n48527 );
and ( n49718 , n48527 , n48529 );
and ( n49719 , n48526 , n48529 );
or ( n49720 , n49717 , n49718 , n49719 );
xor ( n49721 , n49716 , n49720 );
and ( n49722 , n7385 , n14044 );
and ( n49723 , n7808 , n13256 );
xor ( n49724 , n49722 , n49723 );
and ( n49725 , n8079 , n12531 );
xor ( n49726 , n49724 , n49725 );
xor ( n49727 , n49721 , n49726 );
xor ( n49728 , n49712 , n49727 );
and ( n49729 , n48532 , n48533 );
and ( n49730 , n48533 , n48535 );
and ( n49731 , n48532 , n48535 );
or ( n49732 , n49729 , n49730 , n49731 );
and ( n49733 , n6187 , n16550 );
and ( n49734 , n6569 , n15691 );
xor ( n49735 , n49733 , n49734 );
and ( n49736 , n6816 , n14838 );
xor ( n49737 , n49735 , n49736 );
xor ( n49738 , n49732 , n49737 );
and ( n49739 , n4959 , n19222 );
and ( n49740 , n5459 , n18407 );
xor ( n49741 , n49739 , n49740 );
and ( n49742 , n5819 , n17422 );
xor ( n49743 , n49741 , n49742 );
xor ( n49744 , n49738 , n49743 );
xor ( n49745 , n49728 , n49744 );
xor ( n49746 , n49708 , n49745 );
and ( n49747 , n48552 , n48556 );
and ( n49748 , n48556 , n48562 );
and ( n49749 , n48552 , n48562 );
or ( n49750 , n49747 , n49748 , n49749 );
and ( n49751 , n48581 , n48586 );
and ( n49752 , n48586 , n48592 );
and ( n49753 , n48581 , n48592 );
or ( n49754 , n49751 , n49752 , n49753 );
xor ( n49755 , n49750 , n49754 );
and ( n49756 , n48558 , n48559 );
and ( n49757 , n48559 , n48561 );
and ( n49758 , n48558 , n48561 );
or ( n49759 , n49756 , n49757 , n49758 );
and ( n49760 , n48582 , n48583 );
and ( n49761 , n48583 , n48585 );
and ( n49762 , n48582 , n48585 );
or ( n49763 , n49760 , n49761 , n49762 );
xor ( n49764 , n49759 , n49763 );
and ( n49765 , n4132 , n22065 );
and ( n49766 , n4438 , n20976 );
xor ( n49767 , n49765 , n49766 );
and ( n49768 , n4766 , n20156 );
xor ( n49769 , n49767 , n49768 );
xor ( n49770 , n49764 , n49769 );
xor ( n49771 , n49755 , n49770 );
xor ( n49772 , n49746 , n49771 );
xor ( n49773 , n49704 , n49772 );
xor ( n49774 , n49695 , n49773 );
and ( n49775 , n48577 , n48593 );
and ( n49776 , n48593 , n48609 );
and ( n49777 , n48577 , n48609 );
or ( n49778 , n49775 , n49776 , n49777 );
and ( n49779 , n48615 , n48622 );
xor ( n49780 , n49778 , n49779 );
and ( n49781 , n48598 , n48602 );
and ( n49782 , n48602 , n48608 );
and ( n49783 , n48598 , n48608 );
or ( n49784 , n49781 , n49782 , n49783 );
and ( n49785 , n48588 , n48589 );
and ( n49786 , n48589 , n48591 );
and ( n49787 , n48588 , n48591 );
or ( n49788 , n49785 , n49786 , n49787 );
and ( n49789 , n3182 , n25163 );
and ( n49790 , n3545 , n24137 );
xor ( n49791 , n49789 , n49790 );
and ( n49792 , n3801 , n23075 );
xor ( n49793 , n49791 , n49792 );
xor ( n49794 , n49788 , n49793 );
and ( n49795 , n2462 , n28406 );
and ( n49796 , n2779 , n27296 );
xor ( n49797 , n49795 , n49796 );
and ( n49798 , n3024 , n26216 );
xor ( n49799 , n49797 , n49798 );
xor ( n49800 , n49794 , n49799 );
xor ( n49801 , n49784 , n49800 );
and ( n49802 , n48618 , n48619 );
and ( n49803 , n48619 , n48621 );
and ( n49804 , n48618 , n48621 );
or ( n49805 , n49802 , n49803 , n49804 );
and ( n49806 , n48604 , n48605 );
and ( n49807 , n48605 , n48607 );
and ( n49808 , n48604 , n48607 );
or ( n49809 , n49806 , n49807 , n49808 );
xor ( n49810 , n49805 , n49809 );
and ( n49811 , n1933 , n31761 );
and ( n49812 , n2120 , n30629 );
xor ( n49813 , n49811 , n49812 );
and ( n49814 , n2324 , n29508 );
xor ( n49815 , n49813 , n49814 );
xor ( n49816 , n49810 , n49815 );
xor ( n49817 , n49801 , n49816 );
xor ( n49818 , n49780 , n49817 );
not ( n49819 , n1580 );
and ( n49820 , n34193 , n1580 );
nor ( n49821 , n49819 , n49820 );
and ( n49822 , n1694 , n32999 );
xor ( n49823 , n49821 , n49822 );
xor ( n49824 , n49818 , n49823 );
xor ( n49825 , n49774 , n49824 );
xor ( n49826 , n49694 , n49825 );
xor ( n49827 , n49569 , n49826 );
xor ( n49828 , n49487 , n49827 );
xor ( n49829 , n49478 , n49828 );
and ( n49830 , n48267 , n48270 );
and ( n49831 , n48270 , n48628 );
and ( n49832 , n48267 , n48628 );
or ( n49833 , n49830 , n49831 , n49832 );
xor ( n49834 , n49829 , n49833 );
and ( n49835 , n48629 , n48633 );
and ( n49836 , n48634 , n48637 );
or ( n49837 , n49835 , n49836 );
xor ( n49838 , n49834 , n49837 );
buf ( n49839 , n49838 );
buf ( n49840 , n49839 );
not ( n49841 , n49840 );
nor ( n49842 , n49841 , n8739 );
xor ( n49843 , n49470 , n49842 );
and ( n49844 , n48263 , n48642 );
and ( n49845 , n48643 , n48646 );
or ( n49846 , n49844 , n49845 );
xor ( n49847 , n49843 , n49846 );
buf ( n49848 , n49847 );
buf ( n49849 , n49848 );
not ( n49850 , n49849 );
buf ( n49851 , n575 );
not ( n49852 , n49851 );
nor ( n49853 , n49850 , n49852 );
xor ( n49854 , n49096 , n49853 );
xor ( n49855 , n48658 , n49093 );
nor ( n49856 , n48650 , n49852 );
and ( n49857 , n49855 , n49856 );
xor ( n49858 , n49855 , n49856 );
xor ( n49859 , n48662 , n49091 );
nor ( n49860 , n47449 , n49852 );
and ( n49861 , n49859 , n49860 );
xor ( n49862 , n49859 , n49860 );
xor ( n49863 , n48666 , n49089 );
nor ( n49864 , n46248 , n49852 );
and ( n49865 , n49863 , n49864 );
xor ( n49866 , n49863 , n49864 );
xor ( n49867 , n48670 , n49087 );
nor ( n49868 , n45047 , n49852 );
and ( n49869 , n49867 , n49868 );
xor ( n49870 , n49867 , n49868 );
xor ( n49871 , n48674 , n49085 );
nor ( n49872 , n43843 , n49852 );
and ( n49873 , n49871 , n49872 );
xor ( n49874 , n49871 , n49872 );
xor ( n49875 , n48678 , n49083 );
nor ( n49876 , n42641 , n49852 );
and ( n49877 , n49875 , n49876 );
xor ( n49878 , n49875 , n49876 );
xor ( n49879 , n48682 , n49081 );
nor ( n49880 , n41437 , n49852 );
and ( n49881 , n49879 , n49880 );
xor ( n49882 , n49879 , n49880 );
xor ( n49883 , n48686 , n49079 );
nor ( n49884 , n40232 , n49852 );
and ( n49885 , n49883 , n49884 );
xor ( n49886 , n49883 , n49884 );
xor ( n49887 , n48690 , n49077 );
nor ( n49888 , n39027 , n49852 );
and ( n49889 , n49887 , n49888 );
xor ( n49890 , n49887 , n49888 );
xor ( n49891 , n48694 , n49075 );
nor ( n49892 , n37825 , n49852 );
and ( n49893 , n49891 , n49892 );
xor ( n49894 , n49891 , n49892 );
xor ( n49895 , n48698 , n49073 );
nor ( n49896 , n36620 , n49852 );
and ( n49897 , n49895 , n49896 );
xor ( n49898 , n49895 , n49896 );
xor ( n49899 , n48702 , n49071 );
nor ( n49900 , n35419 , n49852 );
and ( n49901 , n49899 , n49900 );
xor ( n49902 , n49899 , n49900 );
xor ( n49903 , n48706 , n49069 );
nor ( n49904 , n34224 , n49852 );
and ( n49905 , n49903 , n49904 );
xor ( n49906 , n49903 , n49904 );
xor ( n49907 , n48710 , n49067 );
nor ( n49908 , n33033 , n49852 );
and ( n49909 , n49907 , n49908 );
xor ( n49910 , n49907 , n49908 );
xor ( n49911 , n48714 , n49065 );
nor ( n49912 , n31867 , n49852 );
and ( n49913 , n49911 , n49912 );
xor ( n49914 , n49911 , n49912 );
xor ( n49915 , n48718 , n49063 );
nor ( n49916 , n30725 , n49852 );
and ( n49917 , n49915 , n49916 );
xor ( n49918 , n49915 , n49916 );
xor ( n49919 , n48722 , n49061 );
nor ( n49920 , n29596 , n49852 );
and ( n49921 , n49919 , n49920 );
xor ( n49922 , n49919 , n49920 );
xor ( n49923 , n48726 , n49059 );
nor ( n49924 , n28487 , n49852 );
and ( n49925 , n49923 , n49924 );
xor ( n49926 , n49923 , n49924 );
xor ( n49927 , n48730 , n49057 );
nor ( n49928 , n27397 , n49852 );
and ( n49929 , n49927 , n49928 );
xor ( n49930 , n49927 , n49928 );
xor ( n49931 , n48734 , n49055 );
nor ( n49932 , n26326 , n49852 );
and ( n49933 , n49931 , n49932 );
xor ( n49934 , n49931 , n49932 );
xor ( n49935 , n48738 , n49053 );
nor ( n49936 , n25272 , n49852 );
and ( n49937 , n49935 , n49936 );
xor ( n49938 , n49935 , n49936 );
xor ( n49939 , n48742 , n49051 );
nor ( n49940 , n24242 , n49852 );
and ( n49941 , n49939 , n49940 );
xor ( n49942 , n49939 , n49940 );
xor ( n49943 , n48746 , n49049 );
nor ( n49944 , n23225 , n49852 );
and ( n49945 , n49943 , n49944 );
xor ( n49946 , n49943 , n49944 );
xor ( n49947 , n48750 , n49047 );
nor ( n49948 , n22231 , n49852 );
and ( n49949 , n49947 , n49948 );
xor ( n49950 , n49947 , n49948 );
xor ( n49951 , n48754 , n49045 );
nor ( n49952 , n21258 , n49852 );
and ( n49953 , n49951 , n49952 );
xor ( n49954 , n49951 , n49952 );
xor ( n49955 , n48758 , n49043 );
nor ( n49956 , n20303 , n49852 );
and ( n49957 , n49955 , n49956 );
xor ( n49958 , n49955 , n49956 );
xor ( n49959 , n48762 , n49041 );
nor ( n49960 , n19365 , n49852 );
and ( n49961 , n49959 , n49960 );
xor ( n49962 , n49959 , n49960 );
xor ( n49963 , n48766 , n49039 );
nor ( n49964 , n18448 , n49852 );
and ( n49965 , n49963 , n49964 );
xor ( n49966 , n49963 , n49964 );
xor ( n49967 , n48770 , n49037 );
nor ( n49968 , n17548 , n49852 );
and ( n49969 , n49967 , n49968 );
xor ( n49970 , n49967 , n49968 );
xor ( n49971 , n48774 , n49035 );
nor ( n49972 , n16669 , n49852 );
and ( n49973 , n49971 , n49972 );
xor ( n49974 , n49971 , n49972 );
xor ( n49975 , n48778 , n49033 );
nor ( n49976 , n15809 , n49852 );
and ( n49977 , n49975 , n49976 );
xor ( n49978 , n49975 , n49976 );
xor ( n49979 , n48782 , n49031 );
nor ( n49980 , n14968 , n49852 );
and ( n49981 , n49979 , n49980 );
xor ( n49982 , n49979 , n49980 );
xor ( n49983 , n48786 , n49029 );
nor ( n49984 , n14147 , n49852 );
and ( n49985 , n49983 , n49984 );
xor ( n49986 , n49983 , n49984 );
xor ( n49987 , n48790 , n49027 );
nor ( n49988 , n13349 , n49852 );
and ( n49989 , n49987 , n49988 );
xor ( n49990 , n49987 , n49988 );
xor ( n49991 , n48794 , n49025 );
nor ( n49992 , n12564 , n49852 );
and ( n49993 , n49991 , n49992 );
xor ( n49994 , n49991 , n49992 );
xor ( n49995 , n48798 , n49023 );
nor ( n49996 , n11799 , n49852 );
and ( n49997 , n49995 , n49996 );
xor ( n49998 , n49995 , n49996 );
xor ( n49999 , n48802 , n49021 );
nor ( n50000 , n11050 , n49852 );
and ( n50001 , n49999 , n50000 );
xor ( n50002 , n49999 , n50000 );
xor ( n50003 , n48806 , n49019 );
nor ( n50004 , n10321 , n49852 );
and ( n50005 , n50003 , n50004 );
xor ( n50006 , n50003 , n50004 );
xor ( n50007 , n48810 , n49017 );
nor ( n50008 , n9429 , n49852 );
and ( n50009 , n50007 , n50008 );
xor ( n50010 , n50007 , n50008 );
xor ( n50011 , n48814 , n49015 );
nor ( n50012 , n8949 , n49852 );
and ( n50013 , n50011 , n50012 );
xor ( n50014 , n50011 , n50012 );
xor ( n50015 , n48818 , n49013 );
nor ( n50016 , n9437 , n49852 );
and ( n50017 , n50015 , n50016 );
xor ( n50018 , n50015 , n50016 );
xor ( n50019 , n48822 , n49011 );
nor ( n50020 , n9446 , n49852 );
and ( n50021 , n50019 , n50020 );
xor ( n50022 , n50019 , n50020 );
xor ( n50023 , n48826 , n49009 );
nor ( n50024 , n9455 , n49852 );
and ( n50025 , n50023 , n50024 );
xor ( n50026 , n50023 , n50024 );
xor ( n50027 , n48830 , n49007 );
nor ( n50028 , n9464 , n49852 );
and ( n50029 , n50027 , n50028 );
xor ( n50030 , n50027 , n50028 );
xor ( n50031 , n48834 , n49005 );
nor ( n50032 , n9473 , n49852 );
and ( n50033 , n50031 , n50032 );
xor ( n50034 , n50031 , n50032 );
xor ( n50035 , n48838 , n49003 );
nor ( n50036 , n9482 , n49852 );
and ( n50037 , n50035 , n50036 );
xor ( n50038 , n50035 , n50036 );
xor ( n50039 , n48842 , n49001 );
nor ( n50040 , n9491 , n49852 );
and ( n50041 , n50039 , n50040 );
xor ( n50042 , n50039 , n50040 );
xor ( n50043 , n48846 , n48999 );
nor ( n50044 , n9500 , n49852 );
and ( n50045 , n50043 , n50044 );
xor ( n50046 , n50043 , n50044 );
xor ( n50047 , n48850 , n48997 );
nor ( n50048 , n9509 , n49852 );
and ( n50049 , n50047 , n50048 );
xor ( n50050 , n50047 , n50048 );
xor ( n50051 , n48854 , n48995 );
nor ( n50052 , n9518 , n49852 );
and ( n50053 , n50051 , n50052 );
xor ( n50054 , n50051 , n50052 );
xor ( n50055 , n48858 , n48993 );
nor ( n50056 , n9527 , n49852 );
and ( n50057 , n50055 , n50056 );
xor ( n50058 , n50055 , n50056 );
xor ( n50059 , n48862 , n48991 );
nor ( n50060 , n9536 , n49852 );
and ( n50061 , n50059 , n50060 );
xor ( n50062 , n50059 , n50060 );
xor ( n50063 , n48866 , n48989 );
nor ( n50064 , n9545 , n49852 );
and ( n50065 , n50063 , n50064 );
xor ( n50066 , n50063 , n50064 );
xor ( n50067 , n48870 , n48987 );
nor ( n50068 , n9554 , n49852 );
and ( n50069 , n50067 , n50068 );
xor ( n50070 , n50067 , n50068 );
xor ( n50071 , n48874 , n48985 );
nor ( n50072 , n9563 , n49852 );
and ( n50073 , n50071 , n50072 );
xor ( n50074 , n50071 , n50072 );
xor ( n50075 , n48878 , n48983 );
nor ( n50076 , n9572 , n49852 );
and ( n50077 , n50075 , n50076 );
xor ( n50078 , n50075 , n50076 );
xor ( n50079 , n48882 , n48981 );
nor ( n50080 , n9581 , n49852 );
and ( n50081 , n50079 , n50080 );
xor ( n50082 , n50079 , n50080 );
xor ( n50083 , n48886 , n48979 );
nor ( n50084 , n9590 , n49852 );
and ( n50085 , n50083 , n50084 );
xor ( n50086 , n50083 , n50084 );
xor ( n50087 , n48890 , n48977 );
nor ( n50088 , n9599 , n49852 );
and ( n50089 , n50087 , n50088 );
xor ( n50090 , n50087 , n50088 );
xor ( n50091 , n48894 , n48975 );
nor ( n50092 , n9608 , n49852 );
and ( n50093 , n50091 , n50092 );
xor ( n50094 , n50091 , n50092 );
xor ( n50095 , n48898 , n48973 );
nor ( n50096 , n9617 , n49852 );
and ( n50097 , n50095 , n50096 );
xor ( n50098 , n50095 , n50096 );
xor ( n50099 , n48902 , n48971 );
nor ( n50100 , n9626 , n49852 );
and ( n50101 , n50099 , n50100 );
xor ( n50102 , n50099 , n50100 );
xor ( n50103 , n48906 , n48969 );
nor ( n50104 , n9635 , n49852 );
and ( n50105 , n50103 , n50104 );
xor ( n50106 , n50103 , n50104 );
xor ( n50107 , n48910 , n48967 );
nor ( n50108 , n9644 , n49852 );
and ( n50109 , n50107 , n50108 );
xor ( n50110 , n50107 , n50108 );
xor ( n50111 , n48914 , n48965 );
nor ( n50112 , n9653 , n49852 );
and ( n50113 , n50111 , n50112 );
xor ( n50114 , n50111 , n50112 );
xor ( n50115 , n48918 , n48963 );
nor ( n50116 , n9662 , n49852 );
and ( n50117 , n50115 , n50116 );
xor ( n50118 , n50115 , n50116 );
xor ( n50119 , n48922 , n48961 );
nor ( n50120 , n9671 , n49852 );
and ( n50121 , n50119 , n50120 );
xor ( n50122 , n50119 , n50120 );
xor ( n50123 , n48926 , n48959 );
nor ( n50124 , n9680 , n49852 );
and ( n50125 , n50123 , n50124 );
xor ( n50126 , n50123 , n50124 );
xor ( n50127 , n48930 , n48957 );
nor ( n50128 , n9689 , n49852 );
and ( n50129 , n50127 , n50128 );
xor ( n50130 , n50127 , n50128 );
xor ( n50131 , n48934 , n48955 );
nor ( n50132 , n9698 , n49852 );
and ( n50133 , n50131 , n50132 );
xor ( n50134 , n50131 , n50132 );
xor ( n50135 , n48938 , n48953 );
nor ( n50136 , n9707 , n49852 );
and ( n50137 , n50135 , n50136 );
xor ( n50138 , n50135 , n50136 );
xor ( n50139 , n48942 , n48951 );
nor ( n50140 , n9716 , n49852 );
and ( n50141 , n50139 , n50140 );
xor ( n50142 , n50139 , n50140 );
xor ( n50143 , n48946 , n48949 );
nor ( n50144 , n9725 , n49852 );
and ( n50145 , n50143 , n50144 );
xor ( n50146 , n50143 , n50144 );
xor ( n50147 , n48947 , n48948 );
nor ( n50148 , n9734 , n49852 );
and ( n50149 , n50147 , n50148 );
xor ( n50150 , n50147 , n50148 );
nor ( n50151 , n9752 , n48652 );
nor ( n50152 , n9743 , n49852 );
and ( n50153 , n50151 , n50152 );
and ( n50154 , n50150 , n50153 );
or ( n50155 , n50149 , n50154 );
and ( n50156 , n50146 , n50155 );
or ( n50157 , n50145 , n50156 );
and ( n50158 , n50142 , n50157 );
or ( n50159 , n50141 , n50158 );
and ( n50160 , n50138 , n50159 );
or ( n50161 , n50137 , n50160 );
and ( n50162 , n50134 , n50161 );
or ( n50163 , n50133 , n50162 );
and ( n50164 , n50130 , n50163 );
or ( n50165 , n50129 , n50164 );
and ( n50166 , n50126 , n50165 );
or ( n50167 , n50125 , n50166 );
and ( n50168 , n50122 , n50167 );
or ( n50169 , n50121 , n50168 );
and ( n50170 , n50118 , n50169 );
or ( n50171 , n50117 , n50170 );
and ( n50172 , n50114 , n50171 );
or ( n50173 , n50113 , n50172 );
and ( n50174 , n50110 , n50173 );
or ( n50175 , n50109 , n50174 );
and ( n50176 , n50106 , n50175 );
or ( n50177 , n50105 , n50176 );
and ( n50178 , n50102 , n50177 );
or ( n50179 , n50101 , n50178 );
and ( n50180 , n50098 , n50179 );
or ( n50181 , n50097 , n50180 );
and ( n50182 , n50094 , n50181 );
or ( n50183 , n50093 , n50182 );
and ( n50184 , n50090 , n50183 );
or ( n50185 , n50089 , n50184 );
and ( n50186 , n50086 , n50185 );
or ( n50187 , n50085 , n50186 );
and ( n50188 , n50082 , n50187 );
or ( n50189 , n50081 , n50188 );
and ( n50190 , n50078 , n50189 );
or ( n50191 , n50077 , n50190 );
and ( n50192 , n50074 , n50191 );
or ( n50193 , n50073 , n50192 );
and ( n50194 , n50070 , n50193 );
or ( n50195 , n50069 , n50194 );
and ( n50196 , n50066 , n50195 );
or ( n50197 , n50065 , n50196 );
and ( n50198 , n50062 , n50197 );
or ( n50199 , n50061 , n50198 );
and ( n50200 , n50058 , n50199 );
or ( n50201 , n50057 , n50200 );
and ( n50202 , n50054 , n50201 );
or ( n50203 , n50053 , n50202 );
and ( n50204 , n50050 , n50203 );
or ( n50205 , n50049 , n50204 );
and ( n50206 , n50046 , n50205 );
or ( n50207 , n50045 , n50206 );
and ( n50208 , n50042 , n50207 );
or ( n50209 , n50041 , n50208 );
and ( n50210 , n50038 , n50209 );
or ( n50211 , n50037 , n50210 );
and ( n50212 , n50034 , n50211 );
or ( n50213 , n50033 , n50212 );
and ( n50214 , n50030 , n50213 );
or ( n50215 , n50029 , n50214 );
and ( n50216 , n50026 , n50215 );
or ( n50217 , n50025 , n50216 );
and ( n50218 , n50022 , n50217 );
or ( n50219 , n50021 , n50218 );
and ( n50220 , n50018 , n50219 );
or ( n50221 , n50017 , n50220 );
and ( n50222 , n50014 , n50221 );
or ( n50223 , n50013 , n50222 );
and ( n50224 , n50010 , n50223 );
or ( n50225 , n50009 , n50224 );
and ( n50226 , n50006 , n50225 );
or ( n50227 , n50005 , n50226 );
and ( n50228 , n50002 , n50227 );
or ( n50229 , n50001 , n50228 );
and ( n50230 , n49998 , n50229 );
or ( n50231 , n49997 , n50230 );
and ( n50232 , n49994 , n50231 );
or ( n50233 , n49993 , n50232 );
and ( n50234 , n49990 , n50233 );
or ( n50235 , n49989 , n50234 );
and ( n50236 , n49986 , n50235 );
or ( n50237 , n49985 , n50236 );
and ( n50238 , n49982 , n50237 );
or ( n50239 , n49981 , n50238 );
and ( n50240 , n49978 , n50239 );
or ( n50241 , n49977 , n50240 );
and ( n50242 , n49974 , n50241 );
or ( n50243 , n49973 , n50242 );
and ( n50244 , n49970 , n50243 );
or ( n50245 , n49969 , n50244 );
and ( n50246 , n49966 , n50245 );
or ( n50247 , n49965 , n50246 );
and ( n50248 , n49962 , n50247 );
or ( n50249 , n49961 , n50248 );
and ( n50250 , n49958 , n50249 );
or ( n50251 , n49957 , n50250 );
and ( n50252 , n49954 , n50251 );
or ( n50253 , n49953 , n50252 );
and ( n50254 , n49950 , n50253 );
or ( n50255 , n49949 , n50254 );
and ( n50256 , n49946 , n50255 );
or ( n50257 , n49945 , n50256 );
and ( n50258 , n49942 , n50257 );
or ( n50259 , n49941 , n50258 );
and ( n50260 , n49938 , n50259 );
or ( n50261 , n49937 , n50260 );
and ( n50262 , n49934 , n50261 );
or ( n50263 , n49933 , n50262 );
and ( n50264 , n49930 , n50263 );
or ( n50265 , n49929 , n50264 );
and ( n50266 , n49926 , n50265 );
or ( n50267 , n49925 , n50266 );
and ( n50268 , n49922 , n50267 );
or ( n50269 , n49921 , n50268 );
and ( n50270 , n49918 , n50269 );
or ( n50271 , n49917 , n50270 );
and ( n50272 , n49914 , n50271 );
or ( n50273 , n49913 , n50272 );
and ( n50274 , n49910 , n50273 );
or ( n50275 , n49909 , n50274 );
and ( n50276 , n49906 , n50275 );
or ( n50277 , n49905 , n50276 );
and ( n50278 , n49902 , n50277 );
or ( n50279 , n49901 , n50278 );
and ( n50280 , n49898 , n50279 );
or ( n50281 , n49897 , n50280 );
and ( n50282 , n49894 , n50281 );
or ( n50283 , n49893 , n50282 );
and ( n50284 , n49890 , n50283 );
or ( n50285 , n49889 , n50284 );
and ( n50286 , n49886 , n50285 );
or ( n50287 , n49885 , n50286 );
and ( n50288 , n49882 , n50287 );
or ( n50289 , n49881 , n50288 );
and ( n50290 , n49878 , n50289 );
or ( n50291 , n49877 , n50290 );
and ( n50292 , n49874 , n50291 );
or ( n50293 , n49873 , n50292 );
and ( n50294 , n49870 , n50293 );
or ( n50295 , n49869 , n50294 );
and ( n50296 , n49866 , n50295 );
or ( n50297 , n49865 , n50296 );
and ( n50298 , n49862 , n50297 );
or ( n50299 , n49861 , n50298 );
and ( n50300 , n49858 , n50299 );
or ( n50301 , n49857 , n50300 );
xor ( n50302 , n49854 , n50301 );
and ( n50303 , n33403 , n1765 );
nor ( n50304 , n1766 , n50303 );
nor ( n50305 , n1945 , n32231 );
xor ( n50306 , n50304 , n50305 );
and ( n50307 , n49098 , n49099 );
and ( n50308 , n49100 , n49103 );
or ( n50309 , n50307 , n50308 );
xor ( n50310 , n50306 , n50309 );
nor ( n50311 , n2137 , n31083 );
xor ( n50312 , n50310 , n50311 );
and ( n50313 , n49104 , n49105 );
and ( n50314 , n49106 , n49109 );
or ( n50315 , n50313 , n50314 );
xor ( n50316 , n50312 , n50315 );
nor ( n50317 , n2343 , n29948 );
xor ( n50318 , n50316 , n50317 );
and ( n50319 , n49110 , n49111 );
and ( n50320 , n49112 , n49115 );
or ( n50321 , n50319 , n50320 );
xor ( n50322 , n50318 , n50321 );
nor ( n50323 , n2566 , n28833 );
xor ( n50324 , n50322 , n50323 );
and ( n50325 , n49116 , n49117 );
and ( n50326 , n49118 , n49121 );
or ( n50327 , n50325 , n50326 );
xor ( n50328 , n50324 , n50327 );
nor ( n50329 , n2797 , n27737 );
xor ( n50330 , n50328 , n50329 );
and ( n50331 , n49122 , n49123 );
and ( n50332 , n49124 , n49127 );
or ( n50333 , n50331 , n50332 );
xor ( n50334 , n50330 , n50333 );
nor ( n50335 , n3043 , n26660 );
xor ( n50336 , n50334 , n50335 );
and ( n50337 , n49128 , n49129 );
and ( n50338 , n49130 , n49133 );
or ( n50339 , n50337 , n50338 );
xor ( n50340 , n50336 , n50339 );
nor ( n50341 , n3300 , n25600 );
xor ( n50342 , n50340 , n50341 );
and ( n50343 , n49134 , n49135 );
and ( n50344 , n49136 , n49139 );
or ( n50345 , n50343 , n50344 );
xor ( n50346 , n50342 , n50345 );
nor ( n50347 , n3570 , n24564 );
xor ( n50348 , n50346 , n50347 );
and ( n50349 , n49140 , n49141 );
and ( n50350 , n49142 , n49145 );
or ( n50351 , n50349 , n50350 );
xor ( n50352 , n50348 , n50351 );
nor ( n50353 , n3853 , n23541 );
xor ( n50354 , n50352 , n50353 );
and ( n50355 , n49146 , n49147 );
and ( n50356 , n49148 , n49151 );
or ( n50357 , n50355 , n50356 );
xor ( n50358 , n50354 , n50357 );
nor ( n50359 , n4151 , n22541 );
xor ( n50360 , n50358 , n50359 );
and ( n50361 , n49152 , n49153 );
and ( n50362 , n49154 , n49157 );
or ( n50363 , n50361 , n50362 );
xor ( n50364 , n50360 , n50363 );
nor ( n50365 , n4458 , n21562 );
xor ( n50366 , n50364 , n50365 );
and ( n50367 , n49158 , n49159 );
and ( n50368 , n49160 , n49163 );
or ( n50369 , n50367 , n50368 );
xor ( n50370 , n50366 , n50369 );
nor ( n50371 , n4786 , n20601 );
xor ( n50372 , n50370 , n50371 );
and ( n50373 , n49164 , n49165 );
and ( n50374 , n49166 , n49169 );
or ( n50375 , n50373 , n50374 );
xor ( n50376 , n50372 , n50375 );
nor ( n50377 , n5126 , n19657 );
xor ( n50378 , n50376 , n50377 );
and ( n50379 , n49170 , n49171 );
and ( n50380 , n49172 , n49175 );
or ( n50381 , n50379 , n50380 );
xor ( n50382 , n50378 , n50381 );
nor ( n50383 , n5477 , n18734 );
xor ( n50384 , n50382 , n50383 );
and ( n50385 , n49176 , n49177 );
and ( n50386 , n49178 , n49181 );
or ( n50387 , n50385 , n50386 );
xor ( n50388 , n50384 , n50387 );
nor ( n50389 , n5838 , n17828 );
xor ( n50390 , n50388 , n50389 );
and ( n50391 , n49182 , n49183 );
and ( n50392 , n49184 , n49187 );
or ( n50393 , n50391 , n50392 );
xor ( n50394 , n50390 , n50393 );
nor ( n50395 , n6212 , n16943 );
xor ( n50396 , n50394 , n50395 );
and ( n50397 , n49188 , n49189 );
and ( n50398 , n49190 , n49193 );
or ( n50399 , n50397 , n50398 );
xor ( n50400 , n50396 , n50399 );
nor ( n50401 , n6596 , n16077 );
xor ( n50402 , n50400 , n50401 );
and ( n50403 , n49194 , n49195 );
and ( n50404 , n49196 , n49199 );
or ( n50405 , n50403 , n50404 );
xor ( n50406 , n50402 , n50405 );
nor ( n50407 , n6997 , n15230 );
xor ( n50408 , n50406 , n50407 );
and ( n50409 , n49200 , n49201 );
and ( n50410 , n49202 , n49205 );
or ( n50411 , n50409 , n50410 );
xor ( n50412 , n50408 , n50411 );
nor ( n50413 , n7413 , n14403 );
xor ( n50414 , n50412 , n50413 );
and ( n50415 , n49206 , n49207 );
and ( n50416 , n49208 , n49211 );
or ( n50417 , n50415 , n50416 );
xor ( n50418 , n50414 , n50417 );
nor ( n50419 , n7841 , n13599 );
xor ( n50420 , n50418 , n50419 );
and ( n50421 , n49212 , n49213 );
and ( n50422 , n49214 , n49217 );
or ( n50423 , n50421 , n50422 );
xor ( n50424 , n50420 , n50423 );
nor ( n50425 , n8281 , n12808 );
xor ( n50426 , n50424 , n50425 );
and ( n50427 , n49218 , n49219 );
and ( n50428 , n49220 , n49223 );
or ( n50429 , n50427 , n50428 );
xor ( n50430 , n50426 , n50429 );
nor ( n50431 , n8737 , n12037 );
xor ( n50432 , n50430 , n50431 );
and ( n50433 , n49224 , n49225 );
and ( n50434 , n49226 , n49229 );
or ( n50435 , n50433 , n50434 );
xor ( n50436 , n50432 , n50435 );
nor ( n50437 , n9420 , n11282 );
xor ( n50438 , n50436 , n50437 );
and ( n50439 , n49230 , n49231 );
and ( n50440 , n49232 , n49235 );
or ( n50441 , n50439 , n50440 );
xor ( n50442 , n50438 , n50441 );
nor ( n50443 , n10312 , n10547 );
xor ( n50444 , n50442 , n50443 );
and ( n50445 , n49236 , n49237 );
and ( n50446 , n49238 , n49241 );
or ( n50447 , n50445 , n50446 );
xor ( n50448 , n50444 , n50447 );
nor ( n50449 , n11041 , n9829 );
xor ( n50450 , n50448 , n50449 );
and ( n50451 , n49242 , n49243 );
and ( n50452 , n49244 , n49247 );
or ( n50453 , n50451 , n50452 );
xor ( n50454 , n50450 , n50453 );
nor ( n50455 , n11790 , n8955 );
xor ( n50456 , n50454 , n50455 );
and ( n50457 , n49248 , n49249 );
and ( n50458 , n49250 , n49253 );
or ( n50459 , n50457 , n50458 );
xor ( n50460 , n50456 , n50459 );
nor ( n50461 , n12555 , n603 );
xor ( n50462 , n50460 , n50461 );
and ( n50463 , n49254 , n49255 );
and ( n50464 , n49256 , n49259 );
or ( n50465 , n50463 , n50464 );
xor ( n50466 , n50462 , n50465 );
nor ( n50467 , n13340 , n652 );
xor ( n50468 , n50466 , n50467 );
and ( n50469 , n49260 , n49261 );
and ( n50470 , n49262 , n49265 );
or ( n50471 , n50469 , n50470 );
xor ( n50472 , n50468 , n50471 );
nor ( n50473 , n14138 , n624 );
xor ( n50474 , n50472 , n50473 );
and ( n50475 , n49266 , n49267 );
and ( n50476 , n49268 , n49271 );
or ( n50477 , n50475 , n50476 );
xor ( n50478 , n50474 , n50477 );
nor ( n50479 , n14959 , n648 );
xor ( n50480 , n50478 , n50479 );
and ( n50481 , n49272 , n49273 );
and ( n50482 , n49274 , n49277 );
or ( n50483 , n50481 , n50482 );
xor ( n50484 , n50480 , n50483 );
nor ( n50485 , n15800 , n686 );
xor ( n50486 , n50484 , n50485 );
and ( n50487 , n49278 , n49279 );
and ( n50488 , n49280 , n49283 );
or ( n50489 , n50487 , n50488 );
xor ( n50490 , n50486 , n50489 );
nor ( n50491 , n16660 , n735 );
xor ( n50492 , n50490 , n50491 );
and ( n50493 , n49284 , n49285 );
and ( n50494 , n49286 , n49289 );
or ( n50495 , n50493 , n50494 );
xor ( n50496 , n50492 , n50495 );
nor ( n50497 , n17539 , n798 );
xor ( n50498 , n50496 , n50497 );
and ( n50499 , n49290 , n49291 );
and ( n50500 , n49292 , n49295 );
or ( n50501 , n50499 , n50500 );
xor ( n50502 , n50498 , n50501 );
nor ( n50503 , n18439 , n870 );
xor ( n50504 , n50502 , n50503 );
and ( n50505 , n49296 , n49297 );
and ( n50506 , n49298 , n49301 );
or ( n50507 , n50505 , n50506 );
xor ( n50508 , n50504 , n50507 );
nor ( n50509 , n19356 , n960 );
xor ( n50510 , n50508 , n50509 );
and ( n50511 , n49302 , n49303 );
and ( n50512 , n49304 , n49307 );
or ( n50513 , n50511 , n50512 );
xor ( n50514 , n50510 , n50513 );
nor ( n50515 , n20294 , n1064 );
xor ( n50516 , n50514 , n50515 );
and ( n50517 , n49308 , n49309 );
and ( n50518 , n49310 , n49313 );
or ( n50519 , n50517 , n50518 );
xor ( n50520 , n50516 , n50519 );
nor ( n50521 , n21249 , n1178 );
xor ( n50522 , n50520 , n50521 );
and ( n50523 , n49314 , n49315 );
and ( n50524 , n49316 , n49319 );
or ( n50525 , n50523 , n50524 );
xor ( n50526 , n50522 , n50525 );
nor ( n50527 , n22222 , n1305 );
xor ( n50528 , n50526 , n50527 );
and ( n50529 , n49320 , n49321 );
and ( n50530 , n49322 , n49325 );
or ( n50531 , n50529 , n50530 );
xor ( n50532 , n50528 , n50531 );
nor ( n50533 , n23216 , n1447 );
xor ( n50534 , n50532 , n50533 );
and ( n50535 , n49326 , n49327 );
and ( n50536 , n49328 , n49331 );
or ( n50537 , n50535 , n50536 );
xor ( n50538 , n50534 , n50537 );
nor ( n50539 , n24233 , n1600 );
xor ( n50540 , n50538 , n50539 );
and ( n50541 , n49332 , n49333 );
and ( n50542 , n49334 , n49337 );
or ( n50543 , n50541 , n50542 );
xor ( n50544 , n50540 , n50543 );
nor ( n50545 , n25263 , n1768 );
xor ( n50546 , n50544 , n50545 );
and ( n50547 , n49338 , n49339 );
and ( n50548 , n49340 , n49343 );
or ( n50549 , n50547 , n50548 );
xor ( n50550 , n50546 , n50549 );
nor ( n50551 , n26317 , n1947 );
xor ( n50552 , n50550 , n50551 );
and ( n50553 , n49344 , n49345 );
and ( n50554 , n49346 , n49349 );
or ( n50555 , n50553 , n50554 );
xor ( n50556 , n50552 , n50555 );
nor ( n50557 , n27388 , n2139 );
xor ( n50558 , n50556 , n50557 );
and ( n50559 , n49350 , n49351 );
and ( n50560 , n49352 , n49355 );
or ( n50561 , n50559 , n50560 );
xor ( n50562 , n50558 , n50561 );
nor ( n50563 , n28478 , n2345 );
xor ( n50564 , n50562 , n50563 );
and ( n50565 , n49356 , n49357 );
and ( n50566 , n49358 , n49361 );
or ( n50567 , n50565 , n50566 );
xor ( n50568 , n50564 , n50567 );
nor ( n50569 , n29587 , n2568 );
xor ( n50570 , n50568 , n50569 );
and ( n50571 , n49362 , n49363 );
and ( n50572 , n49364 , n49367 );
or ( n50573 , n50571 , n50572 );
xor ( n50574 , n50570 , n50573 );
nor ( n50575 , n30716 , n2799 );
xor ( n50576 , n50574 , n50575 );
and ( n50577 , n49368 , n49369 );
and ( n50578 , n49370 , n49373 );
or ( n50579 , n50577 , n50578 );
xor ( n50580 , n50576 , n50579 );
nor ( n50581 , n31858 , n3045 );
xor ( n50582 , n50580 , n50581 );
and ( n50583 , n49374 , n49375 );
and ( n50584 , n49376 , n49379 );
or ( n50585 , n50583 , n50584 );
xor ( n50586 , n50582 , n50585 );
nor ( n50587 , n33024 , n3302 );
xor ( n50588 , n50586 , n50587 );
and ( n50589 , n49380 , n49381 );
and ( n50590 , n49382 , n49385 );
or ( n50591 , n50589 , n50590 );
xor ( n50592 , n50588 , n50591 );
nor ( n50593 , n34215 , n3572 );
xor ( n50594 , n50592 , n50593 );
and ( n50595 , n49386 , n49387 );
and ( n50596 , n49388 , n49391 );
or ( n50597 , n50595 , n50596 );
xor ( n50598 , n50594 , n50597 );
nor ( n50599 , n35410 , n3855 );
xor ( n50600 , n50598 , n50599 );
and ( n50601 , n49392 , n49393 );
and ( n50602 , n49394 , n49397 );
or ( n50603 , n50601 , n50602 );
xor ( n50604 , n50600 , n50603 );
nor ( n50605 , n36611 , n4153 );
xor ( n50606 , n50604 , n50605 );
and ( n50607 , n49398 , n49399 );
and ( n50608 , n49400 , n49403 );
or ( n50609 , n50607 , n50608 );
xor ( n50610 , n50606 , n50609 );
nor ( n50611 , n37816 , n4460 );
xor ( n50612 , n50610 , n50611 );
and ( n50613 , n49404 , n49405 );
and ( n50614 , n49406 , n49409 );
or ( n50615 , n50613 , n50614 );
xor ( n50616 , n50612 , n50615 );
nor ( n50617 , n39018 , n4788 );
xor ( n50618 , n50616 , n50617 );
and ( n50619 , n49410 , n49411 );
and ( n50620 , n49412 , n49415 );
or ( n50621 , n50619 , n50620 );
xor ( n50622 , n50618 , n50621 );
nor ( n50623 , n40223 , n5128 );
xor ( n50624 , n50622 , n50623 );
and ( n50625 , n49416 , n49417 );
and ( n50626 , n49418 , n49421 );
or ( n50627 , n50625 , n50626 );
xor ( n50628 , n50624 , n50627 );
nor ( n50629 , n41428 , n5479 );
xor ( n50630 , n50628 , n50629 );
and ( n50631 , n49422 , n49423 );
and ( n50632 , n49424 , n49427 );
or ( n50633 , n50631 , n50632 );
xor ( n50634 , n50630 , n50633 );
nor ( n50635 , n42632 , n5840 );
xor ( n50636 , n50634 , n50635 );
and ( n50637 , n49428 , n49429 );
and ( n50638 , n49430 , n49433 );
or ( n50639 , n50637 , n50638 );
xor ( n50640 , n50636 , n50639 );
nor ( n50641 , n43834 , n6214 );
xor ( n50642 , n50640 , n50641 );
and ( n50643 , n49434 , n49435 );
and ( n50644 , n49436 , n49439 );
or ( n50645 , n50643 , n50644 );
xor ( n50646 , n50642 , n50645 );
nor ( n50647 , n45038 , n6598 );
xor ( n50648 , n50646 , n50647 );
and ( n50649 , n49440 , n49441 );
and ( n50650 , n49442 , n49445 );
or ( n50651 , n50649 , n50650 );
xor ( n50652 , n50648 , n50651 );
nor ( n50653 , n46239 , n6999 );
xor ( n50654 , n50652 , n50653 );
and ( n50655 , n49446 , n49447 );
and ( n50656 , n49448 , n49451 );
or ( n50657 , n50655 , n50656 );
xor ( n50658 , n50654 , n50657 );
nor ( n50659 , n47440 , n7415 );
xor ( n50660 , n50658 , n50659 );
and ( n50661 , n49452 , n49453 );
and ( n50662 , n49454 , n49457 );
or ( n50663 , n50661 , n50662 );
xor ( n50664 , n50660 , n50663 );
nor ( n50665 , n48641 , n7843 );
xor ( n50666 , n50664 , n50665 );
and ( n50667 , n49458 , n49459 );
and ( n50668 , n49460 , n49463 );
or ( n50669 , n50667 , n50668 );
xor ( n50670 , n50666 , n50669 );
nor ( n50671 , n49841 , n8283 );
xor ( n50672 , n50670 , n50671 );
and ( n50673 , n49464 , n49465 );
and ( n50674 , n49466 , n49469 );
or ( n50675 , n50673 , n50674 );
xor ( n50676 , n50672 , n50675 );
and ( n50677 , n49482 , n49486 );
and ( n50678 , n49486 , n49827 );
and ( n50679 , n49482 , n49827 );
or ( n50680 , n50677 , n50678 , n50679 );
and ( n50681 , n33774 , n1738 );
not ( n50682 , n1738 );
nor ( n50683 , n50681 , n50682 );
xor ( n50684 , n50680 , n50683 );
and ( n50685 , n49495 , n49499 );
and ( n50686 , n49499 , n49567 );
and ( n50687 , n49495 , n49567 );
or ( n50688 , n50685 , n50686 , n50687 );
and ( n50689 , n49491 , n49568 );
and ( n50690 , n49568 , n49826 );
and ( n50691 , n49491 , n49826 );
or ( n50692 , n50689 , n50690 , n50691 );
xor ( n50693 , n50688 , n50692 );
and ( n50694 , n49573 , n49693 );
and ( n50695 , n49693 , n49825 );
and ( n50696 , n49573 , n49825 );
or ( n50697 , n50694 , n50695 , n50696 );
and ( n50698 , n49504 , n49508 );
and ( n50699 , n49508 , n49566 );
and ( n50700 , n49504 , n49566 );
or ( n50701 , n50698 , n50699 , n50700 );
and ( n50702 , n49577 , n49581 );
and ( n50703 , n49581 , n49692 );
and ( n50704 , n49577 , n49692 );
or ( n50705 , n50702 , n50703 , n50704 );
xor ( n50706 , n50701 , n50705 );
and ( n50707 , n49535 , n49539 );
and ( n50708 , n49539 , n49545 );
and ( n50709 , n49535 , n49545 );
or ( n50710 , n50707 , n50708 , n50709 );
and ( n50711 , n49513 , n49517 );
and ( n50712 , n49517 , n49565 );
and ( n50713 , n49513 , n49565 );
or ( n50714 , n50711 , n50712 , n50713 );
xor ( n50715 , n50710 , n50714 );
and ( n50716 , n49522 , n49526 );
and ( n50717 , n49526 , n49564 );
and ( n50718 , n49522 , n49564 );
or ( n50719 , n50716 , n50717 , n50718 );
and ( n50720 , n49590 , n49615 );
and ( n50721 , n49615 , n49653 );
and ( n50722 , n49590 , n49653 );
or ( n50723 , n50720 , n50721 , n50722 );
xor ( n50724 , n50719 , n50723 );
and ( n50725 , n49531 , n49546 );
and ( n50726 , n49546 , n49563 );
and ( n50727 , n49531 , n49563 );
or ( n50728 , n50725 , n50726 , n50727 );
and ( n50729 , n49594 , n49598 );
and ( n50730 , n49598 , n49614 );
and ( n50731 , n49594 , n49614 );
or ( n50732 , n50729 , n50730 , n50731 );
xor ( n50733 , n50728 , n50732 );
and ( n50734 , n49551 , n49556 );
and ( n50735 , n49556 , n49562 );
and ( n50736 , n49551 , n49562 );
or ( n50737 , n50734 , n50735 , n50736 );
and ( n50738 , n49541 , n49542 );
and ( n50739 , n49542 , n49544 );
and ( n50740 , n49541 , n49544 );
or ( n50741 , n50738 , n50739 , n50740 );
and ( n50742 , n49552 , n49553 );
and ( n50743 , n49553 , n49555 );
and ( n50744 , n49552 , n49555 );
or ( n50745 , n50742 , n50743 , n50744 );
xor ( n50746 , n50741 , n50745 );
and ( n50747 , n30695 , n2298 );
and ( n50748 , n31836 , n2100 );
xor ( n50749 , n50747 , n50748 );
and ( n50750 , n32649 , n1882 );
xor ( n50751 , n50749 , n50750 );
xor ( n50752 , n50746 , n50751 );
xor ( n50753 , n50737 , n50752 );
and ( n50754 , n49558 , n49559 );
and ( n50755 , n49559 , n49561 );
and ( n50756 , n49558 , n49561 );
or ( n50757 , n50754 , n50755 , n50756 );
and ( n50758 , n27361 , n2981 );
and ( n50759 , n28456 , n2739 );
xor ( n50760 , n50758 , n50759 );
and ( n50761 , n29559 , n2544 );
xor ( n50762 , n50760 , n50761 );
xor ( n50763 , n50757 , n50762 );
and ( n50764 , n24214 , n3749 );
and ( n50765 , n25243 , n3495 );
xor ( n50766 , n50764 , n50765 );
and ( n50767 , n26296 , n3271 );
xor ( n50768 , n50766 , n50767 );
xor ( n50769 , n50763 , n50768 );
xor ( n50770 , n50753 , n50769 );
xor ( n50771 , n50733 , n50770 );
xor ( n50772 , n50724 , n50771 );
xor ( n50773 , n50715 , n50772 );
xor ( n50774 , n50706 , n50773 );
xor ( n50775 , n50697 , n50774 );
and ( n50776 , n49695 , n49773 );
and ( n50777 , n49773 , n49824 );
and ( n50778 , n49695 , n49824 );
or ( n50779 , n50776 , n50777 , n50778 );
and ( n50780 , n49586 , n49654 );
and ( n50781 , n49654 , n49691 );
and ( n50782 , n49586 , n49691 );
or ( n50783 , n50780 , n50781 , n50782 );
and ( n50784 , n49699 , n49703 );
and ( n50785 , n49703 , n49772 );
and ( n50786 , n49699 , n49772 );
or ( n50787 , n50784 , n50785 , n50786 );
xor ( n50788 , n50783 , n50787 );
and ( n50789 , n49659 , n49663 );
and ( n50790 , n49663 , n49690 );
and ( n50791 , n49659 , n49690 );
or ( n50792 , n50789 , n50790 , n50791 );
and ( n50793 , n49620 , n49636 );
and ( n50794 , n49636 , n49652 );
and ( n50795 , n49620 , n49652 );
or ( n50796 , n50793 , n50794 , n50795 );
and ( n50797 , n49603 , n49607 );
and ( n50798 , n49607 , n49613 );
and ( n50799 , n49603 , n49613 );
or ( n50800 , n50797 , n50798 , n50799 );
and ( n50801 , n49624 , n49629 );
and ( n50802 , n49629 , n49635 );
and ( n50803 , n49624 , n49635 );
or ( n50804 , n50801 , n50802 , n50803 );
xor ( n50805 , n50800 , n50804 );
and ( n50806 , n49609 , n49610 );
and ( n50807 , n49610 , n49612 );
and ( n50808 , n49609 , n49612 );
or ( n50809 , n50806 , n50807 , n50808 );
and ( n50810 , n49625 , n49626 );
and ( n50811 , n49626 , n49628 );
and ( n50812 , n49625 , n49628 );
or ( n50813 , n50810 , n50811 , n50812 );
xor ( n50814 , n50809 , n50813 );
and ( n50815 , n21216 , n4730 );
and ( n50816 , n22186 , n4403 );
xor ( n50817 , n50815 , n50816 );
and ( n50818 , n22892 , n4102 );
xor ( n50819 , n50817 , n50818 );
xor ( n50820 , n50814 , n50819 );
xor ( n50821 , n50805 , n50820 );
xor ( n50822 , n50796 , n50821 );
and ( n50823 , n49641 , n49645 );
and ( n50824 , n49645 , n49651 );
and ( n50825 , n49641 , n49651 );
or ( n50826 , n50823 , n50824 , n50825 );
and ( n50827 , n49631 , n49632 );
and ( n50828 , n49632 , n49634 );
and ( n50829 , n49631 , n49634 );
or ( n50830 , n50827 , n50828 , n50829 );
and ( n50831 , n18144 , n5765 );
and ( n50832 , n19324 , n5408 );
xor ( n50833 , n50831 , n50832 );
and ( n50834 , n20233 , n5103 );
xor ( n50835 , n50833 , n50834 );
xor ( n50836 , n50830 , n50835 );
and ( n50837 , n15758 , n6971 );
and ( n50838 , n16637 , n6504 );
xor ( n50839 , n50837 , n50838 );
and ( n50840 , n17512 , n6132 );
xor ( n50841 , n50839 , n50840 );
xor ( n50842 , n50836 , n50841 );
xor ( n50843 , n50826 , n50842 );
and ( n50844 , n49647 , n49648 );
and ( n50845 , n49648 , n49650 );
and ( n50846 , n49647 , n49650 );
or ( n50847 , n50844 , n50845 , n50846 );
and ( n50848 , n49678 , n49679 );
and ( n50849 , n49679 , n49681 );
and ( n50850 , n49678 , n49681 );
or ( n50851 , n50848 , n50849 , n50850 );
xor ( n50852 , n50847 , n50851 );
and ( n50853 , n13322 , n8243 );
and ( n50854 , n14118 , n7662 );
xor ( n50855 , n50853 , n50854 );
and ( n50856 , n14938 , n7310 );
xor ( n50857 , n50855 , n50856 );
xor ( n50858 , n50852 , n50857 );
xor ( n50859 , n50843 , n50858 );
xor ( n50860 , n50822 , n50859 );
xor ( n50861 , n50792 , n50860 );
and ( n50862 , n49668 , n49672 );
and ( n50863 , n49672 , n49689 );
and ( n50864 , n49668 , n49689 );
or ( n50865 , n50862 , n50863 , n50864 );
and ( n50866 , n49712 , n49727 );
and ( n50867 , n49727 , n49744 );
and ( n50868 , n49712 , n49744 );
or ( n50869 , n50866 , n50867 , n50868 );
xor ( n50870 , n50865 , n50869 );
and ( n50871 , n49677 , n49682 );
and ( n50872 , n49682 , n49688 );
and ( n50873 , n49677 , n49688 );
or ( n50874 , n50871 , n50872 , n50873 );
and ( n50875 , n49716 , n49720 );
and ( n50876 , n49720 , n49726 );
and ( n50877 , n49716 , n49726 );
or ( n50878 , n50875 , n50876 , n50877 );
xor ( n50879 , n50874 , n50878 );
and ( n50880 , n49684 , n49685 );
and ( n50881 , n49685 , n49687 );
and ( n50882 , n49684 , n49687 );
or ( n50883 , n50880 , n50881 , n50882 );
and ( n50884 , n11015 , n10239 );
and ( n50885 , n11769 , n9348 );
xor ( n50886 , n50884 , n50885 );
and ( n50887 , n12320 , n8669 );
xor ( n50888 , n50886 , n50887 );
xor ( n50889 , n50883 , n50888 );
and ( n50890 , n8718 , n12531 );
and ( n50891 , n9400 , n11718 );
xor ( n50892 , n50890 , n50891 );
and ( n50893 , n10291 , n10977 );
xor ( n50894 , n50892 , n50893 );
xor ( n50895 , n50889 , n50894 );
xor ( n50896 , n50879 , n50895 );
xor ( n50897 , n50870 , n50896 );
xor ( n50898 , n50861 , n50897 );
xor ( n50899 , n50788 , n50898 );
xor ( n50900 , n50779 , n50899 );
and ( n50901 , n49818 , n49823 );
and ( n50902 , n49778 , n49779 );
and ( n50903 , n49779 , n49817 );
and ( n50904 , n49778 , n49817 );
or ( n50905 , n50902 , n50903 , n50904 );
and ( n50906 , n49708 , n49745 );
and ( n50907 , n49745 , n49771 );
and ( n50908 , n49708 , n49771 );
or ( n50909 , n50906 , n50907 , n50908 );
xor ( n50910 , n50905 , n50909 );
and ( n50911 , n49750 , n49754 );
and ( n50912 , n49754 , n49770 );
and ( n50913 , n49750 , n49770 );
or ( n50914 , n50911 , n50912 , n50913 );
and ( n50915 , n49732 , n49737 );
and ( n50916 , n49737 , n49743 );
and ( n50917 , n49732 , n49743 );
or ( n50918 , n50915 , n50916 , n50917 );
and ( n50919 , n49722 , n49723 );
and ( n50920 , n49723 , n49725 );
and ( n50921 , n49722 , n49725 );
or ( n50922 , n50919 , n50920 , n50921 );
and ( n50923 , n49733 , n49734 );
and ( n50924 , n49734 , n49736 );
and ( n50925 , n49733 , n49736 );
or ( n50926 , n50923 , n50924 , n50925 );
xor ( n50927 , n50922 , n50926 );
and ( n50928 , n7385 , n14838 );
and ( n50929 , n7808 , n14044 );
xor ( n50930 , n50928 , n50929 );
and ( n50931 , n8079 , n13256 );
xor ( n50932 , n50930 , n50931 );
xor ( n50933 , n50927 , n50932 );
xor ( n50934 , n50918 , n50933 );
and ( n50935 , n49739 , n49740 );
and ( n50936 , n49740 , n49742 );
and ( n50937 , n49739 , n49742 );
or ( n50938 , n50935 , n50936 , n50937 );
and ( n50939 , n6187 , n17422 );
and ( n50940 , n6569 , n16550 );
xor ( n50941 , n50939 , n50940 );
and ( n50942 , n6816 , n15691 );
xor ( n50943 , n50941 , n50942 );
xor ( n50944 , n50938 , n50943 );
and ( n50945 , n4959 , n20156 );
and ( n50946 , n5459 , n19222 );
xor ( n50947 , n50945 , n50946 );
and ( n50948 , n5819 , n18407 );
xor ( n50949 , n50947 , n50948 );
xor ( n50950 , n50944 , n50949 );
xor ( n50951 , n50934 , n50950 );
xor ( n50952 , n50914 , n50951 );
and ( n50953 , n49759 , n49763 );
and ( n50954 , n49763 , n49769 );
and ( n50955 , n49759 , n49769 );
or ( n50956 , n50953 , n50954 , n50955 );
and ( n50957 , n49788 , n49793 );
and ( n50958 , n49793 , n49799 );
and ( n50959 , n49788 , n49799 );
or ( n50960 , n50957 , n50958 , n50959 );
xor ( n50961 , n50956 , n50960 );
and ( n50962 , n49765 , n49766 );
and ( n50963 , n49766 , n49768 );
and ( n50964 , n49765 , n49768 );
or ( n50965 , n50962 , n50963 , n50964 );
and ( n50966 , n49789 , n49790 );
and ( n50967 , n49790 , n49792 );
and ( n50968 , n49789 , n49792 );
or ( n50969 , n50966 , n50967 , n50968 );
xor ( n50970 , n50965 , n50969 );
and ( n50971 , n4132 , n23075 );
and ( n50972 , n4438 , n22065 );
xor ( n50973 , n50971 , n50972 );
and ( n50974 , n4766 , n20976 );
xor ( n50975 , n50973 , n50974 );
xor ( n50976 , n50970 , n50975 );
xor ( n50977 , n50961 , n50976 );
xor ( n50978 , n50952 , n50977 );
xor ( n50979 , n50910 , n50978 );
xor ( n50980 , n50901 , n50979 );
not ( n50981 , n1694 );
and ( n50982 , n34193 , n1694 );
nor ( n50983 , n50981 , n50982 );
and ( n50984 , n49784 , n49800 );
and ( n50985 , n49800 , n49816 );
and ( n50986 , n49784 , n49816 );
or ( n50987 , n50984 , n50985 , n50986 );
and ( n50988 , n49805 , n49809 );
and ( n50989 , n49809 , n49815 );
and ( n50990 , n49805 , n49815 );
or ( n50991 , n50988 , n50989 , n50990 );
and ( n50992 , n49795 , n49796 );
and ( n50993 , n49796 , n49798 );
and ( n50994 , n49795 , n49798 );
or ( n50995 , n50992 , n50993 , n50994 );
and ( n50996 , n3182 , n26216 );
and ( n50997 , n3545 , n25163 );
xor ( n50998 , n50996 , n50997 );
and ( n50999 , n3801 , n24137 );
xor ( n51000 , n50998 , n50999 );
xor ( n51001 , n50995 , n51000 );
and ( n51002 , n2462 , n29508 );
and ( n51003 , n2779 , n28406 );
xor ( n51004 , n51002 , n51003 );
and ( n51005 , n3024 , n27296 );
xor ( n51006 , n51004 , n51005 );
xor ( n51007 , n51001 , n51006 );
xor ( n51008 , n50991 , n51007 );
and ( n51009 , n49811 , n49812 );
and ( n51010 , n49812 , n49814 );
and ( n51011 , n49811 , n49814 );
or ( n51012 , n51009 , n51010 , n51011 );
and ( n51013 , n49821 , n49822 );
xor ( n51014 , n51012 , n51013 );
and ( n51015 , n1933 , n32999 );
and ( n51016 , n2120 , n31761 );
xor ( n51017 , n51015 , n51016 );
and ( n51018 , n2324 , n30629 );
xor ( n51019 , n51017 , n51018 );
xor ( n51020 , n51014 , n51019 );
xor ( n51021 , n51008 , n51020 );
xor ( n51022 , n50987 , n51021 );
xor ( n51023 , n50983 , n51022 );
xor ( n51024 , n50980 , n51023 );
xor ( n51025 , n50900 , n51024 );
xor ( n51026 , n50775 , n51025 );
xor ( n51027 , n50693 , n51026 );
xor ( n51028 , n50684 , n51027 );
and ( n51029 , n49474 , n49477 );
and ( n51030 , n49477 , n49828 );
and ( n51031 , n49474 , n49828 );
or ( n51032 , n51029 , n51030 , n51031 );
xor ( n51033 , n51028 , n51032 );
and ( n51034 , n49829 , n49833 );
and ( n51035 , n49834 , n49837 );
or ( n51036 , n51034 , n51035 );
xor ( n51037 , n51033 , n51036 );
buf ( n51038 , n51037 );
buf ( n51039 , n51038 );
not ( n51040 , n51039 );
nor ( n51041 , n51040 , n8739 );
xor ( n51042 , n50676 , n51041 );
and ( n51043 , n49470 , n49842 );
and ( n51044 , n49843 , n49846 );
or ( n51045 , n51043 , n51044 );
xor ( n51046 , n51042 , n51045 );
buf ( n51047 , n51046 );
buf ( n51048 , n51047 );
not ( n51049 , n51048 );
buf ( n51050 , n576 );
not ( n51051 , n51050 );
nor ( n51052 , n51049 , n51051 );
xor ( n51053 , n50302 , n51052 );
xor ( n51054 , n49858 , n50299 );
nor ( n51055 , n49850 , n51051 );
and ( n51056 , n51054 , n51055 );
xor ( n51057 , n51054 , n51055 );
xor ( n51058 , n49862 , n50297 );
nor ( n51059 , n48650 , n51051 );
and ( n51060 , n51058 , n51059 );
xor ( n51061 , n51058 , n51059 );
xor ( n51062 , n49866 , n50295 );
nor ( n51063 , n47449 , n51051 );
and ( n51064 , n51062 , n51063 );
xor ( n51065 , n51062 , n51063 );
xor ( n51066 , n49870 , n50293 );
nor ( n51067 , n46248 , n51051 );
and ( n51068 , n51066 , n51067 );
xor ( n51069 , n51066 , n51067 );
xor ( n51070 , n49874 , n50291 );
nor ( n51071 , n45047 , n51051 );
and ( n51072 , n51070 , n51071 );
xor ( n51073 , n51070 , n51071 );
xor ( n51074 , n49878 , n50289 );
nor ( n51075 , n43843 , n51051 );
and ( n51076 , n51074 , n51075 );
xor ( n51077 , n51074 , n51075 );
xor ( n51078 , n49882 , n50287 );
nor ( n51079 , n42641 , n51051 );
and ( n51080 , n51078 , n51079 );
xor ( n51081 , n51078 , n51079 );
xor ( n51082 , n49886 , n50285 );
nor ( n51083 , n41437 , n51051 );
and ( n51084 , n51082 , n51083 );
xor ( n51085 , n51082 , n51083 );
xor ( n51086 , n49890 , n50283 );
nor ( n51087 , n40232 , n51051 );
and ( n51088 , n51086 , n51087 );
xor ( n51089 , n51086 , n51087 );
xor ( n51090 , n49894 , n50281 );
nor ( n51091 , n39027 , n51051 );
and ( n51092 , n51090 , n51091 );
xor ( n51093 , n51090 , n51091 );
xor ( n51094 , n49898 , n50279 );
nor ( n51095 , n37825 , n51051 );
and ( n51096 , n51094 , n51095 );
xor ( n51097 , n51094 , n51095 );
xor ( n51098 , n49902 , n50277 );
nor ( n51099 , n36620 , n51051 );
and ( n51100 , n51098 , n51099 );
xor ( n51101 , n51098 , n51099 );
xor ( n51102 , n49906 , n50275 );
nor ( n51103 , n35419 , n51051 );
and ( n51104 , n51102 , n51103 );
xor ( n51105 , n51102 , n51103 );
xor ( n51106 , n49910 , n50273 );
nor ( n51107 , n34224 , n51051 );
and ( n51108 , n51106 , n51107 );
xor ( n51109 , n51106 , n51107 );
xor ( n51110 , n49914 , n50271 );
nor ( n51111 , n33033 , n51051 );
and ( n51112 , n51110 , n51111 );
xor ( n51113 , n51110 , n51111 );
xor ( n51114 , n49918 , n50269 );
nor ( n51115 , n31867 , n51051 );
and ( n51116 , n51114 , n51115 );
xor ( n51117 , n51114 , n51115 );
xor ( n51118 , n49922 , n50267 );
nor ( n51119 , n30725 , n51051 );
and ( n51120 , n51118 , n51119 );
xor ( n51121 , n51118 , n51119 );
xor ( n51122 , n49926 , n50265 );
nor ( n51123 , n29596 , n51051 );
and ( n51124 , n51122 , n51123 );
xor ( n51125 , n51122 , n51123 );
xor ( n51126 , n49930 , n50263 );
nor ( n51127 , n28487 , n51051 );
and ( n51128 , n51126 , n51127 );
xor ( n51129 , n51126 , n51127 );
xor ( n51130 , n49934 , n50261 );
nor ( n51131 , n27397 , n51051 );
and ( n51132 , n51130 , n51131 );
xor ( n51133 , n51130 , n51131 );
xor ( n51134 , n49938 , n50259 );
nor ( n51135 , n26326 , n51051 );
and ( n51136 , n51134 , n51135 );
xor ( n51137 , n51134 , n51135 );
xor ( n51138 , n49942 , n50257 );
nor ( n51139 , n25272 , n51051 );
and ( n51140 , n51138 , n51139 );
xor ( n51141 , n51138 , n51139 );
xor ( n51142 , n49946 , n50255 );
nor ( n51143 , n24242 , n51051 );
and ( n51144 , n51142 , n51143 );
xor ( n51145 , n51142 , n51143 );
xor ( n51146 , n49950 , n50253 );
nor ( n51147 , n23225 , n51051 );
and ( n51148 , n51146 , n51147 );
xor ( n51149 , n51146 , n51147 );
xor ( n51150 , n49954 , n50251 );
nor ( n51151 , n22231 , n51051 );
and ( n51152 , n51150 , n51151 );
xor ( n51153 , n51150 , n51151 );
xor ( n51154 , n49958 , n50249 );
nor ( n51155 , n21258 , n51051 );
and ( n51156 , n51154 , n51155 );
xor ( n51157 , n51154 , n51155 );
xor ( n51158 , n49962 , n50247 );
nor ( n51159 , n20303 , n51051 );
and ( n51160 , n51158 , n51159 );
xor ( n51161 , n51158 , n51159 );
xor ( n51162 , n49966 , n50245 );
nor ( n51163 , n19365 , n51051 );
and ( n51164 , n51162 , n51163 );
xor ( n51165 , n51162 , n51163 );
xor ( n51166 , n49970 , n50243 );
nor ( n51167 , n18448 , n51051 );
and ( n51168 , n51166 , n51167 );
xor ( n51169 , n51166 , n51167 );
xor ( n51170 , n49974 , n50241 );
nor ( n51171 , n17548 , n51051 );
and ( n51172 , n51170 , n51171 );
xor ( n51173 , n51170 , n51171 );
xor ( n51174 , n49978 , n50239 );
nor ( n51175 , n16669 , n51051 );
and ( n51176 , n51174 , n51175 );
xor ( n51177 , n51174 , n51175 );
xor ( n51178 , n49982 , n50237 );
nor ( n51179 , n15809 , n51051 );
and ( n51180 , n51178 , n51179 );
xor ( n51181 , n51178 , n51179 );
xor ( n51182 , n49986 , n50235 );
nor ( n51183 , n14968 , n51051 );
and ( n51184 , n51182 , n51183 );
xor ( n51185 , n51182 , n51183 );
xor ( n51186 , n49990 , n50233 );
nor ( n51187 , n14147 , n51051 );
and ( n51188 , n51186 , n51187 );
xor ( n51189 , n51186 , n51187 );
xor ( n51190 , n49994 , n50231 );
nor ( n51191 , n13349 , n51051 );
and ( n51192 , n51190 , n51191 );
xor ( n51193 , n51190 , n51191 );
xor ( n51194 , n49998 , n50229 );
nor ( n51195 , n12564 , n51051 );
and ( n51196 , n51194 , n51195 );
xor ( n51197 , n51194 , n51195 );
xor ( n51198 , n50002 , n50227 );
nor ( n51199 , n11799 , n51051 );
and ( n51200 , n51198 , n51199 );
xor ( n51201 , n51198 , n51199 );
xor ( n51202 , n50006 , n50225 );
nor ( n51203 , n11050 , n51051 );
and ( n51204 , n51202 , n51203 );
xor ( n51205 , n51202 , n51203 );
xor ( n51206 , n50010 , n50223 );
nor ( n51207 , n10321 , n51051 );
and ( n51208 , n51206 , n51207 );
xor ( n51209 , n51206 , n51207 );
xor ( n51210 , n50014 , n50221 );
nor ( n51211 , n9429 , n51051 );
and ( n51212 , n51210 , n51211 );
xor ( n51213 , n51210 , n51211 );
xor ( n51214 , n50018 , n50219 );
nor ( n51215 , n8949 , n51051 );
and ( n51216 , n51214 , n51215 );
xor ( n51217 , n51214 , n51215 );
xor ( n51218 , n50022 , n50217 );
nor ( n51219 , n9437 , n51051 );
and ( n51220 , n51218 , n51219 );
xor ( n51221 , n51218 , n51219 );
xor ( n51222 , n50026 , n50215 );
nor ( n51223 , n9446 , n51051 );
and ( n51224 , n51222 , n51223 );
xor ( n51225 , n51222 , n51223 );
xor ( n51226 , n50030 , n50213 );
nor ( n51227 , n9455 , n51051 );
and ( n51228 , n51226 , n51227 );
xor ( n51229 , n51226 , n51227 );
xor ( n51230 , n50034 , n50211 );
nor ( n51231 , n9464 , n51051 );
and ( n51232 , n51230 , n51231 );
xor ( n51233 , n51230 , n51231 );
xor ( n51234 , n50038 , n50209 );
nor ( n51235 , n9473 , n51051 );
and ( n51236 , n51234 , n51235 );
xor ( n51237 , n51234 , n51235 );
xor ( n51238 , n50042 , n50207 );
nor ( n51239 , n9482 , n51051 );
and ( n51240 , n51238 , n51239 );
xor ( n51241 , n51238 , n51239 );
xor ( n51242 , n50046 , n50205 );
nor ( n51243 , n9491 , n51051 );
and ( n51244 , n51242 , n51243 );
xor ( n51245 , n51242 , n51243 );
xor ( n51246 , n50050 , n50203 );
nor ( n51247 , n9500 , n51051 );
and ( n51248 , n51246 , n51247 );
xor ( n51249 , n51246 , n51247 );
xor ( n51250 , n50054 , n50201 );
nor ( n51251 , n9509 , n51051 );
and ( n51252 , n51250 , n51251 );
xor ( n51253 , n51250 , n51251 );
xor ( n51254 , n50058 , n50199 );
nor ( n51255 , n9518 , n51051 );
and ( n51256 , n51254 , n51255 );
xor ( n51257 , n51254 , n51255 );
xor ( n51258 , n50062 , n50197 );
nor ( n51259 , n9527 , n51051 );
and ( n51260 , n51258 , n51259 );
xor ( n51261 , n51258 , n51259 );
xor ( n51262 , n50066 , n50195 );
nor ( n51263 , n9536 , n51051 );
and ( n51264 , n51262 , n51263 );
xor ( n51265 , n51262 , n51263 );
xor ( n51266 , n50070 , n50193 );
nor ( n51267 , n9545 , n51051 );
and ( n51268 , n51266 , n51267 );
xor ( n51269 , n51266 , n51267 );
xor ( n51270 , n50074 , n50191 );
nor ( n51271 , n9554 , n51051 );
and ( n51272 , n51270 , n51271 );
xor ( n51273 , n51270 , n51271 );
xor ( n51274 , n50078 , n50189 );
nor ( n51275 , n9563 , n51051 );
and ( n51276 , n51274 , n51275 );
xor ( n51277 , n51274 , n51275 );
xor ( n51278 , n50082 , n50187 );
nor ( n51279 , n9572 , n51051 );
and ( n51280 , n51278 , n51279 );
xor ( n51281 , n51278 , n51279 );
xor ( n51282 , n50086 , n50185 );
nor ( n51283 , n9581 , n51051 );
and ( n51284 , n51282 , n51283 );
xor ( n51285 , n51282 , n51283 );
xor ( n51286 , n50090 , n50183 );
nor ( n51287 , n9590 , n51051 );
and ( n51288 , n51286 , n51287 );
xor ( n51289 , n51286 , n51287 );
xor ( n51290 , n50094 , n50181 );
nor ( n51291 , n9599 , n51051 );
and ( n51292 , n51290 , n51291 );
xor ( n51293 , n51290 , n51291 );
xor ( n51294 , n50098 , n50179 );
nor ( n51295 , n9608 , n51051 );
and ( n51296 , n51294 , n51295 );
xor ( n51297 , n51294 , n51295 );
xor ( n51298 , n50102 , n50177 );
nor ( n51299 , n9617 , n51051 );
and ( n51300 , n51298 , n51299 );
xor ( n51301 , n51298 , n51299 );
xor ( n51302 , n50106 , n50175 );
nor ( n51303 , n9626 , n51051 );
and ( n51304 , n51302 , n51303 );
xor ( n51305 , n51302 , n51303 );
xor ( n51306 , n50110 , n50173 );
nor ( n51307 , n9635 , n51051 );
and ( n51308 , n51306 , n51307 );
xor ( n51309 , n51306 , n51307 );
xor ( n51310 , n50114 , n50171 );
nor ( n51311 , n9644 , n51051 );
and ( n51312 , n51310 , n51311 );
xor ( n51313 , n51310 , n51311 );
xor ( n51314 , n50118 , n50169 );
nor ( n51315 , n9653 , n51051 );
and ( n51316 , n51314 , n51315 );
xor ( n51317 , n51314 , n51315 );
xor ( n51318 , n50122 , n50167 );
nor ( n51319 , n9662 , n51051 );
and ( n51320 , n51318 , n51319 );
xor ( n51321 , n51318 , n51319 );
xor ( n51322 , n50126 , n50165 );
nor ( n51323 , n9671 , n51051 );
and ( n51324 , n51322 , n51323 );
xor ( n51325 , n51322 , n51323 );
xor ( n51326 , n50130 , n50163 );
nor ( n51327 , n9680 , n51051 );
and ( n51328 , n51326 , n51327 );
xor ( n51329 , n51326 , n51327 );
xor ( n51330 , n50134 , n50161 );
nor ( n51331 , n9689 , n51051 );
and ( n51332 , n51330 , n51331 );
xor ( n51333 , n51330 , n51331 );
xor ( n51334 , n50138 , n50159 );
nor ( n51335 , n9698 , n51051 );
and ( n51336 , n51334 , n51335 );
xor ( n51337 , n51334 , n51335 );
xor ( n51338 , n50142 , n50157 );
nor ( n51339 , n9707 , n51051 );
and ( n51340 , n51338 , n51339 );
xor ( n51341 , n51338 , n51339 );
xor ( n51342 , n50146 , n50155 );
nor ( n51343 , n9716 , n51051 );
and ( n51344 , n51342 , n51343 );
xor ( n51345 , n51342 , n51343 );
xor ( n51346 , n50150 , n50153 );
nor ( n51347 , n9725 , n51051 );
and ( n51348 , n51346 , n51347 );
xor ( n51349 , n51346 , n51347 );
xor ( n51350 , n50151 , n50152 );
nor ( n51351 , n9734 , n51051 );
and ( n51352 , n51350 , n51351 );
xor ( n51353 , n51350 , n51351 );
nor ( n51354 , n9752 , n49852 );
nor ( n51355 , n9743 , n51051 );
and ( n51356 , n51354 , n51355 );
and ( n51357 , n51353 , n51356 );
or ( n51358 , n51352 , n51357 );
and ( n51359 , n51349 , n51358 );
or ( n51360 , n51348 , n51359 );
and ( n51361 , n51345 , n51360 );
or ( n51362 , n51344 , n51361 );
and ( n51363 , n51341 , n51362 );
or ( n51364 , n51340 , n51363 );
and ( n51365 , n51337 , n51364 );
or ( n51366 , n51336 , n51365 );
and ( n51367 , n51333 , n51366 );
or ( n51368 , n51332 , n51367 );
and ( n51369 , n51329 , n51368 );
or ( n51370 , n51328 , n51369 );
and ( n51371 , n51325 , n51370 );
or ( n51372 , n51324 , n51371 );
and ( n51373 , n51321 , n51372 );
or ( n51374 , n51320 , n51373 );
and ( n51375 , n51317 , n51374 );
or ( n51376 , n51316 , n51375 );
and ( n51377 , n51313 , n51376 );
or ( n51378 , n51312 , n51377 );
and ( n51379 , n51309 , n51378 );
or ( n51380 , n51308 , n51379 );
and ( n51381 , n51305 , n51380 );
or ( n51382 , n51304 , n51381 );
and ( n51383 , n51301 , n51382 );
or ( n51384 , n51300 , n51383 );
and ( n51385 , n51297 , n51384 );
or ( n51386 , n51296 , n51385 );
and ( n51387 , n51293 , n51386 );
or ( n51388 , n51292 , n51387 );
and ( n51389 , n51289 , n51388 );
or ( n51390 , n51288 , n51389 );
and ( n51391 , n51285 , n51390 );
or ( n51392 , n51284 , n51391 );
and ( n51393 , n51281 , n51392 );
or ( n51394 , n51280 , n51393 );
and ( n51395 , n51277 , n51394 );
or ( n51396 , n51276 , n51395 );
and ( n51397 , n51273 , n51396 );
or ( n51398 , n51272 , n51397 );
and ( n51399 , n51269 , n51398 );
or ( n51400 , n51268 , n51399 );
and ( n51401 , n51265 , n51400 );
or ( n51402 , n51264 , n51401 );
and ( n51403 , n51261 , n51402 );
or ( n51404 , n51260 , n51403 );
and ( n51405 , n51257 , n51404 );
or ( n51406 , n51256 , n51405 );
and ( n51407 , n51253 , n51406 );
or ( n51408 , n51252 , n51407 );
and ( n51409 , n51249 , n51408 );
or ( n51410 , n51248 , n51409 );
and ( n51411 , n51245 , n51410 );
or ( n51412 , n51244 , n51411 );
and ( n51413 , n51241 , n51412 );
or ( n51414 , n51240 , n51413 );
and ( n51415 , n51237 , n51414 );
or ( n51416 , n51236 , n51415 );
and ( n51417 , n51233 , n51416 );
or ( n51418 , n51232 , n51417 );
and ( n51419 , n51229 , n51418 );
or ( n51420 , n51228 , n51419 );
and ( n51421 , n51225 , n51420 );
or ( n51422 , n51224 , n51421 );
and ( n51423 , n51221 , n51422 );
or ( n51424 , n51220 , n51423 );
and ( n51425 , n51217 , n51424 );
or ( n51426 , n51216 , n51425 );
and ( n51427 , n51213 , n51426 );
or ( n51428 , n51212 , n51427 );
and ( n51429 , n51209 , n51428 );
or ( n51430 , n51208 , n51429 );
and ( n51431 , n51205 , n51430 );
or ( n51432 , n51204 , n51431 );
and ( n51433 , n51201 , n51432 );
or ( n51434 , n51200 , n51433 );
and ( n51435 , n51197 , n51434 );
or ( n51436 , n51196 , n51435 );
and ( n51437 , n51193 , n51436 );
or ( n51438 , n51192 , n51437 );
and ( n51439 , n51189 , n51438 );
or ( n51440 , n51188 , n51439 );
and ( n51441 , n51185 , n51440 );
or ( n51442 , n51184 , n51441 );
and ( n51443 , n51181 , n51442 );
or ( n51444 , n51180 , n51443 );
and ( n51445 , n51177 , n51444 );
or ( n51446 , n51176 , n51445 );
and ( n51447 , n51173 , n51446 );
or ( n51448 , n51172 , n51447 );
and ( n51449 , n51169 , n51448 );
or ( n51450 , n51168 , n51449 );
and ( n51451 , n51165 , n51450 );
or ( n51452 , n51164 , n51451 );
and ( n51453 , n51161 , n51452 );
or ( n51454 , n51160 , n51453 );
and ( n51455 , n51157 , n51454 );
or ( n51456 , n51156 , n51455 );
and ( n51457 , n51153 , n51456 );
or ( n51458 , n51152 , n51457 );
and ( n51459 , n51149 , n51458 );
or ( n51460 , n51148 , n51459 );
and ( n51461 , n51145 , n51460 );
or ( n51462 , n51144 , n51461 );
and ( n51463 , n51141 , n51462 );
or ( n51464 , n51140 , n51463 );
and ( n51465 , n51137 , n51464 );
or ( n51466 , n51136 , n51465 );
and ( n51467 , n51133 , n51466 );
or ( n51468 , n51132 , n51467 );
and ( n51469 , n51129 , n51468 );
or ( n51470 , n51128 , n51469 );
and ( n51471 , n51125 , n51470 );
or ( n51472 , n51124 , n51471 );
and ( n51473 , n51121 , n51472 );
or ( n51474 , n51120 , n51473 );
and ( n51475 , n51117 , n51474 );
or ( n51476 , n51116 , n51475 );
and ( n51477 , n51113 , n51476 );
or ( n51478 , n51112 , n51477 );
and ( n51479 , n51109 , n51478 );
or ( n51480 , n51108 , n51479 );
and ( n51481 , n51105 , n51480 );
or ( n51482 , n51104 , n51481 );
and ( n51483 , n51101 , n51482 );
or ( n51484 , n51100 , n51483 );
and ( n51485 , n51097 , n51484 );
or ( n51486 , n51096 , n51485 );
and ( n51487 , n51093 , n51486 );
or ( n51488 , n51092 , n51487 );
and ( n51489 , n51089 , n51488 );
or ( n51490 , n51088 , n51489 );
and ( n51491 , n51085 , n51490 );
or ( n51492 , n51084 , n51491 );
and ( n51493 , n51081 , n51492 );
or ( n51494 , n51080 , n51493 );
and ( n51495 , n51077 , n51494 );
or ( n51496 , n51076 , n51495 );
and ( n51497 , n51073 , n51496 );
or ( n51498 , n51072 , n51497 );
and ( n51499 , n51069 , n51498 );
or ( n51500 , n51068 , n51499 );
and ( n51501 , n51065 , n51500 );
or ( n51502 , n51064 , n51501 );
and ( n51503 , n51061 , n51502 );
or ( n51504 , n51060 , n51503 );
and ( n51505 , n51057 , n51504 );
or ( n51506 , n51056 , n51505 );
xor ( n51507 , n51053 , n51506 );
and ( n51508 , n33403 , n1944 );
nor ( n51509 , n1945 , n51508 );
nor ( n51510 , n2137 , n32231 );
xor ( n51511 , n51509 , n51510 );
and ( n51512 , n50304 , n50305 );
and ( n51513 , n50306 , n50309 );
or ( n51514 , n51512 , n51513 );
xor ( n51515 , n51511 , n51514 );
nor ( n51516 , n2343 , n31083 );
xor ( n51517 , n51515 , n51516 );
and ( n51518 , n50310 , n50311 );
and ( n51519 , n50312 , n50315 );
or ( n51520 , n51518 , n51519 );
xor ( n51521 , n51517 , n51520 );
nor ( n51522 , n2566 , n29948 );
xor ( n51523 , n51521 , n51522 );
and ( n51524 , n50316 , n50317 );
and ( n51525 , n50318 , n50321 );
or ( n51526 , n51524 , n51525 );
xor ( n51527 , n51523 , n51526 );
nor ( n51528 , n2797 , n28833 );
xor ( n51529 , n51527 , n51528 );
and ( n51530 , n50322 , n50323 );
and ( n51531 , n50324 , n50327 );
or ( n51532 , n51530 , n51531 );
xor ( n51533 , n51529 , n51532 );
nor ( n51534 , n3043 , n27737 );
xor ( n51535 , n51533 , n51534 );
and ( n51536 , n50328 , n50329 );
and ( n51537 , n50330 , n50333 );
or ( n51538 , n51536 , n51537 );
xor ( n51539 , n51535 , n51538 );
nor ( n51540 , n3300 , n26660 );
xor ( n51541 , n51539 , n51540 );
and ( n51542 , n50334 , n50335 );
and ( n51543 , n50336 , n50339 );
or ( n51544 , n51542 , n51543 );
xor ( n51545 , n51541 , n51544 );
nor ( n51546 , n3570 , n25600 );
xor ( n51547 , n51545 , n51546 );
and ( n51548 , n50340 , n50341 );
and ( n51549 , n50342 , n50345 );
or ( n51550 , n51548 , n51549 );
xor ( n51551 , n51547 , n51550 );
nor ( n51552 , n3853 , n24564 );
xor ( n51553 , n51551 , n51552 );
and ( n51554 , n50346 , n50347 );
and ( n51555 , n50348 , n50351 );
or ( n51556 , n51554 , n51555 );
xor ( n51557 , n51553 , n51556 );
nor ( n51558 , n4151 , n23541 );
xor ( n51559 , n51557 , n51558 );
and ( n51560 , n50352 , n50353 );
and ( n51561 , n50354 , n50357 );
or ( n51562 , n51560 , n51561 );
xor ( n51563 , n51559 , n51562 );
nor ( n51564 , n4458 , n22541 );
xor ( n51565 , n51563 , n51564 );
and ( n51566 , n50358 , n50359 );
and ( n51567 , n50360 , n50363 );
or ( n51568 , n51566 , n51567 );
xor ( n51569 , n51565 , n51568 );
nor ( n51570 , n4786 , n21562 );
xor ( n51571 , n51569 , n51570 );
and ( n51572 , n50364 , n50365 );
and ( n51573 , n50366 , n50369 );
or ( n51574 , n51572 , n51573 );
xor ( n51575 , n51571 , n51574 );
nor ( n51576 , n5126 , n20601 );
xor ( n51577 , n51575 , n51576 );
and ( n51578 , n50370 , n50371 );
and ( n51579 , n50372 , n50375 );
or ( n51580 , n51578 , n51579 );
xor ( n51581 , n51577 , n51580 );
nor ( n51582 , n5477 , n19657 );
xor ( n51583 , n51581 , n51582 );
and ( n51584 , n50376 , n50377 );
and ( n51585 , n50378 , n50381 );
or ( n51586 , n51584 , n51585 );
xor ( n51587 , n51583 , n51586 );
nor ( n51588 , n5838 , n18734 );
xor ( n51589 , n51587 , n51588 );
and ( n51590 , n50382 , n50383 );
and ( n51591 , n50384 , n50387 );
or ( n51592 , n51590 , n51591 );
xor ( n51593 , n51589 , n51592 );
nor ( n51594 , n6212 , n17828 );
xor ( n51595 , n51593 , n51594 );
and ( n51596 , n50388 , n50389 );
and ( n51597 , n50390 , n50393 );
or ( n51598 , n51596 , n51597 );
xor ( n51599 , n51595 , n51598 );
nor ( n51600 , n6596 , n16943 );
xor ( n51601 , n51599 , n51600 );
and ( n51602 , n50394 , n50395 );
and ( n51603 , n50396 , n50399 );
or ( n51604 , n51602 , n51603 );
xor ( n51605 , n51601 , n51604 );
nor ( n51606 , n6997 , n16077 );
xor ( n51607 , n51605 , n51606 );
and ( n51608 , n50400 , n50401 );
and ( n51609 , n50402 , n50405 );
or ( n51610 , n51608 , n51609 );
xor ( n51611 , n51607 , n51610 );
nor ( n51612 , n7413 , n15230 );
xor ( n51613 , n51611 , n51612 );
and ( n51614 , n50406 , n50407 );
and ( n51615 , n50408 , n50411 );
or ( n51616 , n51614 , n51615 );
xor ( n51617 , n51613 , n51616 );
nor ( n51618 , n7841 , n14403 );
xor ( n51619 , n51617 , n51618 );
and ( n51620 , n50412 , n50413 );
and ( n51621 , n50414 , n50417 );
or ( n51622 , n51620 , n51621 );
xor ( n51623 , n51619 , n51622 );
nor ( n51624 , n8281 , n13599 );
xor ( n51625 , n51623 , n51624 );
and ( n51626 , n50418 , n50419 );
and ( n51627 , n50420 , n50423 );
or ( n51628 , n51626 , n51627 );
xor ( n51629 , n51625 , n51628 );
nor ( n51630 , n8737 , n12808 );
xor ( n51631 , n51629 , n51630 );
and ( n51632 , n50424 , n50425 );
and ( n51633 , n50426 , n50429 );
or ( n51634 , n51632 , n51633 );
xor ( n51635 , n51631 , n51634 );
nor ( n51636 , n9420 , n12037 );
xor ( n51637 , n51635 , n51636 );
and ( n51638 , n50430 , n50431 );
and ( n51639 , n50432 , n50435 );
or ( n51640 , n51638 , n51639 );
xor ( n51641 , n51637 , n51640 );
nor ( n51642 , n10312 , n11282 );
xor ( n51643 , n51641 , n51642 );
and ( n51644 , n50436 , n50437 );
and ( n51645 , n50438 , n50441 );
or ( n51646 , n51644 , n51645 );
xor ( n51647 , n51643 , n51646 );
nor ( n51648 , n11041 , n10547 );
xor ( n51649 , n51647 , n51648 );
and ( n51650 , n50442 , n50443 );
and ( n51651 , n50444 , n50447 );
or ( n51652 , n51650 , n51651 );
xor ( n51653 , n51649 , n51652 );
nor ( n51654 , n11790 , n9829 );
xor ( n51655 , n51653 , n51654 );
and ( n51656 , n50448 , n50449 );
and ( n51657 , n50450 , n50453 );
or ( n51658 , n51656 , n51657 );
xor ( n51659 , n51655 , n51658 );
nor ( n51660 , n12555 , n8955 );
xor ( n51661 , n51659 , n51660 );
and ( n51662 , n50454 , n50455 );
and ( n51663 , n50456 , n50459 );
or ( n51664 , n51662 , n51663 );
xor ( n51665 , n51661 , n51664 );
nor ( n51666 , n13340 , n603 );
xor ( n51667 , n51665 , n51666 );
and ( n51668 , n50460 , n50461 );
and ( n51669 , n50462 , n50465 );
or ( n51670 , n51668 , n51669 );
xor ( n51671 , n51667 , n51670 );
nor ( n51672 , n14138 , n652 );
xor ( n51673 , n51671 , n51672 );
and ( n51674 , n50466 , n50467 );
and ( n51675 , n50468 , n50471 );
or ( n51676 , n51674 , n51675 );
xor ( n51677 , n51673 , n51676 );
nor ( n51678 , n14959 , n624 );
xor ( n51679 , n51677 , n51678 );
and ( n51680 , n50472 , n50473 );
and ( n51681 , n50474 , n50477 );
or ( n51682 , n51680 , n51681 );
xor ( n51683 , n51679 , n51682 );
nor ( n51684 , n15800 , n648 );
xor ( n51685 , n51683 , n51684 );
and ( n51686 , n50478 , n50479 );
and ( n51687 , n50480 , n50483 );
or ( n51688 , n51686 , n51687 );
xor ( n51689 , n51685 , n51688 );
nor ( n51690 , n16660 , n686 );
xor ( n51691 , n51689 , n51690 );
and ( n51692 , n50484 , n50485 );
and ( n51693 , n50486 , n50489 );
or ( n51694 , n51692 , n51693 );
xor ( n51695 , n51691 , n51694 );
nor ( n51696 , n17539 , n735 );
xor ( n51697 , n51695 , n51696 );
and ( n51698 , n50490 , n50491 );
and ( n51699 , n50492 , n50495 );
or ( n51700 , n51698 , n51699 );
xor ( n51701 , n51697 , n51700 );
nor ( n51702 , n18439 , n798 );
xor ( n51703 , n51701 , n51702 );
and ( n51704 , n50496 , n50497 );
and ( n51705 , n50498 , n50501 );
or ( n51706 , n51704 , n51705 );
xor ( n51707 , n51703 , n51706 );
nor ( n51708 , n19356 , n870 );
xor ( n51709 , n51707 , n51708 );
and ( n51710 , n50502 , n50503 );
and ( n51711 , n50504 , n50507 );
or ( n51712 , n51710 , n51711 );
xor ( n51713 , n51709 , n51712 );
nor ( n51714 , n20294 , n960 );
xor ( n51715 , n51713 , n51714 );
and ( n51716 , n50508 , n50509 );
and ( n51717 , n50510 , n50513 );
or ( n51718 , n51716 , n51717 );
xor ( n51719 , n51715 , n51718 );
nor ( n51720 , n21249 , n1064 );
xor ( n51721 , n51719 , n51720 );
and ( n51722 , n50514 , n50515 );
and ( n51723 , n50516 , n50519 );
or ( n51724 , n51722 , n51723 );
xor ( n51725 , n51721 , n51724 );
nor ( n51726 , n22222 , n1178 );
xor ( n51727 , n51725 , n51726 );
and ( n51728 , n50520 , n50521 );
and ( n51729 , n50522 , n50525 );
or ( n51730 , n51728 , n51729 );
xor ( n51731 , n51727 , n51730 );
nor ( n51732 , n23216 , n1305 );
xor ( n51733 , n51731 , n51732 );
and ( n51734 , n50526 , n50527 );
and ( n51735 , n50528 , n50531 );
or ( n51736 , n51734 , n51735 );
xor ( n51737 , n51733 , n51736 );
nor ( n51738 , n24233 , n1447 );
xor ( n51739 , n51737 , n51738 );
and ( n51740 , n50532 , n50533 );
and ( n51741 , n50534 , n50537 );
or ( n51742 , n51740 , n51741 );
xor ( n51743 , n51739 , n51742 );
nor ( n51744 , n25263 , n1600 );
xor ( n51745 , n51743 , n51744 );
and ( n51746 , n50538 , n50539 );
and ( n51747 , n50540 , n50543 );
or ( n51748 , n51746 , n51747 );
xor ( n51749 , n51745 , n51748 );
nor ( n51750 , n26317 , n1768 );
xor ( n51751 , n51749 , n51750 );
and ( n51752 , n50544 , n50545 );
and ( n51753 , n50546 , n50549 );
or ( n51754 , n51752 , n51753 );
xor ( n51755 , n51751 , n51754 );
nor ( n51756 , n27388 , n1947 );
xor ( n51757 , n51755 , n51756 );
and ( n51758 , n50550 , n50551 );
and ( n51759 , n50552 , n50555 );
or ( n51760 , n51758 , n51759 );
xor ( n51761 , n51757 , n51760 );
nor ( n51762 , n28478 , n2139 );
xor ( n51763 , n51761 , n51762 );
and ( n51764 , n50556 , n50557 );
and ( n51765 , n50558 , n50561 );
or ( n51766 , n51764 , n51765 );
xor ( n51767 , n51763 , n51766 );
nor ( n51768 , n29587 , n2345 );
xor ( n51769 , n51767 , n51768 );
and ( n51770 , n50562 , n50563 );
and ( n51771 , n50564 , n50567 );
or ( n51772 , n51770 , n51771 );
xor ( n51773 , n51769 , n51772 );
nor ( n51774 , n30716 , n2568 );
xor ( n51775 , n51773 , n51774 );
and ( n51776 , n50568 , n50569 );
and ( n51777 , n50570 , n50573 );
or ( n51778 , n51776 , n51777 );
xor ( n51779 , n51775 , n51778 );
nor ( n51780 , n31858 , n2799 );
xor ( n51781 , n51779 , n51780 );
and ( n51782 , n50574 , n50575 );
and ( n51783 , n50576 , n50579 );
or ( n51784 , n51782 , n51783 );
xor ( n51785 , n51781 , n51784 );
nor ( n51786 , n33024 , n3045 );
xor ( n51787 , n51785 , n51786 );
and ( n51788 , n50580 , n50581 );
and ( n51789 , n50582 , n50585 );
or ( n51790 , n51788 , n51789 );
xor ( n51791 , n51787 , n51790 );
nor ( n51792 , n34215 , n3302 );
xor ( n51793 , n51791 , n51792 );
and ( n51794 , n50586 , n50587 );
and ( n51795 , n50588 , n50591 );
or ( n51796 , n51794 , n51795 );
xor ( n51797 , n51793 , n51796 );
nor ( n51798 , n35410 , n3572 );
xor ( n51799 , n51797 , n51798 );
and ( n51800 , n50592 , n50593 );
and ( n51801 , n50594 , n50597 );
or ( n51802 , n51800 , n51801 );
xor ( n51803 , n51799 , n51802 );
nor ( n51804 , n36611 , n3855 );
xor ( n51805 , n51803 , n51804 );
and ( n51806 , n50598 , n50599 );
and ( n51807 , n50600 , n50603 );
or ( n51808 , n51806 , n51807 );
xor ( n51809 , n51805 , n51808 );
nor ( n51810 , n37816 , n4153 );
xor ( n51811 , n51809 , n51810 );
and ( n51812 , n50604 , n50605 );
and ( n51813 , n50606 , n50609 );
or ( n51814 , n51812 , n51813 );
xor ( n51815 , n51811 , n51814 );
nor ( n51816 , n39018 , n4460 );
xor ( n51817 , n51815 , n51816 );
and ( n51818 , n50610 , n50611 );
and ( n51819 , n50612 , n50615 );
or ( n51820 , n51818 , n51819 );
xor ( n51821 , n51817 , n51820 );
nor ( n51822 , n40223 , n4788 );
xor ( n51823 , n51821 , n51822 );
and ( n51824 , n50616 , n50617 );
and ( n51825 , n50618 , n50621 );
or ( n51826 , n51824 , n51825 );
xor ( n51827 , n51823 , n51826 );
nor ( n51828 , n41428 , n5128 );
xor ( n51829 , n51827 , n51828 );
and ( n51830 , n50622 , n50623 );
and ( n51831 , n50624 , n50627 );
or ( n51832 , n51830 , n51831 );
xor ( n51833 , n51829 , n51832 );
nor ( n51834 , n42632 , n5479 );
xor ( n51835 , n51833 , n51834 );
and ( n51836 , n50628 , n50629 );
and ( n51837 , n50630 , n50633 );
or ( n51838 , n51836 , n51837 );
xor ( n51839 , n51835 , n51838 );
nor ( n51840 , n43834 , n5840 );
xor ( n51841 , n51839 , n51840 );
and ( n51842 , n50634 , n50635 );
and ( n51843 , n50636 , n50639 );
or ( n51844 , n51842 , n51843 );
xor ( n51845 , n51841 , n51844 );
nor ( n51846 , n45038 , n6214 );
xor ( n51847 , n51845 , n51846 );
and ( n51848 , n50640 , n50641 );
and ( n51849 , n50642 , n50645 );
or ( n51850 , n51848 , n51849 );
xor ( n51851 , n51847 , n51850 );
nor ( n51852 , n46239 , n6598 );
xor ( n51853 , n51851 , n51852 );
and ( n51854 , n50646 , n50647 );
and ( n51855 , n50648 , n50651 );
or ( n51856 , n51854 , n51855 );
xor ( n51857 , n51853 , n51856 );
nor ( n51858 , n47440 , n6999 );
xor ( n51859 , n51857 , n51858 );
and ( n51860 , n50652 , n50653 );
and ( n51861 , n50654 , n50657 );
or ( n51862 , n51860 , n51861 );
xor ( n51863 , n51859 , n51862 );
nor ( n51864 , n48641 , n7415 );
xor ( n51865 , n51863 , n51864 );
and ( n51866 , n50658 , n50659 );
and ( n51867 , n50660 , n50663 );
or ( n51868 , n51866 , n51867 );
xor ( n51869 , n51865 , n51868 );
nor ( n51870 , n49841 , n7843 );
xor ( n51871 , n51869 , n51870 );
and ( n51872 , n50664 , n50665 );
and ( n51873 , n50666 , n50669 );
or ( n51874 , n51872 , n51873 );
xor ( n51875 , n51871 , n51874 );
nor ( n51876 , n51040 , n8283 );
xor ( n51877 , n51875 , n51876 );
and ( n51878 , n50670 , n50671 );
and ( n51879 , n50672 , n50675 );
or ( n51880 , n51878 , n51879 );
xor ( n51881 , n51877 , n51880 );
and ( n51882 , n50688 , n50692 );
and ( n51883 , n50692 , n51026 );
and ( n51884 , n50688 , n51026 );
or ( n51885 , n51882 , n51883 , n51884 );
and ( n51886 , n33774 , n1882 );
not ( n51887 , n1882 );
nor ( n51888 , n51886 , n51887 );
xor ( n51889 , n51885 , n51888 );
and ( n51890 , n50701 , n50705 );
and ( n51891 , n50705 , n50773 );
and ( n51892 , n50701 , n50773 );
or ( n51893 , n51890 , n51891 , n51892 );
and ( n51894 , n50697 , n50774 );
and ( n51895 , n50774 , n51025 );
and ( n51896 , n50697 , n51025 );
or ( n51897 , n51894 , n51895 , n51896 );
xor ( n51898 , n51893 , n51897 );
and ( n51899 , n50779 , n50899 );
and ( n51900 , n50899 , n51024 );
and ( n51901 , n50779 , n51024 );
or ( n51902 , n51899 , n51900 , n51901 );
and ( n51903 , n50710 , n50714 );
and ( n51904 , n50714 , n50772 );
and ( n51905 , n50710 , n50772 );
or ( n51906 , n51903 , n51904 , n51905 );
and ( n51907 , n50783 , n50787 );
and ( n51908 , n50787 , n50898 );
and ( n51909 , n50783 , n50898 );
or ( n51910 , n51907 , n51908 , n51909 );
xor ( n51911 , n51906 , n51910 );
and ( n51912 , n50741 , n50745 );
and ( n51913 , n50745 , n50751 );
and ( n51914 , n50741 , n50751 );
or ( n51915 , n51912 , n51913 , n51914 );
and ( n51916 , n50719 , n50723 );
and ( n51917 , n50723 , n50771 );
and ( n51918 , n50719 , n50771 );
or ( n51919 , n51916 , n51917 , n51918 );
xor ( n51920 , n51915 , n51919 );
and ( n51921 , n50728 , n50732 );
and ( n51922 , n50732 , n50770 );
and ( n51923 , n50728 , n50770 );
or ( n51924 , n51921 , n51922 , n51923 );
and ( n51925 , n50796 , n50821 );
and ( n51926 , n50821 , n50859 );
and ( n51927 , n50796 , n50859 );
or ( n51928 , n51925 , n51926 , n51927 );
xor ( n51929 , n51924 , n51928 );
and ( n51930 , n50737 , n50752 );
and ( n51931 , n50752 , n50769 );
and ( n51932 , n50737 , n50769 );
or ( n51933 , n51930 , n51931 , n51932 );
and ( n51934 , n50800 , n50804 );
and ( n51935 , n50804 , n50820 );
and ( n51936 , n50800 , n50820 );
or ( n51937 , n51934 , n51935 , n51936 );
xor ( n51938 , n51933 , n51937 );
and ( n51939 , n50757 , n50762 );
and ( n51940 , n50762 , n50768 );
and ( n51941 , n50757 , n50768 );
or ( n51942 , n51939 , n51940 , n51941 );
and ( n51943 , n50747 , n50748 );
and ( n51944 , n50748 , n50750 );
and ( n51945 , n50747 , n50750 );
or ( n51946 , n51943 , n51944 , n51945 );
and ( n51947 , n50758 , n50759 );
and ( n51948 , n50759 , n50761 );
and ( n51949 , n50758 , n50761 );
or ( n51950 , n51947 , n51948 , n51949 );
xor ( n51951 , n51946 , n51950 );
and ( n51952 , n30695 , n2544 );
and ( n51953 , n31836 , n2298 );
xor ( n51954 , n51952 , n51953 );
and ( n51955 , n32649 , n2100 );
xor ( n51956 , n51954 , n51955 );
xor ( n51957 , n51951 , n51956 );
xor ( n51958 , n51942 , n51957 );
and ( n51959 , n50764 , n50765 );
and ( n51960 , n50765 , n50767 );
and ( n51961 , n50764 , n50767 );
or ( n51962 , n51959 , n51960 , n51961 );
and ( n51963 , n27361 , n3271 );
and ( n51964 , n28456 , n2981 );
xor ( n51965 , n51963 , n51964 );
and ( n51966 , n29559 , n2739 );
xor ( n51967 , n51965 , n51966 );
xor ( n51968 , n51962 , n51967 );
and ( n51969 , n24214 , n4102 );
and ( n51970 , n25243 , n3749 );
xor ( n51971 , n51969 , n51970 );
and ( n51972 , n26296 , n3495 );
xor ( n51973 , n51971 , n51972 );
xor ( n51974 , n51968 , n51973 );
xor ( n51975 , n51958 , n51974 );
xor ( n51976 , n51938 , n51975 );
xor ( n51977 , n51929 , n51976 );
xor ( n51978 , n51920 , n51977 );
xor ( n51979 , n51911 , n51978 );
xor ( n51980 , n51902 , n51979 );
and ( n51981 , n50901 , n50979 );
and ( n51982 , n50979 , n51023 );
and ( n51983 , n50901 , n51023 );
or ( n51984 , n51981 , n51982 , n51983 );
and ( n51985 , n50792 , n50860 );
and ( n51986 , n50860 , n50897 );
and ( n51987 , n50792 , n50897 );
or ( n51988 , n51985 , n51986 , n51987 );
and ( n51989 , n50905 , n50909 );
and ( n51990 , n50909 , n50978 );
and ( n51991 , n50905 , n50978 );
or ( n51992 , n51989 , n51990 , n51991 );
xor ( n51993 , n51988 , n51992 );
and ( n51994 , n50865 , n50869 );
and ( n51995 , n50869 , n50896 );
and ( n51996 , n50865 , n50896 );
or ( n51997 , n51994 , n51995 , n51996 );
and ( n51998 , n50826 , n50842 );
and ( n51999 , n50842 , n50858 );
and ( n52000 , n50826 , n50858 );
or ( n52001 , n51998 , n51999 , n52000 );
and ( n52002 , n50809 , n50813 );
and ( n52003 , n50813 , n50819 );
and ( n52004 , n50809 , n50819 );
or ( n52005 , n52002 , n52003 , n52004 );
and ( n52006 , n50830 , n50835 );
and ( n52007 , n50835 , n50841 );
and ( n52008 , n50830 , n50841 );
or ( n52009 , n52006 , n52007 , n52008 );
xor ( n52010 , n52005 , n52009 );
and ( n52011 , n50815 , n50816 );
and ( n52012 , n50816 , n50818 );
and ( n52013 , n50815 , n50818 );
or ( n52014 , n52011 , n52012 , n52013 );
and ( n52015 , n50831 , n50832 );
and ( n52016 , n50832 , n50834 );
and ( n52017 , n50831 , n50834 );
or ( n52018 , n52015 , n52016 , n52017 );
xor ( n52019 , n52014 , n52018 );
and ( n52020 , n21216 , n5103 );
and ( n52021 , n22186 , n4730 );
xor ( n52022 , n52020 , n52021 );
and ( n52023 , n22892 , n4403 );
xor ( n52024 , n52022 , n52023 );
xor ( n52025 , n52019 , n52024 );
xor ( n52026 , n52010 , n52025 );
xor ( n52027 , n52001 , n52026 );
and ( n52028 , n50847 , n50851 );
and ( n52029 , n50851 , n50857 );
and ( n52030 , n50847 , n50857 );
or ( n52031 , n52028 , n52029 , n52030 );
and ( n52032 , n50837 , n50838 );
and ( n52033 , n50838 , n50840 );
and ( n52034 , n50837 , n50840 );
or ( n52035 , n52032 , n52033 , n52034 );
and ( n52036 , n18144 , n6132 );
and ( n52037 , n19324 , n5765 );
xor ( n52038 , n52036 , n52037 );
and ( n52039 , n20233 , n5408 );
xor ( n52040 , n52038 , n52039 );
xor ( n52041 , n52035 , n52040 );
and ( n52042 , n15758 , n7310 );
and ( n52043 , n16637 , n6971 );
xor ( n52044 , n52042 , n52043 );
and ( n52045 , n17512 , n6504 );
xor ( n52046 , n52044 , n52045 );
xor ( n52047 , n52041 , n52046 );
xor ( n52048 , n52031 , n52047 );
and ( n52049 , n50853 , n50854 );
and ( n52050 , n50854 , n50856 );
and ( n52051 , n50853 , n50856 );
or ( n52052 , n52049 , n52050 , n52051 );
and ( n52053 , n50884 , n50885 );
and ( n52054 , n50885 , n50887 );
and ( n52055 , n50884 , n50887 );
or ( n52056 , n52053 , n52054 , n52055 );
xor ( n52057 , n52052 , n52056 );
and ( n52058 , n13322 , n8669 );
and ( n52059 , n14118 , n8243 );
xor ( n52060 , n52058 , n52059 );
and ( n52061 , n14938 , n7662 );
xor ( n52062 , n52060 , n52061 );
xor ( n52063 , n52057 , n52062 );
xor ( n52064 , n52048 , n52063 );
xor ( n52065 , n52027 , n52064 );
xor ( n52066 , n51997 , n52065 );
and ( n52067 , n50874 , n50878 );
and ( n52068 , n50878 , n50895 );
and ( n52069 , n50874 , n50895 );
or ( n52070 , n52067 , n52068 , n52069 );
and ( n52071 , n50918 , n50933 );
and ( n52072 , n50933 , n50950 );
and ( n52073 , n50918 , n50950 );
or ( n52074 , n52071 , n52072 , n52073 );
xor ( n52075 , n52070 , n52074 );
and ( n52076 , n50883 , n50888 );
and ( n52077 , n50888 , n50894 );
and ( n52078 , n50883 , n50894 );
or ( n52079 , n52076 , n52077 , n52078 );
and ( n52080 , n50922 , n50926 );
and ( n52081 , n50926 , n50932 );
and ( n52082 , n50922 , n50932 );
or ( n52083 , n52080 , n52081 , n52082 );
xor ( n52084 , n52079 , n52083 );
and ( n52085 , n50890 , n50891 );
and ( n52086 , n50891 , n50893 );
and ( n52087 , n50890 , n50893 );
or ( n52088 , n52085 , n52086 , n52087 );
buf ( n52089 , n11015 );
and ( n52090 , n11769 , n10239 );
xor ( n52091 , n52089 , n52090 );
and ( n52092 , n12320 , n9348 );
xor ( n52093 , n52091 , n52092 );
xor ( n52094 , n52088 , n52093 );
and ( n52095 , n8718 , n13256 );
and ( n52096 , n9400 , n12531 );
xor ( n52097 , n52095 , n52096 );
and ( n52098 , n10291 , n11718 );
xor ( n52099 , n52097 , n52098 );
xor ( n52100 , n52094 , n52099 );
xor ( n52101 , n52084 , n52100 );
xor ( n52102 , n52075 , n52101 );
xor ( n52103 , n52066 , n52102 );
xor ( n52104 , n51993 , n52103 );
xor ( n52105 , n51984 , n52104 );
and ( n52106 , n50983 , n51022 );
and ( n52107 , n50914 , n50951 );
and ( n52108 , n50951 , n50977 );
and ( n52109 , n50914 , n50977 );
or ( n52110 , n52107 , n52108 , n52109 );
and ( n52111 , n50987 , n51021 );
xor ( n52112 , n52110 , n52111 );
and ( n52113 , n50956 , n50960 );
and ( n52114 , n50960 , n50976 );
and ( n52115 , n50956 , n50976 );
or ( n52116 , n52113 , n52114 , n52115 );
and ( n52117 , n50938 , n50943 );
and ( n52118 , n50943 , n50949 );
and ( n52119 , n50938 , n50949 );
or ( n52120 , n52117 , n52118 , n52119 );
and ( n52121 , n50928 , n50929 );
and ( n52122 , n50929 , n50931 );
and ( n52123 , n50928 , n50931 );
or ( n52124 , n52121 , n52122 , n52123 );
and ( n52125 , n50939 , n50940 );
and ( n52126 , n50940 , n50942 );
and ( n52127 , n50939 , n50942 );
or ( n52128 , n52125 , n52126 , n52127 );
xor ( n52129 , n52124 , n52128 );
and ( n52130 , n7385 , n15691 );
and ( n52131 , n7808 , n14838 );
xor ( n52132 , n52130 , n52131 );
and ( n52133 , n8079 , n14044 );
xor ( n52134 , n52132 , n52133 );
xor ( n52135 , n52129 , n52134 );
xor ( n52136 , n52120 , n52135 );
and ( n52137 , n50945 , n50946 );
and ( n52138 , n50946 , n50948 );
and ( n52139 , n50945 , n50948 );
or ( n52140 , n52137 , n52138 , n52139 );
and ( n52141 , n6187 , n18407 );
and ( n52142 , n6569 , n17422 );
xor ( n52143 , n52141 , n52142 );
and ( n52144 , n6816 , n16550 );
xor ( n52145 , n52143 , n52144 );
xor ( n52146 , n52140 , n52145 );
and ( n52147 , n4959 , n20976 );
and ( n52148 , n5459 , n20156 );
xor ( n52149 , n52147 , n52148 );
and ( n52150 , n5819 , n19222 );
xor ( n52151 , n52149 , n52150 );
xor ( n52152 , n52146 , n52151 );
xor ( n52153 , n52136 , n52152 );
xor ( n52154 , n52116 , n52153 );
and ( n52155 , n50965 , n50969 );
and ( n52156 , n50969 , n50975 );
and ( n52157 , n50965 , n50975 );
or ( n52158 , n52155 , n52156 , n52157 );
and ( n52159 , n50995 , n51000 );
and ( n52160 , n51000 , n51006 );
and ( n52161 , n50995 , n51006 );
or ( n52162 , n52159 , n52160 , n52161 );
xor ( n52163 , n52158 , n52162 );
and ( n52164 , n50971 , n50972 );
and ( n52165 , n50972 , n50974 );
and ( n52166 , n50971 , n50974 );
or ( n52167 , n52164 , n52165 , n52166 );
and ( n52168 , n50996 , n50997 );
and ( n52169 , n50997 , n50999 );
and ( n52170 , n50996 , n50999 );
or ( n52171 , n52168 , n52169 , n52170 );
xor ( n52172 , n52167 , n52171 );
and ( n52173 , n4132 , n24137 );
and ( n52174 , n4438 , n23075 );
xor ( n52175 , n52173 , n52174 );
and ( n52176 , n4766 , n22065 );
xor ( n52177 , n52175 , n52176 );
xor ( n52178 , n52172 , n52177 );
xor ( n52179 , n52163 , n52178 );
xor ( n52180 , n52154 , n52179 );
xor ( n52181 , n52112 , n52180 );
xor ( n52182 , n52106 , n52181 );
and ( n52183 , n50991 , n51007 );
and ( n52184 , n51007 , n51020 );
and ( n52185 , n50991 , n51020 );
or ( n52186 , n52183 , n52184 , n52185 );
and ( n52187 , n51012 , n51013 );
and ( n52188 , n51013 , n51019 );
and ( n52189 , n51012 , n51019 );
or ( n52190 , n52187 , n52188 , n52189 );
and ( n52191 , n51002 , n51003 );
and ( n52192 , n51003 , n51005 );
and ( n52193 , n51002 , n51005 );
or ( n52194 , n52191 , n52192 , n52193 );
and ( n52195 , n3182 , n27296 );
and ( n52196 , n3545 , n26216 );
xor ( n52197 , n52195 , n52196 );
and ( n52198 , n3801 , n25163 );
xor ( n52199 , n52197 , n52198 );
xor ( n52200 , n52194 , n52199 );
and ( n52201 , n2462 , n30629 );
and ( n52202 , n2779 , n29508 );
xor ( n52203 , n52201 , n52202 );
and ( n52204 , n3024 , n28406 );
xor ( n52205 , n52203 , n52204 );
xor ( n52206 , n52200 , n52205 );
xor ( n52207 , n52190 , n52206 );
and ( n52208 , n51015 , n51016 );
and ( n52209 , n51016 , n51018 );
and ( n52210 , n51015 , n51018 );
or ( n52211 , n52208 , n52209 , n52210 );
not ( n52212 , n1933 );
and ( n52213 , n34193 , n1933 );
nor ( n52214 , n52212 , n52213 );
and ( n52215 , n2120 , n32999 );
xor ( n52216 , n52214 , n52215 );
and ( n52217 , n2324 , n31761 );
xor ( n52218 , n52216 , n52217 );
xor ( n52219 , n52211 , n52218 );
xor ( n52220 , n52207 , n52219 );
xor ( n52221 , n52186 , n52220 );
xor ( n52222 , n52182 , n52221 );
xor ( n52223 , n52105 , n52222 );
xor ( n52224 , n51980 , n52223 );
xor ( n52225 , n51898 , n52224 );
xor ( n52226 , n51889 , n52225 );
and ( n52227 , n50680 , n50683 );
and ( n52228 , n50683 , n51027 );
and ( n52229 , n50680 , n51027 );
or ( n52230 , n52227 , n52228 , n52229 );
xor ( n52231 , n52226 , n52230 );
and ( n52232 , n51028 , n51032 );
and ( n52233 , n51033 , n51036 );
or ( n52234 , n52232 , n52233 );
xor ( n52235 , n52231 , n52234 );
buf ( n52236 , n52235 );
buf ( n52237 , n52236 );
not ( n52238 , n52237 );
nor ( n52239 , n52238 , n8739 );
xor ( n52240 , n51881 , n52239 );
and ( n52241 , n50676 , n51041 );
and ( n52242 , n51042 , n51045 );
or ( n52243 , n52241 , n52242 );
xor ( n52244 , n52240 , n52243 );
buf ( n52245 , n52244 );
buf ( n52246 , n52245 );
not ( n52247 , n52246 );
buf ( n52248 , n577 );
not ( n52249 , n52248 );
nor ( n52250 , n52247 , n52249 );
xor ( n52251 , n51507 , n52250 );
xor ( n52252 , n51057 , n51504 );
nor ( n52253 , n51049 , n52249 );
and ( n52254 , n52252 , n52253 );
xor ( n52255 , n52252 , n52253 );
xor ( n52256 , n51061 , n51502 );
nor ( n52257 , n49850 , n52249 );
and ( n52258 , n52256 , n52257 );
xor ( n52259 , n52256 , n52257 );
xor ( n52260 , n51065 , n51500 );
nor ( n52261 , n48650 , n52249 );
and ( n52262 , n52260 , n52261 );
xor ( n52263 , n52260 , n52261 );
xor ( n52264 , n51069 , n51498 );
nor ( n52265 , n47449 , n52249 );
and ( n52266 , n52264 , n52265 );
xor ( n52267 , n52264 , n52265 );
xor ( n52268 , n51073 , n51496 );
nor ( n52269 , n46248 , n52249 );
and ( n52270 , n52268 , n52269 );
xor ( n52271 , n52268 , n52269 );
xor ( n52272 , n51077 , n51494 );
nor ( n52273 , n45047 , n52249 );
and ( n52274 , n52272 , n52273 );
xor ( n52275 , n52272 , n52273 );
xor ( n52276 , n51081 , n51492 );
nor ( n52277 , n43843 , n52249 );
and ( n52278 , n52276 , n52277 );
xor ( n52279 , n52276 , n52277 );
xor ( n52280 , n51085 , n51490 );
nor ( n52281 , n42641 , n52249 );
and ( n52282 , n52280 , n52281 );
xor ( n52283 , n52280 , n52281 );
xor ( n52284 , n51089 , n51488 );
nor ( n52285 , n41437 , n52249 );
and ( n52286 , n52284 , n52285 );
xor ( n52287 , n52284 , n52285 );
xor ( n52288 , n51093 , n51486 );
nor ( n52289 , n40232 , n52249 );
and ( n52290 , n52288 , n52289 );
xor ( n52291 , n52288 , n52289 );
xor ( n52292 , n51097 , n51484 );
nor ( n52293 , n39027 , n52249 );
and ( n52294 , n52292 , n52293 );
xor ( n52295 , n52292 , n52293 );
xor ( n52296 , n51101 , n51482 );
nor ( n52297 , n37825 , n52249 );
and ( n52298 , n52296 , n52297 );
xor ( n52299 , n52296 , n52297 );
xor ( n52300 , n51105 , n51480 );
nor ( n52301 , n36620 , n52249 );
and ( n52302 , n52300 , n52301 );
xor ( n52303 , n52300 , n52301 );
xor ( n52304 , n51109 , n51478 );
nor ( n52305 , n35419 , n52249 );
and ( n52306 , n52304 , n52305 );
xor ( n52307 , n52304 , n52305 );
xor ( n52308 , n51113 , n51476 );
nor ( n52309 , n34224 , n52249 );
and ( n52310 , n52308 , n52309 );
xor ( n52311 , n52308 , n52309 );
xor ( n52312 , n51117 , n51474 );
nor ( n52313 , n33033 , n52249 );
and ( n52314 , n52312 , n52313 );
xor ( n52315 , n52312 , n52313 );
xor ( n52316 , n51121 , n51472 );
nor ( n52317 , n31867 , n52249 );
and ( n52318 , n52316 , n52317 );
xor ( n52319 , n52316 , n52317 );
xor ( n52320 , n51125 , n51470 );
nor ( n52321 , n30725 , n52249 );
and ( n52322 , n52320 , n52321 );
xor ( n52323 , n52320 , n52321 );
xor ( n52324 , n51129 , n51468 );
nor ( n52325 , n29596 , n52249 );
and ( n52326 , n52324 , n52325 );
xor ( n52327 , n52324 , n52325 );
xor ( n52328 , n51133 , n51466 );
nor ( n52329 , n28487 , n52249 );
and ( n52330 , n52328 , n52329 );
xor ( n52331 , n52328 , n52329 );
xor ( n52332 , n51137 , n51464 );
nor ( n52333 , n27397 , n52249 );
and ( n52334 , n52332 , n52333 );
xor ( n52335 , n52332 , n52333 );
xor ( n52336 , n51141 , n51462 );
nor ( n52337 , n26326 , n52249 );
and ( n52338 , n52336 , n52337 );
xor ( n52339 , n52336 , n52337 );
xor ( n52340 , n51145 , n51460 );
nor ( n52341 , n25272 , n52249 );
and ( n52342 , n52340 , n52341 );
xor ( n52343 , n52340 , n52341 );
xor ( n52344 , n51149 , n51458 );
nor ( n52345 , n24242 , n52249 );
and ( n52346 , n52344 , n52345 );
xor ( n52347 , n52344 , n52345 );
xor ( n52348 , n51153 , n51456 );
nor ( n52349 , n23225 , n52249 );
and ( n52350 , n52348 , n52349 );
xor ( n52351 , n52348 , n52349 );
xor ( n52352 , n51157 , n51454 );
nor ( n52353 , n22231 , n52249 );
and ( n52354 , n52352 , n52353 );
xor ( n52355 , n52352 , n52353 );
xor ( n52356 , n51161 , n51452 );
nor ( n52357 , n21258 , n52249 );
and ( n52358 , n52356 , n52357 );
xor ( n52359 , n52356 , n52357 );
xor ( n52360 , n51165 , n51450 );
nor ( n52361 , n20303 , n52249 );
and ( n52362 , n52360 , n52361 );
xor ( n52363 , n52360 , n52361 );
xor ( n52364 , n51169 , n51448 );
nor ( n52365 , n19365 , n52249 );
and ( n52366 , n52364 , n52365 );
xor ( n52367 , n52364 , n52365 );
xor ( n52368 , n51173 , n51446 );
nor ( n52369 , n18448 , n52249 );
and ( n52370 , n52368 , n52369 );
xor ( n52371 , n52368 , n52369 );
xor ( n52372 , n51177 , n51444 );
nor ( n52373 , n17548 , n52249 );
and ( n52374 , n52372 , n52373 );
xor ( n52375 , n52372 , n52373 );
xor ( n52376 , n51181 , n51442 );
nor ( n52377 , n16669 , n52249 );
and ( n52378 , n52376 , n52377 );
xor ( n52379 , n52376 , n52377 );
xor ( n52380 , n51185 , n51440 );
nor ( n52381 , n15809 , n52249 );
and ( n52382 , n52380 , n52381 );
xor ( n52383 , n52380 , n52381 );
xor ( n52384 , n51189 , n51438 );
nor ( n52385 , n14968 , n52249 );
and ( n52386 , n52384 , n52385 );
xor ( n52387 , n52384 , n52385 );
xor ( n52388 , n51193 , n51436 );
nor ( n52389 , n14147 , n52249 );
and ( n52390 , n52388 , n52389 );
xor ( n52391 , n52388 , n52389 );
xor ( n52392 , n51197 , n51434 );
nor ( n52393 , n13349 , n52249 );
and ( n52394 , n52392 , n52393 );
xor ( n52395 , n52392 , n52393 );
xor ( n52396 , n51201 , n51432 );
nor ( n52397 , n12564 , n52249 );
and ( n52398 , n52396 , n52397 );
xor ( n52399 , n52396 , n52397 );
xor ( n52400 , n51205 , n51430 );
nor ( n52401 , n11799 , n52249 );
and ( n52402 , n52400 , n52401 );
xor ( n52403 , n52400 , n52401 );
xor ( n52404 , n51209 , n51428 );
nor ( n52405 , n11050 , n52249 );
and ( n52406 , n52404 , n52405 );
xor ( n52407 , n52404 , n52405 );
xor ( n52408 , n51213 , n51426 );
nor ( n52409 , n10321 , n52249 );
and ( n52410 , n52408 , n52409 );
xor ( n52411 , n52408 , n52409 );
xor ( n52412 , n51217 , n51424 );
nor ( n52413 , n9429 , n52249 );
and ( n52414 , n52412 , n52413 );
xor ( n52415 , n52412 , n52413 );
xor ( n52416 , n51221 , n51422 );
nor ( n52417 , n8949 , n52249 );
and ( n52418 , n52416 , n52417 );
xor ( n52419 , n52416 , n52417 );
xor ( n52420 , n51225 , n51420 );
nor ( n52421 , n9437 , n52249 );
and ( n52422 , n52420 , n52421 );
xor ( n52423 , n52420 , n52421 );
xor ( n52424 , n51229 , n51418 );
nor ( n52425 , n9446 , n52249 );
and ( n52426 , n52424 , n52425 );
xor ( n52427 , n52424 , n52425 );
xor ( n52428 , n51233 , n51416 );
nor ( n52429 , n9455 , n52249 );
and ( n52430 , n52428 , n52429 );
xor ( n52431 , n52428 , n52429 );
xor ( n52432 , n51237 , n51414 );
nor ( n52433 , n9464 , n52249 );
and ( n52434 , n52432 , n52433 );
xor ( n52435 , n52432 , n52433 );
xor ( n52436 , n51241 , n51412 );
nor ( n52437 , n9473 , n52249 );
and ( n52438 , n52436 , n52437 );
xor ( n52439 , n52436 , n52437 );
xor ( n52440 , n51245 , n51410 );
nor ( n52441 , n9482 , n52249 );
and ( n52442 , n52440 , n52441 );
xor ( n52443 , n52440 , n52441 );
xor ( n52444 , n51249 , n51408 );
nor ( n52445 , n9491 , n52249 );
and ( n52446 , n52444 , n52445 );
xor ( n52447 , n52444 , n52445 );
xor ( n52448 , n51253 , n51406 );
nor ( n52449 , n9500 , n52249 );
and ( n52450 , n52448 , n52449 );
xor ( n52451 , n52448 , n52449 );
xor ( n52452 , n51257 , n51404 );
nor ( n52453 , n9509 , n52249 );
and ( n52454 , n52452 , n52453 );
xor ( n52455 , n52452 , n52453 );
xor ( n52456 , n51261 , n51402 );
nor ( n52457 , n9518 , n52249 );
and ( n52458 , n52456 , n52457 );
xor ( n52459 , n52456 , n52457 );
xor ( n52460 , n51265 , n51400 );
nor ( n52461 , n9527 , n52249 );
and ( n52462 , n52460 , n52461 );
xor ( n52463 , n52460 , n52461 );
xor ( n52464 , n51269 , n51398 );
nor ( n52465 , n9536 , n52249 );
and ( n52466 , n52464 , n52465 );
xor ( n52467 , n52464 , n52465 );
xor ( n52468 , n51273 , n51396 );
nor ( n52469 , n9545 , n52249 );
and ( n52470 , n52468 , n52469 );
xor ( n52471 , n52468 , n52469 );
xor ( n52472 , n51277 , n51394 );
nor ( n52473 , n9554 , n52249 );
and ( n52474 , n52472 , n52473 );
xor ( n52475 , n52472 , n52473 );
xor ( n52476 , n51281 , n51392 );
nor ( n52477 , n9563 , n52249 );
and ( n52478 , n52476 , n52477 );
xor ( n52479 , n52476 , n52477 );
xor ( n52480 , n51285 , n51390 );
nor ( n52481 , n9572 , n52249 );
and ( n52482 , n52480 , n52481 );
xor ( n52483 , n52480 , n52481 );
xor ( n52484 , n51289 , n51388 );
nor ( n52485 , n9581 , n52249 );
and ( n52486 , n52484 , n52485 );
xor ( n52487 , n52484 , n52485 );
xor ( n52488 , n51293 , n51386 );
nor ( n52489 , n9590 , n52249 );
and ( n52490 , n52488 , n52489 );
xor ( n52491 , n52488 , n52489 );
xor ( n52492 , n51297 , n51384 );
nor ( n52493 , n9599 , n52249 );
and ( n52494 , n52492 , n52493 );
xor ( n52495 , n52492 , n52493 );
xor ( n52496 , n51301 , n51382 );
nor ( n52497 , n9608 , n52249 );
and ( n52498 , n52496 , n52497 );
xor ( n52499 , n52496 , n52497 );
xor ( n52500 , n51305 , n51380 );
nor ( n52501 , n9617 , n52249 );
and ( n52502 , n52500 , n52501 );
xor ( n52503 , n52500 , n52501 );
xor ( n52504 , n51309 , n51378 );
nor ( n52505 , n9626 , n52249 );
and ( n52506 , n52504 , n52505 );
xor ( n52507 , n52504 , n52505 );
xor ( n52508 , n51313 , n51376 );
nor ( n52509 , n9635 , n52249 );
and ( n52510 , n52508 , n52509 );
xor ( n52511 , n52508 , n52509 );
xor ( n52512 , n51317 , n51374 );
nor ( n52513 , n9644 , n52249 );
and ( n52514 , n52512 , n52513 );
xor ( n52515 , n52512 , n52513 );
xor ( n52516 , n51321 , n51372 );
nor ( n52517 , n9653 , n52249 );
and ( n52518 , n52516 , n52517 );
xor ( n52519 , n52516 , n52517 );
xor ( n52520 , n51325 , n51370 );
nor ( n52521 , n9662 , n52249 );
and ( n52522 , n52520 , n52521 );
xor ( n52523 , n52520 , n52521 );
xor ( n52524 , n51329 , n51368 );
nor ( n52525 , n9671 , n52249 );
and ( n52526 , n52524 , n52525 );
xor ( n52527 , n52524 , n52525 );
xor ( n52528 , n51333 , n51366 );
nor ( n52529 , n9680 , n52249 );
and ( n52530 , n52528 , n52529 );
xor ( n52531 , n52528 , n52529 );
xor ( n52532 , n51337 , n51364 );
nor ( n52533 , n9689 , n52249 );
and ( n52534 , n52532 , n52533 );
xor ( n52535 , n52532 , n52533 );
xor ( n52536 , n51341 , n51362 );
nor ( n52537 , n9698 , n52249 );
and ( n52538 , n52536 , n52537 );
xor ( n52539 , n52536 , n52537 );
xor ( n52540 , n51345 , n51360 );
nor ( n52541 , n9707 , n52249 );
and ( n52542 , n52540 , n52541 );
xor ( n52543 , n52540 , n52541 );
xor ( n52544 , n51349 , n51358 );
nor ( n52545 , n9716 , n52249 );
and ( n52546 , n52544 , n52545 );
xor ( n52547 , n52544 , n52545 );
xor ( n52548 , n51353 , n51356 );
nor ( n52549 , n9725 , n52249 );
and ( n52550 , n52548 , n52549 );
xor ( n52551 , n52548 , n52549 );
xor ( n52552 , n51354 , n51355 );
nor ( n52553 , n9734 , n52249 );
and ( n52554 , n52552 , n52553 );
xor ( n52555 , n52552 , n52553 );
nor ( n52556 , n9752 , n51051 );
nor ( n52557 , n9743 , n52249 );
and ( n52558 , n52556 , n52557 );
and ( n52559 , n52555 , n52558 );
or ( n52560 , n52554 , n52559 );
and ( n52561 , n52551 , n52560 );
or ( n52562 , n52550 , n52561 );
and ( n52563 , n52547 , n52562 );
or ( n52564 , n52546 , n52563 );
and ( n52565 , n52543 , n52564 );
or ( n52566 , n52542 , n52565 );
and ( n52567 , n52539 , n52566 );
or ( n52568 , n52538 , n52567 );
and ( n52569 , n52535 , n52568 );
or ( n52570 , n52534 , n52569 );
and ( n52571 , n52531 , n52570 );
or ( n52572 , n52530 , n52571 );
and ( n52573 , n52527 , n52572 );
or ( n52574 , n52526 , n52573 );
and ( n52575 , n52523 , n52574 );
or ( n52576 , n52522 , n52575 );
and ( n52577 , n52519 , n52576 );
or ( n52578 , n52518 , n52577 );
and ( n52579 , n52515 , n52578 );
or ( n52580 , n52514 , n52579 );
and ( n52581 , n52511 , n52580 );
or ( n52582 , n52510 , n52581 );
and ( n52583 , n52507 , n52582 );
or ( n52584 , n52506 , n52583 );
and ( n52585 , n52503 , n52584 );
or ( n52586 , n52502 , n52585 );
and ( n52587 , n52499 , n52586 );
or ( n52588 , n52498 , n52587 );
and ( n52589 , n52495 , n52588 );
or ( n52590 , n52494 , n52589 );
and ( n52591 , n52491 , n52590 );
or ( n52592 , n52490 , n52591 );
and ( n52593 , n52487 , n52592 );
or ( n52594 , n52486 , n52593 );
and ( n52595 , n52483 , n52594 );
or ( n52596 , n52482 , n52595 );
and ( n52597 , n52479 , n52596 );
or ( n52598 , n52478 , n52597 );
and ( n52599 , n52475 , n52598 );
or ( n52600 , n52474 , n52599 );
and ( n52601 , n52471 , n52600 );
or ( n52602 , n52470 , n52601 );
and ( n52603 , n52467 , n52602 );
or ( n52604 , n52466 , n52603 );
and ( n52605 , n52463 , n52604 );
or ( n52606 , n52462 , n52605 );
and ( n52607 , n52459 , n52606 );
or ( n52608 , n52458 , n52607 );
and ( n52609 , n52455 , n52608 );
or ( n52610 , n52454 , n52609 );
and ( n52611 , n52451 , n52610 );
or ( n52612 , n52450 , n52611 );
and ( n52613 , n52447 , n52612 );
or ( n52614 , n52446 , n52613 );
and ( n52615 , n52443 , n52614 );
or ( n52616 , n52442 , n52615 );
and ( n52617 , n52439 , n52616 );
or ( n52618 , n52438 , n52617 );
and ( n52619 , n52435 , n52618 );
or ( n52620 , n52434 , n52619 );
and ( n52621 , n52431 , n52620 );
or ( n52622 , n52430 , n52621 );
and ( n52623 , n52427 , n52622 );
or ( n52624 , n52426 , n52623 );
and ( n52625 , n52423 , n52624 );
or ( n52626 , n52422 , n52625 );
and ( n52627 , n52419 , n52626 );
or ( n52628 , n52418 , n52627 );
and ( n52629 , n52415 , n52628 );
or ( n52630 , n52414 , n52629 );
and ( n52631 , n52411 , n52630 );
or ( n52632 , n52410 , n52631 );
and ( n52633 , n52407 , n52632 );
or ( n52634 , n52406 , n52633 );
and ( n52635 , n52403 , n52634 );
or ( n52636 , n52402 , n52635 );
and ( n52637 , n52399 , n52636 );
or ( n52638 , n52398 , n52637 );
and ( n52639 , n52395 , n52638 );
or ( n52640 , n52394 , n52639 );
and ( n52641 , n52391 , n52640 );
or ( n52642 , n52390 , n52641 );
and ( n52643 , n52387 , n52642 );
or ( n52644 , n52386 , n52643 );
and ( n52645 , n52383 , n52644 );
or ( n52646 , n52382 , n52645 );
and ( n52647 , n52379 , n52646 );
or ( n52648 , n52378 , n52647 );
and ( n52649 , n52375 , n52648 );
or ( n52650 , n52374 , n52649 );
and ( n52651 , n52371 , n52650 );
or ( n52652 , n52370 , n52651 );
and ( n52653 , n52367 , n52652 );
or ( n52654 , n52366 , n52653 );
and ( n52655 , n52363 , n52654 );
or ( n52656 , n52362 , n52655 );
and ( n52657 , n52359 , n52656 );
or ( n52658 , n52358 , n52657 );
and ( n52659 , n52355 , n52658 );
or ( n52660 , n52354 , n52659 );
and ( n52661 , n52351 , n52660 );
or ( n52662 , n52350 , n52661 );
and ( n52663 , n52347 , n52662 );
or ( n52664 , n52346 , n52663 );
and ( n52665 , n52343 , n52664 );
or ( n52666 , n52342 , n52665 );
and ( n52667 , n52339 , n52666 );
or ( n52668 , n52338 , n52667 );
and ( n52669 , n52335 , n52668 );
or ( n52670 , n52334 , n52669 );
and ( n52671 , n52331 , n52670 );
or ( n52672 , n52330 , n52671 );
and ( n52673 , n52327 , n52672 );
or ( n52674 , n52326 , n52673 );
and ( n52675 , n52323 , n52674 );
or ( n52676 , n52322 , n52675 );
and ( n52677 , n52319 , n52676 );
or ( n52678 , n52318 , n52677 );
and ( n52679 , n52315 , n52678 );
or ( n52680 , n52314 , n52679 );
and ( n52681 , n52311 , n52680 );
or ( n52682 , n52310 , n52681 );
and ( n52683 , n52307 , n52682 );
or ( n52684 , n52306 , n52683 );
and ( n52685 , n52303 , n52684 );
or ( n52686 , n52302 , n52685 );
and ( n52687 , n52299 , n52686 );
or ( n52688 , n52298 , n52687 );
and ( n52689 , n52295 , n52688 );
or ( n52690 , n52294 , n52689 );
and ( n52691 , n52291 , n52690 );
or ( n52692 , n52290 , n52691 );
and ( n52693 , n52287 , n52692 );
or ( n52694 , n52286 , n52693 );
and ( n52695 , n52283 , n52694 );
or ( n52696 , n52282 , n52695 );
and ( n52697 , n52279 , n52696 );
or ( n52698 , n52278 , n52697 );
and ( n52699 , n52275 , n52698 );
or ( n52700 , n52274 , n52699 );
and ( n52701 , n52271 , n52700 );
or ( n52702 , n52270 , n52701 );
and ( n52703 , n52267 , n52702 );
or ( n52704 , n52266 , n52703 );
and ( n52705 , n52263 , n52704 );
or ( n52706 , n52262 , n52705 );
and ( n52707 , n52259 , n52706 );
or ( n52708 , n52258 , n52707 );
and ( n52709 , n52255 , n52708 );
or ( n52710 , n52254 , n52709 );
xor ( n52711 , n52251 , n52710 );
and ( n52712 , n33403 , n2136 );
nor ( n52713 , n2137 , n52712 );
nor ( n52714 , n2343 , n32231 );
xor ( n52715 , n52713 , n52714 );
and ( n52716 , n51509 , n51510 );
and ( n52717 , n51511 , n51514 );
or ( n52718 , n52716 , n52717 );
xor ( n52719 , n52715 , n52718 );
nor ( n52720 , n2566 , n31083 );
xor ( n52721 , n52719 , n52720 );
and ( n52722 , n51515 , n51516 );
and ( n52723 , n51517 , n51520 );
or ( n52724 , n52722 , n52723 );
xor ( n52725 , n52721 , n52724 );
nor ( n52726 , n2797 , n29948 );
xor ( n52727 , n52725 , n52726 );
and ( n52728 , n51521 , n51522 );
and ( n52729 , n51523 , n51526 );
or ( n52730 , n52728 , n52729 );
xor ( n52731 , n52727 , n52730 );
nor ( n52732 , n3043 , n28833 );
xor ( n52733 , n52731 , n52732 );
and ( n52734 , n51527 , n51528 );
and ( n52735 , n51529 , n51532 );
or ( n52736 , n52734 , n52735 );
xor ( n52737 , n52733 , n52736 );
nor ( n52738 , n3300 , n27737 );
xor ( n52739 , n52737 , n52738 );
and ( n52740 , n51533 , n51534 );
and ( n52741 , n51535 , n51538 );
or ( n52742 , n52740 , n52741 );
xor ( n52743 , n52739 , n52742 );
nor ( n52744 , n3570 , n26660 );
xor ( n52745 , n52743 , n52744 );
and ( n52746 , n51539 , n51540 );
and ( n52747 , n51541 , n51544 );
or ( n52748 , n52746 , n52747 );
xor ( n52749 , n52745 , n52748 );
nor ( n52750 , n3853 , n25600 );
xor ( n52751 , n52749 , n52750 );
and ( n52752 , n51545 , n51546 );
and ( n52753 , n51547 , n51550 );
or ( n52754 , n52752 , n52753 );
xor ( n52755 , n52751 , n52754 );
nor ( n52756 , n4151 , n24564 );
xor ( n52757 , n52755 , n52756 );
and ( n52758 , n51551 , n51552 );
and ( n52759 , n51553 , n51556 );
or ( n52760 , n52758 , n52759 );
xor ( n52761 , n52757 , n52760 );
nor ( n52762 , n4458 , n23541 );
xor ( n52763 , n52761 , n52762 );
and ( n52764 , n51557 , n51558 );
and ( n52765 , n51559 , n51562 );
or ( n52766 , n52764 , n52765 );
xor ( n52767 , n52763 , n52766 );
nor ( n52768 , n4786 , n22541 );
xor ( n52769 , n52767 , n52768 );
and ( n52770 , n51563 , n51564 );
and ( n52771 , n51565 , n51568 );
or ( n52772 , n52770 , n52771 );
xor ( n52773 , n52769 , n52772 );
nor ( n52774 , n5126 , n21562 );
xor ( n52775 , n52773 , n52774 );
and ( n52776 , n51569 , n51570 );
and ( n52777 , n51571 , n51574 );
or ( n52778 , n52776 , n52777 );
xor ( n52779 , n52775 , n52778 );
nor ( n52780 , n5477 , n20601 );
xor ( n52781 , n52779 , n52780 );
and ( n52782 , n51575 , n51576 );
and ( n52783 , n51577 , n51580 );
or ( n52784 , n52782 , n52783 );
xor ( n52785 , n52781 , n52784 );
nor ( n52786 , n5838 , n19657 );
xor ( n52787 , n52785 , n52786 );
and ( n52788 , n51581 , n51582 );
and ( n52789 , n51583 , n51586 );
or ( n52790 , n52788 , n52789 );
xor ( n52791 , n52787 , n52790 );
nor ( n52792 , n6212 , n18734 );
xor ( n52793 , n52791 , n52792 );
and ( n52794 , n51587 , n51588 );
and ( n52795 , n51589 , n51592 );
or ( n52796 , n52794 , n52795 );
xor ( n52797 , n52793 , n52796 );
nor ( n52798 , n6596 , n17828 );
xor ( n52799 , n52797 , n52798 );
and ( n52800 , n51593 , n51594 );
and ( n52801 , n51595 , n51598 );
or ( n52802 , n52800 , n52801 );
xor ( n52803 , n52799 , n52802 );
nor ( n52804 , n6997 , n16943 );
xor ( n52805 , n52803 , n52804 );
and ( n52806 , n51599 , n51600 );
and ( n52807 , n51601 , n51604 );
or ( n52808 , n52806 , n52807 );
xor ( n52809 , n52805 , n52808 );
nor ( n52810 , n7413 , n16077 );
xor ( n52811 , n52809 , n52810 );
and ( n52812 , n51605 , n51606 );
and ( n52813 , n51607 , n51610 );
or ( n52814 , n52812 , n52813 );
xor ( n52815 , n52811 , n52814 );
nor ( n52816 , n7841 , n15230 );
xor ( n52817 , n52815 , n52816 );
and ( n52818 , n51611 , n51612 );
and ( n52819 , n51613 , n51616 );
or ( n52820 , n52818 , n52819 );
xor ( n52821 , n52817 , n52820 );
nor ( n52822 , n8281 , n14403 );
xor ( n52823 , n52821 , n52822 );
and ( n52824 , n51617 , n51618 );
and ( n52825 , n51619 , n51622 );
or ( n52826 , n52824 , n52825 );
xor ( n52827 , n52823 , n52826 );
nor ( n52828 , n8737 , n13599 );
xor ( n52829 , n52827 , n52828 );
and ( n52830 , n51623 , n51624 );
and ( n52831 , n51625 , n51628 );
or ( n52832 , n52830 , n52831 );
xor ( n52833 , n52829 , n52832 );
nor ( n52834 , n9420 , n12808 );
xor ( n52835 , n52833 , n52834 );
and ( n52836 , n51629 , n51630 );
and ( n52837 , n51631 , n51634 );
or ( n52838 , n52836 , n52837 );
xor ( n52839 , n52835 , n52838 );
nor ( n52840 , n10312 , n12037 );
xor ( n52841 , n52839 , n52840 );
and ( n52842 , n51635 , n51636 );
and ( n52843 , n51637 , n51640 );
or ( n52844 , n52842 , n52843 );
xor ( n52845 , n52841 , n52844 );
nor ( n52846 , n11041 , n11282 );
xor ( n52847 , n52845 , n52846 );
and ( n52848 , n51641 , n51642 );
and ( n52849 , n51643 , n51646 );
or ( n52850 , n52848 , n52849 );
xor ( n52851 , n52847 , n52850 );
nor ( n52852 , n11790 , n10547 );
xor ( n52853 , n52851 , n52852 );
and ( n52854 , n51647 , n51648 );
and ( n52855 , n51649 , n51652 );
or ( n52856 , n52854 , n52855 );
xor ( n52857 , n52853 , n52856 );
nor ( n52858 , n12555 , n9829 );
xor ( n52859 , n52857 , n52858 );
and ( n52860 , n51653 , n51654 );
and ( n52861 , n51655 , n51658 );
or ( n52862 , n52860 , n52861 );
xor ( n52863 , n52859 , n52862 );
nor ( n52864 , n13340 , n8955 );
xor ( n52865 , n52863 , n52864 );
and ( n52866 , n51659 , n51660 );
and ( n52867 , n51661 , n51664 );
or ( n52868 , n52866 , n52867 );
xor ( n52869 , n52865 , n52868 );
nor ( n52870 , n14138 , n603 );
xor ( n52871 , n52869 , n52870 );
and ( n52872 , n51665 , n51666 );
and ( n52873 , n51667 , n51670 );
or ( n52874 , n52872 , n52873 );
xor ( n52875 , n52871 , n52874 );
nor ( n52876 , n14959 , n652 );
xor ( n52877 , n52875 , n52876 );
and ( n52878 , n51671 , n51672 );
and ( n52879 , n51673 , n51676 );
or ( n52880 , n52878 , n52879 );
xor ( n52881 , n52877 , n52880 );
nor ( n52882 , n15800 , n624 );
xor ( n52883 , n52881 , n52882 );
and ( n52884 , n51677 , n51678 );
and ( n52885 , n51679 , n51682 );
or ( n52886 , n52884 , n52885 );
xor ( n52887 , n52883 , n52886 );
nor ( n52888 , n16660 , n648 );
xor ( n52889 , n52887 , n52888 );
and ( n52890 , n51683 , n51684 );
and ( n52891 , n51685 , n51688 );
or ( n52892 , n52890 , n52891 );
xor ( n52893 , n52889 , n52892 );
nor ( n52894 , n17539 , n686 );
xor ( n52895 , n52893 , n52894 );
and ( n52896 , n51689 , n51690 );
and ( n52897 , n51691 , n51694 );
or ( n52898 , n52896 , n52897 );
xor ( n52899 , n52895 , n52898 );
nor ( n52900 , n18439 , n735 );
xor ( n52901 , n52899 , n52900 );
and ( n52902 , n51695 , n51696 );
and ( n52903 , n51697 , n51700 );
or ( n52904 , n52902 , n52903 );
xor ( n52905 , n52901 , n52904 );
nor ( n52906 , n19356 , n798 );
xor ( n52907 , n52905 , n52906 );
and ( n52908 , n51701 , n51702 );
and ( n52909 , n51703 , n51706 );
or ( n52910 , n52908 , n52909 );
xor ( n52911 , n52907 , n52910 );
nor ( n52912 , n20294 , n870 );
xor ( n52913 , n52911 , n52912 );
and ( n52914 , n51707 , n51708 );
and ( n52915 , n51709 , n51712 );
or ( n52916 , n52914 , n52915 );
xor ( n52917 , n52913 , n52916 );
nor ( n52918 , n21249 , n960 );
xor ( n52919 , n52917 , n52918 );
and ( n52920 , n51713 , n51714 );
and ( n52921 , n51715 , n51718 );
or ( n52922 , n52920 , n52921 );
xor ( n52923 , n52919 , n52922 );
nor ( n52924 , n22222 , n1064 );
xor ( n52925 , n52923 , n52924 );
and ( n52926 , n51719 , n51720 );
and ( n52927 , n51721 , n51724 );
or ( n52928 , n52926 , n52927 );
xor ( n52929 , n52925 , n52928 );
nor ( n52930 , n23216 , n1178 );
xor ( n52931 , n52929 , n52930 );
and ( n52932 , n51725 , n51726 );
and ( n52933 , n51727 , n51730 );
or ( n52934 , n52932 , n52933 );
xor ( n52935 , n52931 , n52934 );
nor ( n52936 , n24233 , n1305 );
xor ( n52937 , n52935 , n52936 );
and ( n52938 , n51731 , n51732 );
and ( n52939 , n51733 , n51736 );
or ( n52940 , n52938 , n52939 );
xor ( n52941 , n52937 , n52940 );
nor ( n52942 , n25263 , n1447 );
xor ( n52943 , n52941 , n52942 );
and ( n52944 , n51737 , n51738 );
and ( n52945 , n51739 , n51742 );
or ( n52946 , n52944 , n52945 );
xor ( n52947 , n52943 , n52946 );
nor ( n52948 , n26317 , n1600 );
xor ( n52949 , n52947 , n52948 );
and ( n52950 , n51743 , n51744 );
and ( n52951 , n51745 , n51748 );
or ( n52952 , n52950 , n52951 );
xor ( n52953 , n52949 , n52952 );
nor ( n52954 , n27388 , n1768 );
xor ( n52955 , n52953 , n52954 );
and ( n52956 , n51749 , n51750 );
and ( n52957 , n51751 , n51754 );
or ( n52958 , n52956 , n52957 );
xor ( n52959 , n52955 , n52958 );
nor ( n52960 , n28478 , n1947 );
xor ( n52961 , n52959 , n52960 );
and ( n52962 , n51755 , n51756 );
and ( n52963 , n51757 , n51760 );
or ( n52964 , n52962 , n52963 );
xor ( n52965 , n52961 , n52964 );
nor ( n52966 , n29587 , n2139 );
xor ( n52967 , n52965 , n52966 );
and ( n52968 , n51761 , n51762 );
and ( n52969 , n51763 , n51766 );
or ( n52970 , n52968 , n52969 );
xor ( n52971 , n52967 , n52970 );
nor ( n52972 , n30716 , n2345 );
xor ( n52973 , n52971 , n52972 );
and ( n52974 , n51767 , n51768 );
and ( n52975 , n51769 , n51772 );
or ( n52976 , n52974 , n52975 );
xor ( n52977 , n52973 , n52976 );
nor ( n52978 , n31858 , n2568 );
xor ( n52979 , n52977 , n52978 );
and ( n52980 , n51773 , n51774 );
and ( n52981 , n51775 , n51778 );
or ( n52982 , n52980 , n52981 );
xor ( n52983 , n52979 , n52982 );
nor ( n52984 , n33024 , n2799 );
xor ( n52985 , n52983 , n52984 );
and ( n52986 , n51779 , n51780 );
and ( n52987 , n51781 , n51784 );
or ( n52988 , n52986 , n52987 );
xor ( n52989 , n52985 , n52988 );
nor ( n52990 , n34215 , n3045 );
xor ( n52991 , n52989 , n52990 );
and ( n52992 , n51785 , n51786 );
and ( n52993 , n51787 , n51790 );
or ( n52994 , n52992 , n52993 );
xor ( n52995 , n52991 , n52994 );
nor ( n52996 , n35410 , n3302 );
xor ( n52997 , n52995 , n52996 );
and ( n52998 , n51791 , n51792 );
and ( n52999 , n51793 , n51796 );
or ( n53000 , n52998 , n52999 );
xor ( n53001 , n52997 , n53000 );
nor ( n53002 , n36611 , n3572 );
xor ( n53003 , n53001 , n53002 );
and ( n53004 , n51797 , n51798 );
and ( n53005 , n51799 , n51802 );
or ( n53006 , n53004 , n53005 );
xor ( n53007 , n53003 , n53006 );
nor ( n53008 , n37816 , n3855 );
xor ( n53009 , n53007 , n53008 );
and ( n53010 , n51803 , n51804 );
and ( n53011 , n51805 , n51808 );
or ( n53012 , n53010 , n53011 );
xor ( n53013 , n53009 , n53012 );
nor ( n53014 , n39018 , n4153 );
xor ( n53015 , n53013 , n53014 );
and ( n53016 , n51809 , n51810 );
and ( n53017 , n51811 , n51814 );
or ( n53018 , n53016 , n53017 );
xor ( n53019 , n53015 , n53018 );
nor ( n53020 , n40223 , n4460 );
xor ( n53021 , n53019 , n53020 );
and ( n53022 , n51815 , n51816 );
and ( n53023 , n51817 , n51820 );
or ( n53024 , n53022 , n53023 );
xor ( n53025 , n53021 , n53024 );
nor ( n53026 , n41428 , n4788 );
xor ( n53027 , n53025 , n53026 );
and ( n53028 , n51821 , n51822 );
and ( n53029 , n51823 , n51826 );
or ( n53030 , n53028 , n53029 );
xor ( n53031 , n53027 , n53030 );
nor ( n53032 , n42632 , n5128 );
xor ( n53033 , n53031 , n53032 );
and ( n53034 , n51827 , n51828 );
and ( n53035 , n51829 , n51832 );
or ( n53036 , n53034 , n53035 );
xor ( n53037 , n53033 , n53036 );
nor ( n53038 , n43834 , n5479 );
xor ( n53039 , n53037 , n53038 );
and ( n53040 , n51833 , n51834 );
and ( n53041 , n51835 , n51838 );
or ( n53042 , n53040 , n53041 );
xor ( n53043 , n53039 , n53042 );
nor ( n53044 , n45038 , n5840 );
xor ( n53045 , n53043 , n53044 );
and ( n53046 , n51839 , n51840 );
and ( n53047 , n51841 , n51844 );
or ( n53048 , n53046 , n53047 );
xor ( n53049 , n53045 , n53048 );
nor ( n53050 , n46239 , n6214 );
xor ( n53051 , n53049 , n53050 );
and ( n53052 , n51845 , n51846 );
and ( n53053 , n51847 , n51850 );
or ( n53054 , n53052 , n53053 );
xor ( n53055 , n53051 , n53054 );
nor ( n53056 , n47440 , n6598 );
xor ( n53057 , n53055 , n53056 );
and ( n53058 , n51851 , n51852 );
and ( n53059 , n51853 , n51856 );
or ( n53060 , n53058 , n53059 );
xor ( n53061 , n53057 , n53060 );
nor ( n53062 , n48641 , n6999 );
xor ( n53063 , n53061 , n53062 );
and ( n53064 , n51857 , n51858 );
and ( n53065 , n51859 , n51862 );
or ( n53066 , n53064 , n53065 );
xor ( n53067 , n53063 , n53066 );
nor ( n53068 , n49841 , n7415 );
xor ( n53069 , n53067 , n53068 );
and ( n53070 , n51863 , n51864 );
and ( n53071 , n51865 , n51868 );
or ( n53072 , n53070 , n53071 );
xor ( n53073 , n53069 , n53072 );
nor ( n53074 , n51040 , n7843 );
xor ( n53075 , n53073 , n53074 );
and ( n53076 , n51869 , n51870 );
and ( n53077 , n51871 , n51874 );
or ( n53078 , n53076 , n53077 );
xor ( n53079 , n53075 , n53078 );
nor ( n53080 , n52238 , n8283 );
xor ( n53081 , n53079 , n53080 );
and ( n53082 , n51875 , n51876 );
and ( n53083 , n51877 , n51880 );
or ( n53084 , n53082 , n53083 );
xor ( n53085 , n53081 , n53084 );
and ( n53086 , n51893 , n51897 );
and ( n53087 , n51897 , n52224 );
and ( n53088 , n51893 , n52224 );
or ( n53089 , n53086 , n53087 , n53088 );
and ( n53090 , n33774 , n2100 );
not ( n53091 , n2100 );
nor ( n53092 , n53090 , n53091 );
xor ( n53093 , n53089 , n53092 );
and ( n53094 , n51906 , n51910 );
and ( n53095 , n51910 , n51978 );
and ( n53096 , n51906 , n51978 );
or ( n53097 , n53094 , n53095 , n53096 );
and ( n53098 , n51902 , n51979 );
and ( n53099 , n51979 , n52223 );
and ( n53100 , n51902 , n52223 );
or ( n53101 , n53098 , n53099 , n53100 );
xor ( n53102 , n53097 , n53101 );
and ( n53103 , n51984 , n52104 );
and ( n53104 , n52104 , n52222 );
and ( n53105 , n51984 , n52222 );
or ( n53106 , n53103 , n53104 , n53105 );
and ( n53107 , n51915 , n51919 );
and ( n53108 , n51919 , n51977 );
and ( n53109 , n51915 , n51977 );
or ( n53110 , n53107 , n53108 , n53109 );
and ( n53111 , n51988 , n51992 );
and ( n53112 , n51992 , n52103 );
and ( n53113 , n51988 , n52103 );
or ( n53114 , n53111 , n53112 , n53113 );
xor ( n53115 , n53110 , n53114 );
and ( n53116 , n51946 , n51950 );
and ( n53117 , n51950 , n51956 );
and ( n53118 , n51946 , n51956 );
or ( n53119 , n53116 , n53117 , n53118 );
and ( n53120 , n51924 , n51928 );
and ( n53121 , n51928 , n51976 );
and ( n53122 , n51924 , n51976 );
or ( n53123 , n53120 , n53121 , n53122 );
xor ( n53124 , n53119 , n53123 );
and ( n53125 , n51933 , n51937 );
and ( n53126 , n51937 , n51975 );
and ( n53127 , n51933 , n51975 );
or ( n53128 , n53125 , n53126 , n53127 );
and ( n53129 , n52001 , n52026 );
and ( n53130 , n52026 , n52064 );
and ( n53131 , n52001 , n52064 );
or ( n53132 , n53129 , n53130 , n53131 );
xor ( n53133 , n53128 , n53132 );
and ( n53134 , n51942 , n51957 );
and ( n53135 , n51957 , n51974 );
and ( n53136 , n51942 , n51974 );
or ( n53137 , n53134 , n53135 , n53136 );
and ( n53138 , n52005 , n52009 );
and ( n53139 , n52009 , n52025 );
and ( n53140 , n52005 , n52025 );
or ( n53141 , n53138 , n53139 , n53140 );
xor ( n53142 , n53137 , n53141 );
and ( n53143 , n51962 , n51967 );
and ( n53144 , n51967 , n51973 );
and ( n53145 , n51962 , n51973 );
or ( n53146 , n53143 , n53144 , n53145 );
and ( n53147 , n51952 , n51953 );
and ( n53148 , n51953 , n51955 );
and ( n53149 , n51952 , n51955 );
or ( n53150 , n53147 , n53148 , n53149 );
and ( n53151 , n51963 , n51964 );
and ( n53152 , n51964 , n51966 );
and ( n53153 , n51963 , n51966 );
or ( n53154 , n53151 , n53152 , n53153 );
xor ( n53155 , n53150 , n53154 );
and ( n53156 , n30695 , n2739 );
and ( n53157 , n31836 , n2544 );
xor ( n53158 , n53156 , n53157 );
and ( n53159 , n32649 , n2298 );
xor ( n53160 , n53158 , n53159 );
xor ( n53161 , n53155 , n53160 );
xor ( n53162 , n53146 , n53161 );
and ( n53163 , n51969 , n51970 );
and ( n53164 , n51970 , n51972 );
and ( n53165 , n51969 , n51972 );
or ( n53166 , n53163 , n53164 , n53165 );
and ( n53167 , n27361 , n3495 );
and ( n53168 , n28456 , n3271 );
xor ( n53169 , n53167 , n53168 );
and ( n53170 , n29559 , n2981 );
xor ( n53171 , n53169 , n53170 );
xor ( n53172 , n53166 , n53171 );
and ( n53173 , n24214 , n4403 );
and ( n53174 , n25243 , n4102 );
xor ( n53175 , n53173 , n53174 );
and ( n53176 , n26296 , n3749 );
xor ( n53177 , n53175 , n53176 );
xor ( n53178 , n53172 , n53177 );
xor ( n53179 , n53162 , n53178 );
xor ( n53180 , n53142 , n53179 );
xor ( n53181 , n53133 , n53180 );
xor ( n53182 , n53124 , n53181 );
xor ( n53183 , n53115 , n53182 );
xor ( n53184 , n53106 , n53183 );
and ( n53185 , n52106 , n52181 );
and ( n53186 , n52181 , n52221 );
and ( n53187 , n52106 , n52221 );
or ( n53188 , n53185 , n53186 , n53187 );
and ( n53189 , n51997 , n52065 );
and ( n53190 , n52065 , n52102 );
and ( n53191 , n51997 , n52102 );
or ( n53192 , n53189 , n53190 , n53191 );
and ( n53193 , n52110 , n52111 );
and ( n53194 , n52111 , n52180 );
and ( n53195 , n52110 , n52180 );
or ( n53196 , n53193 , n53194 , n53195 );
xor ( n53197 , n53192 , n53196 );
and ( n53198 , n52070 , n52074 );
and ( n53199 , n52074 , n52101 );
and ( n53200 , n52070 , n52101 );
or ( n53201 , n53198 , n53199 , n53200 );
and ( n53202 , n52031 , n52047 );
and ( n53203 , n52047 , n52063 );
and ( n53204 , n52031 , n52063 );
or ( n53205 , n53202 , n53203 , n53204 );
and ( n53206 , n52014 , n52018 );
and ( n53207 , n52018 , n52024 );
and ( n53208 , n52014 , n52024 );
or ( n53209 , n53206 , n53207 , n53208 );
and ( n53210 , n52035 , n52040 );
and ( n53211 , n52040 , n52046 );
and ( n53212 , n52035 , n52046 );
or ( n53213 , n53210 , n53211 , n53212 );
xor ( n53214 , n53209 , n53213 );
and ( n53215 , n52020 , n52021 );
and ( n53216 , n52021 , n52023 );
and ( n53217 , n52020 , n52023 );
or ( n53218 , n53215 , n53216 , n53217 );
and ( n53219 , n52036 , n52037 );
and ( n53220 , n52037 , n52039 );
and ( n53221 , n52036 , n52039 );
or ( n53222 , n53219 , n53220 , n53221 );
xor ( n53223 , n53218 , n53222 );
and ( n53224 , n21216 , n5408 );
and ( n53225 , n22186 , n5103 );
xor ( n53226 , n53224 , n53225 );
and ( n53227 , n22892 , n4730 );
xor ( n53228 , n53226 , n53227 );
xor ( n53229 , n53223 , n53228 );
xor ( n53230 , n53214 , n53229 );
xor ( n53231 , n53205 , n53230 );
and ( n53232 , n52052 , n52056 );
and ( n53233 , n52056 , n52062 );
and ( n53234 , n52052 , n52062 );
or ( n53235 , n53232 , n53233 , n53234 );
and ( n53236 , n52042 , n52043 );
and ( n53237 , n52043 , n52045 );
and ( n53238 , n52042 , n52045 );
or ( n53239 , n53236 , n53237 , n53238 );
and ( n53240 , n18144 , n6504 );
and ( n53241 , n19324 , n6132 );
xor ( n53242 , n53240 , n53241 );
and ( n53243 , n20233 , n5765 );
xor ( n53244 , n53242 , n53243 );
xor ( n53245 , n53239 , n53244 );
and ( n53246 , n15758 , n7662 );
and ( n53247 , n16637 , n7310 );
xor ( n53248 , n53246 , n53247 );
and ( n53249 , n17512 , n6971 );
xor ( n53250 , n53248 , n53249 );
xor ( n53251 , n53245 , n53250 );
xor ( n53252 , n53235 , n53251 );
and ( n53253 , n52058 , n52059 );
and ( n53254 , n52059 , n52061 );
and ( n53255 , n52058 , n52061 );
or ( n53256 , n53253 , n53254 , n53255 );
and ( n53257 , n52089 , n52090 );
and ( n53258 , n52090 , n52092 );
and ( n53259 , n52089 , n52092 );
or ( n53260 , n53257 , n53258 , n53259 );
xor ( n53261 , n53256 , n53260 );
and ( n53262 , n13322 , n9348 );
and ( n53263 , n14118 , n8669 );
xor ( n53264 , n53262 , n53263 );
and ( n53265 , n14938 , n8243 );
xor ( n53266 , n53264 , n53265 );
xor ( n53267 , n53261 , n53266 );
xor ( n53268 , n53252 , n53267 );
xor ( n53269 , n53231 , n53268 );
xor ( n53270 , n53201 , n53269 );
and ( n53271 , n52079 , n52083 );
and ( n53272 , n52083 , n52100 );
and ( n53273 , n52079 , n52100 );
or ( n53274 , n53271 , n53272 , n53273 );
and ( n53275 , n52120 , n52135 );
and ( n53276 , n52135 , n52152 );
and ( n53277 , n52120 , n52152 );
or ( n53278 , n53275 , n53276 , n53277 );
xor ( n53279 , n53274 , n53278 );
and ( n53280 , n52088 , n52093 );
and ( n53281 , n52093 , n52099 );
and ( n53282 , n52088 , n52099 );
or ( n53283 , n53280 , n53281 , n53282 );
and ( n53284 , n52124 , n52128 );
and ( n53285 , n52128 , n52134 );
and ( n53286 , n52124 , n52134 );
or ( n53287 , n53284 , n53285 , n53286 );
xor ( n53288 , n53283 , n53287 );
and ( n53289 , n52095 , n52096 );
and ( n53290 , n52096 , n52098 );
and ( n53291 , n52095 , n52098 );
or ( n53292 , n53289 , n53290 , n53291 );
and ( n53293 , n12320 , n10239 );
buf ( n53294 , n53293 );
xor ( n53295 , n53292 , n53294 );
and ( n53296 , n8718 , n14044 );
and ( n53297 , n9400 , n13256 );
xor ( n53298 , n53296 , n53297 );
and ( n53299 , n10291 , n12531 );
xor ( n53300 , n53298 , n53299 );
xor ( n53301 , n53295 , n53300 );
xor ( n53302 , n53288 , n53301 );
xor ( n53303 , n53279 , n53302 );
xor ( n53304 , n53270 , n53303 );
xor ( n53305 , n53197 , n53304 );
xor ( n53306 , n53188 , n53305 );
and ( n53307 , n52116 , n52153 );
and ( n53308 , n52153 , n52179 );
and ( n53309 , n52116 , n52179 );
or ( n53310 , n53307 , n53308 , n53309 );
and ( n53311 , n52186 , n52220 );
xor ( n53312 , n53310 , n53311 );
and ( n53313 , n52158 , n52162 );
and ( n53314 , n52162 , n52178 );
and ( n53315 , n52158 , n52178 );
or ( n53316 , n53313 , n53314 , n53315 );
and ( n53317 , n52140 , n52145 );
and ( n53318 , n52145 , n52151 );
and ( n53319 , n52140 , n52151 );
or ( n53320 , n53317 , n53318 , n53319 );
and ( n53321 , n52130 , n52131 );
and ( n53322 , n52131 , n52133 );
and ( n53323 , n52130 , n52133 );
or ( n53324 , n53321 , n53322 , n53323 );
and ( n53325 , n52141 , n52142 );
and ( n53326 , n52142 , n52144 );
and ( n53327 , n52141 , n52144 );
or ( n53328 , n53325 , n53326 , n53327 );
xor ( n53329 , n53324 , n53328 );
and ( n53330 , n7385 , n16550 );
and ( n53331 , n7808 , n15691 );
xor ( n53332 , n53330 , n53331 );
and ( n53333 , n8079 , n14838 );
xor ( n53334 , n53332 , n53333 );
xor ( n53335 , n53329 , n53334 );
xor ( n53336 , n53320 , n53335 );
and ( n53337 , n52147 , n52148 );
and ( n53338 , n52148 , n52150 );
and ( n53339 , n52147 , n52150 );
or ( n53340 , n53337 , n53338 , n53339 );
and ( n53341 , n6187 , n19222 );
and ( n53342 , n6569 , n18407 );
xor ( n53343 , n53341 , n53342 );
and ( n53344 , n6816 , n17422 );
xor ( n53345 , n53343 , n53344 );
xor ( n53346 , n53340 , n53345 );
and ( n53347 , n4959 , n22065 );
and ( n53348 , n5459 , n20976 );
xor ( n53349 , n53347 , n53348 );
and ( n53350 , n5819 , n20156 );
xor ( n53351 , n53349 , n53350 );
xor ( n53352 , n53346 , n53351 );
xor ( n53353 , n53336 , n53352 );
xor ( n53354 , n53316 , n53353 );
and ( n53355 , n52167 , n52171 );
and ( n53356 , n52171 , n52177 );
and ( n53357 , n52167 , n52177 );
or ( n53358 , n53355 , n53356 , n53357 );
and ( n53359 , n52194 , n52199 );
and ( n53360 , n52199 , n52205 );
and ( n53361 , n52194 , n52205 );
or ( n53362 , n53359 , n53360 , n53361 );
xor ( n53363 , n53358 , n53362 );
and ( n53364 , n52173 , n52174 );
and ( n53365 , n52174 , n52176 );
and ( n53366 , n52173 , n52176 );
or ( n53367 , n53364 , n53365 , n53366 );
and ( n53368 , n52195 , n52196 );
and ( n53369 , n52196 , n52198 );
and ( n53370 , n52195 , n52198 );
or ( n53371 , n53368 , n53369 , n53370 );
xor ( n53372 , n53367 , n53371 );
and ( n53373 , n4132 , n25163 );
and ( n53374 , n4438 , n24137 );
xor ( n53375 , n53373 , n53374 );
and ( n53376 , n4766 , n23075 );
xor ( n53377 , n53375 , n53376 );
xor ( n53378 , n53372 , n53377 );
xor ( n53379 , n53363 , n53378 );
xor ( n53380 , n53354 , n53379 );
xor ( n53381 , n53312 , n53380 );
and ( n53382 , n52190 , n52206 );
and ( n53383 , n52206 , n52219 );
and ( n53384 , n52190 , n52219 );
or ( n53385 , n53382 , n53383 , n53384 );
and ( n53386 , n52211 , n52218 );
and ( n53387 , n52201 , n52202 );
and ( n53388 , n52202 , n52204 );
and ( n53389 , n52201 , n52204 );
or ( n53390 , n53387 , n53388 , n53389 );
and ( n53391 , n2462 , n31761 );
and ( n53392 , n2779 , n30629 );
xor ( n53393 , n53391 , n53392 );
and ( n53394 , n3024 , n29508 );
xor ( n53395 , n53393 , n53394 );
xor ( n53396 , n53390 , n53395 );
and ( n53397 , n3182 , n28406 );
and ( n53398 , n3545 , n27296 );
xor ( n53399 , n53397 , n53398 );
and ( n53400 , n3801 , n26216 );
xor ( n53401 , n53399 , n53400 );
xor ( n53402 , n53396 , n53401 );
xor ( n53403 , n53386 , n53402 );
and ( n53404 , n52214 , n52215 );
and ( n53405 , n52215 , n52217 );
and ( n53406 , n52214 , n52217 );
or ( n53407 , n53404 , n53405 , n53406 );
not ( n53408 , n2120 );
and ( n53409 , n34193 , n2120 );
nor ( n53410 , n53408 , n53409 );
and ( n53411 , n2324 , n32999 );
xor ( n53412 , n53410 , n53411 );
xor ( n53413 , n53407 , n53412 );
xor ( n53414 , n53403 , n53413 );
xor ( n53415 , n53385 , n53414 );
xor ( n53416 , n53381 , n53415 );
xor ( n53417 , n53306 , n53416 );
xor ( n53418 , n53184 , n53417 );
xor ( n53419 , n53102 , n53418 );
xor ( n53420 , n53093 , n53419 );
and ( n53421 , n51885 , n51888 );
and ( n53422 , n51888 , n52225 );
and ( n53423 , n51885 , n52225 );
or ( n53424 , n53421 , n53422 , n53423 );
xor ( n53425 , n53420 , n53424 );
and ( n53426 , n52226 , n52230 );
and ( n53427 , n52231 , n52234 );
or ( n53428 , n53426 , n53427 );
xor ( n53429 , n53425 , n53428 );
buf ( n53430 , n53429 );
buf ( n53431 , n53430 );
not ( n53432 , n53431 );
nor ( n53433 , n53432 , n8739 );
xor ( n53434 , n53085 , n53433 );
and ( n53435 , n51881 , n52239 );
and ( n53436 , n52240 , n52243 );
or ( n53437 , n53435 , n53436 );
xor ( n53438 , n53434 , n53437 );
buf ( n53439 , n53438 );
buf ( n53440 , n53439 );
not ( n53441 , n53440 );
buf ( n53442 , n578 );
not ( n53443 , n53442 );
nor ( n53444 , n53441 , n53443 );
xor ( n53445 , n52711 , n53444 );
xor ( n53446 , n52255 , n52708 );
nor ( n53447 , n52247 , n53443 );
and ( n53448 , n53446 , n53447 );
xor ( n53449 , n53446 , n53447 );
xor ( n53450 , n52259 , n52706 );
nor ( n53451 , n51049 , n53443 );
and ( n53452 , n53450 , n53451 );
xor ( n53453 , n53450 , n53451 );
xor ( n53454 , n52263 , n52704 );
nor ( n53455 , n49850 , n53443 );
and ( n53456 , n53454 , n53455 );
xor ( n53457 , n53454 , n53455 );
xor ( n53458 , n52267 , n52702 );
nor ( n53459 , n48650 , n53443 );
and ( n53460 , n53458 , n53459 );
xor ( n53461 , n53458 , n53459 );
xor ( n53462 , n52271 , n52700 );
nor ( n53463 , n47449 , n53443 );
and ( n53464 , n53462 , n53463 );
xor ( n53465 , n53462 , n53463 );
xor ( n53466 , n52275 , n52698 );
nor ( n53467 , n46248 , n53443 );
and ( n53468 , n53466 , n53467 );
xor ( n53469 , n53466 , n53467 );
xor ( n53470 , n52279 , n52696 );
nor ( n53471 , n45047 , n53443 );
and ( n53472 , n53470 , n53471 );
xor ( n53473 , n53470 , n53471 );
xor ( n53474 , n52283 , n52694 );
nor ( n53475 , n43843 , n53443 );
and ( n53476 , n53474 , n53475 );
xor ( n53477 , n53474 , n53475 );
xor ( n53478 , n52287 , n52692 );
nor ( n53479 , n42641 , n53443 );
and ( n53480 , n53478 , n53479 );
xor ( n53481 , n53478 , n53479 );
xor ( n53482 , n52291 , n52690 );
nor ( n53483 , n41437 , n53443 );
and ( n53484 , n53482 , n53483 );
xor ( n53485 , n53482 , n53483 );
xor ( n53486 , n52295 , n52688 );
nor ( n53487 , n40232 , n53443 );
and ( n53488 , n53486 , n53487 );
xor ( n53489 , n53486 , n53487 );
xor ( n53490 , n52299 , n52686 );
nor ( n53491 , n39027 , n53443 );
and ( n53492 , n53490 , n53491 );
xor ( n53493 , n53490 , n53491 );
xor ( n53494 , n52303 , n52684 );
nor ( n53495 , n37825 , n53443 );
and ( n53496 , n53494 , n53495 );
xor ( n53497 , n53494 , n53495 );
xor ( n53498 , n52307 , n52682 );
nor ( n53499 , n36620 , n53443 );
and ( n53500 , n53498 , n53499 );
xor ( n53501 , n53498 , n53499 );
xor ( n53502 , n52311 , n52680 );
nor ( n53503 , n35419 , n53443 );
and ( n53504 , n53502 , n53503 );
xor ( n53505 , n53502 , n53503 );
xor ( n53506 , n52315 , n52678 );
nor ( n53507 , n34224 , n53443 );
and ( n53508 , n53506 , n53507 );
xor ( n53509 , n53506 , n53507 );
xor ( n53510 , n52319 , n52676 );
nor ( n53511 , n33033 , n53443 );
and ( n53512 , n53510 , n53511 );
xor ( n53513 , n53510 , n53511 );
xor ( n53514 , n52323 , n52674 );
nor ( n53515 , n31867 , n53443 );
and ( n53516 , n53514 , n53515 );
xor ( n53517 , n53514 , n53515 );
xor ( n53518 , n52327 , n52672 );
nor ( n53519 , n30725 , n53443 );
and ( n53520 , n53518 , n53519 );
xor ( n53521 , n53518 , n53519 );
xor ( n53522 , n52331 , n52670 );
nor ( n53523 , n29596 , n53443 );
and ( n53524 , n53522 , n53523 );
xor ( n53525 , n53522 , n53523 );
xor ( n53526 , n52335 , n52668 );
nor ( n53527 , n28487 , n53443 );
and ( n53528 , n53526 , n53527 );
xor ( n53529 , n53526 , n53527 );
xor ( n53530 , n52339 , n52666 );
nor ( n53531 , n27397 , n53443 );
and ( n53532 , n53530 , n53531 );
xor ( n53533 , n53530 , n53531 );
xor ( n53534 , n52343 , n52664 );
nor ( n53535 , n26326 , n53443 );
and ( n53536 , n53534 , n53535 );
xor ( n53537 , n53534 , n53535 );
xor ( n53538 , n52347 , n52662 );
nor ( n53539 , n25272 , n53443 );
and ( n53540 , n53538 , n53539 );
xor ( n53541 , n53538 , n53539 );
xor ( n53542 , n52351 , n52660 );
nor ( n53543 , n24242 , n53443 );
and ( n53544 , n53542 , n53543 );
xor ( n53545 , n53542 , n53543 );
xor ( n53546 , n52355 , n52658 );
nor ( n53547 , n23225 , n53443 );
and ( n53548 , n53546 , n53547 );
xor ( n53549 , n53546 , n53547 );
xor ( n53550 , n52359 , n52656 );
nor ( n53551 , n22231 , n53443 );
and ( n53552 , n53550 , n53551 );
xor ( n53553 , n53550 , n53551 );
xor ( n53554 , n52363 , n52654 );
nor ( n53555 , n21258 , n53443 );
and ( n53556 , n53554 , n53555 );
xor ( n53557 , n53554 , n53555 );
xor ( n53558 , n52367 , n52652 );
nor ( n53559 , n20303 , n53443 );
and ( n53560 , n53558 , n53559 );
xor ( n53561 , n53558 , n53559 );
xor ( n53562 , n52371 , n52650 );
nor ( n53563 , n19365 , n53443 );
and ( n53564 , n53562 , n53563 );
xor ( n53565 , n53562 , n53563 );
xor ( n53566 , n52375 , n52648 );
nor ( n53567 , n18448 , n53443 );
and ( n53568 , n53566 , n53567 );
xor ( n53569 , n53566 , n53567 );
xor ( n53570 , n52379 , n52646 );
nor ( n53571 , n17548 , n53443 );
and ( n53572 , n53570 , n53571 );
xor ( n53573 , n53570 , n53571 );
xor ( n53574 , n52383 , n52644 );
nor ( n53575 , n16669 , n53443 );
and ( n53576 , n53574 , n53575 );
xor ( n53577 , n53574 , n53575 );
xor ( n53578 , n52387 , n52642 );
nor ( n53579 , n15809 , n53443 );
and ( n53580 , n53578 , n53579 );
xor ( n53581 , n53578 , n53579 );
xor ( n53582 , n52391 , n52640 );
nor ( n53583 , n14968 , n53443 );
and ( n53584 , n53582 , n53583 );
xor ( n53585 , n53582 , n53583 );
xor ( n53586 , n52395 , n52638 );
nor ( n53587 , n14147 , n53443 );
and ( n53588 , n53586 , n53587 );
xor ( n53589 , n53586 , n53587 );
xor ( n53590 , n52399 , n52636 );
nor ( n53591 , n13349 , n53443 );
and ( n53592 , n53590 , n53591 );
xor ( n53593 , n53590 , n53591 );
xor ( n53594 , n52403 , n52634 );
nor ( n53595 , n12564 , n53443 );
and ( n53596 , n53594 , n53595 );
xor ( n53597 , n53594 , n53595 );
xor ( n53598 , n52407 , n52632 );
nor ( n53599 , n11799 , n53443 );
and ( n53600 , n53598 , n53599 );
xor ( n53601 , n53598 , n53599 );
xor ( n53602 , n52411 , n52630 );
nor ( n53603 , n11050 , n53443 );
and ( n53604 , n53602 , n53603 );
xor ( n53605 , n53602 , n53603 );
xor ( n53606 , n52415 , n52628 );
nor ( n53607 , n10321 , n53443 );
and ( n53608 , n53606 , n53607 );
xor ( n53609 , n53606 , n53607 );
xor ( n53610 , n52419 , n52626 );
nor ( n53611 , n9429 , n53443 );
and ( n53612 , n53610 , n53611 );
xor ( n53613 , n53610 , n53611 );
xor ( n53614 , n52423 , n52624 );
nor ( n53615 , n8949 , n53443 );
and ( n53616 , n53614 , n53615 );
xor ( n53617 , n53614 , n53615 );
xor ( n53618 , n52427 , n52622 );
nor ( n53619 , n9437 , n53443 );
and ( n53620 , n53618 , n53619 );
xor ( n53621 , n53618 , n53619 );
xor ( n53622 , n52431 , n52620 );
nor ( n53623 , n9446 , n53443 );
and ( n53624 , n53622 , n53623 );
xor ( n53625 , n53622 , n53623 );
xor ( n53626 , n52435 , n52618 );
nor ( n53627 , n9455 , n53443 );
and ( n53628 , n53626 , n53627 );
xor ( n53629 , n53626 , n53627 );
xor ( n53630 , n52439 , n52616 );
nor ( n53631 , n9464 , n53443 );
and ( n53632 , n53630 , n53631 );
xor ( n53633 , n53630 , n53631 );
xor ( n53634 , n52443 , n52614 );
nor ( n53635 , n9473 , n53443 );
and ( n53636 , n53634 , n53635 );
xor ( n53637 , n53634 , n53635 );
xor ( n53638 , n52447 , n52612 );
nor ( n53639 , n9482 , n53443 );
and ( n53640 , n53638 , n53639 );
xor ( n53641 , n53638 , n53639 );
xor ( n53642 , n52451 , n52610 );
nor ( n53643 , n9491 , n53443 );
and ( n53644 , n53642 , n53643 );
xor ( n53645 , n53642 , n53643 );
xor ( n53646 , n52455 , n52608 );
nor ( n53647 , n9500 , n53443 );
and ( n53648 , n53646 , n53647 );
xor ( n53649 , n53646 , n53647 );
xor ( n53650 , n52459 , n52606 );
nor ( n53651 , n9509 , n53443 );
and ( n53652 , n53650 , n53651 );
xor ( n53653 , n53650 , n53651 );
xor ( n53654 , n52463 , n52604 );
nor ( n53655 , n9518 , n53443 );
and ( n53656 , n53654 , n53655 );
xor ( n53657 , n53654 , n53655 );
xor ( n53658 , n52467 , n52602 );
nor ( n53659 , n9527 , n53443 );
and ( n53660 , n53658 , n53659 );
xor ( n53661 , n53658 , n53659 );
xor ( n53662 , n52471 , n52600 );
nor ( n53663 , n9536 , n53443 );
and ( n53664 , n53662 , n53663 );
xor ( n53665 , n53662 , n53663 );
xor ( n53666 , n52475 , n52598 );
nor ( n53667 , n9545 , n53443 );
and ( n53668 , n53666 , n53667 );
xor ( n53669 , n53666 , n53667 );
xor ( n53670 , n52479 , n52596 );
nor ( n53671 , n9554 , n53443 );
and ( n53672 , n53670 , n53671 );
xor ( n53673 , n53670 , n53671 );
xor ( n53674 , n52483 , n52594 );
nor ( n53675 , n9563 , n53443 );
and ( n53676 , n53674 , n53675 );
xor ( n53677 , n53674 , n53675 );
xor ( n53678 , n52487 , n52592 );
nor ( n53679 , n9572 , n53443 );
and ( n53680 , n53678 , n53679 );
xor ( n53681 , n53678 , n53679 );
xor ( n53682 , n52491 , n52590 );
nor ( n53683 , n9581 , n53443 );
and ( n53684 , n53682 , n53683 );
xor ( n53685 , n53682 , n53683 );
xor ( n53686 , n52495 , n52588 );
nor ( n53687 , n9590 , n53443 );
and ( n53688 , n53686 , n53687 );
xor ( n53689 , n53686 , n53687 );
xor ( n53690 , n52499 , n52586 );
nor ( n53691 , n9599 , n53443 );
and ( n53692 , n53690 , n53691 );
xor ( n53693 , n53690 , n53691 );
xor ( n53694 , n52503 , n52584 );
nor ( n53695 , n9608 , n53443 );
and ( n53696 , n53694 , n53695 );
xor ( n53697 , n53694 , n53695 );
xor ( n53698 , n52507 , n52582 );
nor ( n53699 , n9617 , n53443 );
and ( n53700 , n53698 , n53699 );
xor ( n53701 , n53698 , n53699 );
xor ( n53702 , n52511 , n52580 );
nor ( n53703 , n9626 , n53443 );
and ( n53704 , n53702 , n53703 );
xor ( n53705 , n53702 , n53703 );
xor ( n53706 , n52515 , n52578 );
nor ( n53707 , n9635 , n53443 );
and ( n53708 , n53706 , n53707 );
xor ( n53709 , n53706 , n53707 );
xor ( n53710 , n52519 , n52576 );
nor ( n53711 , n9644 , n53443 );
and ( n53712 , n53710 , n53711 );
xor ( n53713 , n53710 , n53711 );
xor ( n53714 , n52523 , n52574 );
nor ( n53715 , n9653 , n53443 );
and ( n53716 , n53714 , n53715 );
xor ( n53717 , n53714 , n53715 );
xor ( n53718 , n52527 , n52572 );
nor ( n53719 , n9662 , n53443 );
and ( n53720 , n53718 , n53719 );
xor ( n53721 , n53718 , n53719 );
xor ( n53722 , n52531 , n52570 );
nor ( n53723 , n9671 , n53443 );
and ( n53724 , n53722 , n53723 );
xor ( n53725 , n53722 , n53723 );
xor ( n53726 , n52535 , n52568 );
nor ( n53727 , n9680 , n53443 );
and ( n53728 , n53726 , n53727 );
xor ( n53729 , n53726 , n53727 );
xor ( n53730 , n52539 , n52566 );
nor ( n53731 , n9689 , n53443 );
and ( n53732 , n53730 , n53731 );
xor ( n53733 , n53730 , n53731 );
xor ( n53734 , n52543 , n52564 );
nor ( n53735 , n9698 , n53443 );
and ( n53736 , n53734 , n53735 );
xor ( n53737 , n53734 , n53735 );
xor ( n53738 , n52547 , n52562 );
nor ( n53739 , n9707 , n53443 );
and ( n53740 , n53738 , n53739 );
xor ( n53741 , n53738 , n53739 );
xor ( n53742 , n52551 , n52560 );
nor ( n53743 , n9716 , n53443 );
and ( n53744 , n53742 , n53743 );
xor ( n53745 , n53742 , n53743 );
xor ( n53746 , n52555 , n52558 );
nor ( n53747 , n9725 , n53443 );
and ( n53748 , n53746 , n53747 );
xor ( n53749 , n53746 , n53747 );
xor ( n53750 , n52556 , n52557 );
nor ( n53751 , n9734 , n53443 );
and ( n53752 , n53750 , n53751 );
xor ( n53753 , n53750 , n53751 );
nor ( n53754 , n9752 , n52249 );
nor ( n53755 , n9743 , n53443 );
and ( n53756 , n53754 , n53755 );
and ( n53757 , n53753 , n53756 );
or ( n53758 , n53752 , n53757 );
and ( n53759 , n53749 , n53758 );
or ( n53760 , n53748 , n53759 );
and ( n53761 , n53745 , n53760 );
or ( n53762 , n53744 , n53761 );
and ( n53763 , n53741 , n53762 );
or ( n53764 , n53740 , n53763 );
and ( n53765 , n53737 , n53764 );
or ( n53766 , n53736 , n53765 );
and ( n53767 , n53733 , n53766 );
or ( n53768 , n53732 , n53767 );
and ( n53769 , n53729 , n53768 );
or ( n53770 , n53728 , n53769 );
and ( n53771 , n53725 , n53770 );
or ( n53772 , n53724 , n53771 );
and ( n53773 , n53721 , n53772 );
or ( n53774 , n53720 , n53773 );
and ( n53775 , n53717 , n53774 );
or ( n53776 , n53716 , n53775 );
and ( n53777 , n53713 , n53776 );
or ( n53778 , n53712 , n53777 );
and ( n53779 , n53709 , n53778 );
or ( n53780 , n53708 , n53779 );
and ( n53781 , n53705 , n53780 );
or ( n53782 , n53704 , n53781 );
and ( n53783 , n53701 , n53782 );
or ( n53784 , n53700 , n53783 );
and ( n53785 , n53697 , n53784 );
or ( n53786 , n53696 , n53785 );
and ( n53787 , n53693 , n53786 );
or ( n53788 , n53692 , n53787 );
and ( n53789 , n53689 , n53788 );
or ( n53790 , n53688 , n53789 );
and ( n53791 , n53685 , n53790 );
or ( n53792 , n53684 , n53791 );
and ( n53793 , n53681 , n53792 );
or ( n53794 , n53680 , n53793 );
and ( n53795 , n53677 , n53794 );
or ( n53796 , n53676 , n53795 );
and ( n53797 , n53673 , n53796 );
or ( n53798 , n53672 , n53797 );
and ( n53799 , n53669 , n53798 );
or ( n53800 , n53668 , n53799 );
and ( n53801 , n53665 , n53800 );
or ( n53802 , n53664 , n53801 );
and ( n53803 , n53661 , n53802 );
or ( n53804 , n53660 , n53803 );
and ( n53805 , n53657 , n53804 );
or ( n53806 , n53656 , n53805 );
and ( n53807 , n53653 , n53806 );
or ( n53808 , n53652 , n53807 );
and ( n53809 , n53649 , n53808 );
or ( n53810 , n53648 , n53809 );
and ( n53811 , n53645 , n53810 );
or ( n53812 , n53644 , n53811 );
and ( n53813 , n53641 , n53812 );
or ( n53814 , n53640 , n53813 );
and ( n53815 , n53637 , n53814 );
or ( n53816 , n53636 , n53815 );
and ( n53817 , n53633 , n53816 );
or ( n53818 , n53632 , n53817 );
and ( n53819 , n53629 , n53818 );
or ( n53820 , n53628 , n53819 );
and ( n53821 , n53625 , n53820 );
or ( n53822 , n53624 , n53821 );
and ( n53823 , n53621 , n53822 );
or ( n53824 , n53620 , n53823 );
and ( n53825 , n53617 , n53824 );
or ( n53826 , n53616 , n53825 );
and ( n53827 , n53613 , n53826 );
or ( n53828 , n53612 , n53827 );
and ( n53829 , n53609 , n53828 );
or ( n53830 , n53608 , n53829 );
and ( n53831 , n53605 , n53830 );
or ( n53832 , n53604 , n53831 );
and ( n53833 , n53601 , n53832 );
or ( n53834 , n53600 , n53833 );
and ( n53835 , n53597 , n53834 );
or ( n53836 , n53596 , n53835 );
and ( n53837 , n53593 , n53836 );
or ( n53838 , n53592 , n53837 );
and ( n53839 , n53589 , n53838 );
or ( n53840 , n53588 , n53839 );
and ( n53841 , n53585 , n53840 );
or ( n53842 , n53584 , n53841 );
and ( n53843 , n53581 , n53842 );
or ( n53844 , n53580 , n53843 );
and ( n53845 , n53577 , n53844 );
or ( n53846 , n53576 , n53845 );
and ( n53847 , n53573 , n53846 );
or ( n53848 , n53572 , n53847 );
and ( n53849 , n53569 , n53848 );
or ( n53850 , n53568 , n53849 );
and ( n53851 , n53565 , n53850 );
or ( n53852 , n53564 , n53851 );
and ( n53853 , n53561 , n53852 );
or ( n53854 , n53560 , n53853 );
and ( n53855 , n53557 , n53854 );
or ( n53856 , n53556 , n53855 );
and ( n53857 , n53553 , n53856 );
or ( n53858 , n53552 , n53857 );
and ( n53859 , n53549 , n53858 );
or ( n53860 , n53548 , n53859 );
and ( n53861 , n53545 , n53860 );
or ( n53862 , n53544 , n53861 );
and ( n53863 , n53541 , n53862 );
or ( n53864 , n53540 , n53863 );
and ( n53865 , n53537 , n53864 );
or ( n53866 , n53536 , n53865 );
and ( n53867 , n53533 , n53866 );
or ( n53868 , n53532 , n53867 );
and ( n53869 , n53529 , n53868 );
or ( n53870 , n53528 , n53869 );
and ( n53871 , n53525 , n53870 );
or ( n53872 , n53524 , n53871 );
and ( n53873 , n53521 , n53872 );
or ( n53874 , n53520 , n53873 );
and ( n53875 , n53517 , n53874 );
or ( n53876 , n53516 , n53875 );
and ( n53877 , n53513 , n53876 );
or ( n53878 , n53512 , n53877 );
and ( n53879 , n53509 , n53878 );
or ( n53880 , n53508 , n53879 );
and ( n53881 , n53505 , n53880 );
or ( n53882 , n53504 , n53881 );
and ( n53883 , n53501 , n53882 );
or ( n53884 , n53500 , n53883 );
and ( n53885 , n53497 , n53884 );
or ( n53886 , n53496 , n53885 );
and ( n53887 , n53493 , n53886 );
or ( n53888 , n53492 , n53887 );
and ( n53889 , n53489 , n53888 );
or ( n53890 , n53488 , n53889 );
and ( n53891 , n53485 , n53890 );
or ( n53892 , n53484 , n53891 );
and ( n53893 , n53481 , n53892 );
or ( n53894 , n53480 , n53893 );
and ( n53895 , n53477 , n53894 );
or ( n53896 , n53476 , n53895 );
and ( n53897 , n53473 , n53896 );
or ( n53898 , n53472 , n53897 );
and ( n53899 , n53469 , n53898 );
or ( n53900 , n53468 , n53899 );
and ( n53901 , n53465 , n53900 );
or ( n53902 , n53464 , n53901 );
and ( n53903 , n53461 , n53902 );
or ( n53904 , n53460 , n53903 );
and ( n53905 , n53457 , n53904 );
or ( n53906 , n53456 , n53905 );
and ( n53907 , n53453 , n53906 );
or ( n53908 , n53452 , n53907 );
and ( n53909 , n53449 , n53908 );
or ( n53910 , n53448 , n53909 );
xor ( n53911 , n53445 , n53910 );
and ( n53912 , n33403 , n2342 );
nor ( n53913 , n2343 , n53912 );
nor ( n53914 , n2566 , n32231 );
xor ( n53915 , n53913 , n53914 );
and ( n53916 , n52713 , n52714 );
and ( n53917 , n52715 , n52718 );
or ( n53918 , n53916 , n53917 );
xor ( n53919 , n53915 , n53918 );
nor ( n53920 , n2797 , n31083 );
xor ( n53921 , n53919 , n53920 );
and ( n53922 , n52719 , n52720 );
and ( n53923 , n52721 , n52724 );
or ( n53924 , n53922 , n53923 );
xor ( n53925 , n53921 , n53924 );
nor ( n53926 , n3043 , n29948 );
xor ( n53927 , n53925 , n53926 );
and ( n53928 , n52725 , n52726 );
and ( n53929 , n52727 , n52730 );
or ( n53930 , n53928 , n53929 );
xor ( n53931 , n53927 , n53930 );
nor ( n53932 , n3300 , n28833 );
xor ( n53933 , n53931 , n53932 );
and ( n53934 , n52731 , n52732 );
and ( n53935 , n52733 , n52736 );
or ( n53936 , n53934 , n53935 );
xor ( n53937 , n53933 , n53936 );
nor ( n53938 , n3570 , n27737 );
xor ( n53939 , n53937 , n53938 );
and ( n53940 , n52737 , n52738 );
and ( n53941 , n52739 , n52742 );
or ( n53942 , n53940 , n53941 );
xor ( n53943 , n53939 , n53942 );
nor ( n53944 , n3853 , n26660 );
xor ( n53945 , n53943 , n53944 );
and ( n53946 , n52743 , n52744 );
and ( n53947 , n52745 , n52748 );
or ( n53948 , n53946 , n53947 );
xor ( n53949 , n53945 , n53948 );
nor ( n53950 , n4151 , n25600 );
xor ( n53951 , n53949 , n53950 );
and ( n53952 , n52749 , n52750 );
and ( n53953 , n52751 , n52754 );
or ( n53954 , n53952 , n53953 );
xor ( n53955 , n53951 , n53954 );
nor ( n53956 , n4458 , n24564 );
xor ( n53957 , n53955 , n53956 );
and ( n53958 , n52755 , n52756 );
and ( n53959 , n52757 , n52760 );
or ( n53960 , n53958 , n53959 );
xor ( n53961 , n53957 , n53960 );
nor ( n53962 , n4786 , n23541 );
xor ( n53963 , n53961 , n53962 );
and ( n53964 , n52761 , n52762 );
and ( n53965 , n52763 , n52766 );
or ( n53966 , n53964 , n53965 );
xor ( n53967 , n53963 , n53966 );
nor ( n53968 , n5126 , n22541 );
xor ( n53969 , n53967 , n53968 );
and ( n53970 , n52767 , n52768 );
and ( n53971 , n52769 , n52772 );
or ( n53972 , n53970 , n53971 );
xor ( n53973 , n53969 , n53972 );
nor ( n53974 , n5477 , n21562 );
xor ( n53975 , n53973 , n53974 );
and ( n53976 , n52773 , n52774 );
and ( n53977 , n52775 , n52778 );
or ( n53978 , n53976 , n53977 );
xor ( n53979 , n53975 , n53978 );
nor ( n53980 , n5838 , n20601 );
xor ( n53981 , n53979 , n53980 );
and ( n53982 , n52779 , n52780 );
and ( n53983 , n52781 , n52784 );
or ( n53984 , n53982 , n53983 );
xor ( n53985 , n53981 , n53984 );
nor ( n53986 , n6212 , n19657 );
xor ( n53987 , n53985 , n53986 );
and ( n53988 , n52785 , n52786 );
and ( n53989 , n52787 , n52790 );
or ( n53990 , n53988 , n53989 );
xor ( n53991 , n53987 , n53990 );
nor ( n53992 , n6596 , n18734 );
xor ( n53993 , n53991 , n53992 );
and ( n53994 , n52791 , n52792 );
and ( n53995 , n52793 , n52796 );
or ( n53996 , n53994 , n53995 );
xor ( n53997 , n53993 , n53996 );
nor ( n53998 , n6997 , n17828 );
xor ( n53999 , n53997 , n53998 );
and ( n54000 , n52797 , n52798 );
and ( n54001 , n52799 , n52802 );
or ( n54002 , n54000 , n54001 );
xor ( n54003 , n53999 , n54002 );
nor ( n54004 , n7413 , n16943 );
xor ( n54005 , n54003 , n54004 );
and ( n54006 , n52803 , n52804 );
and ( n54007 , n52805 , n52808 );
or ( n54008 , n54006 , n54007 );
xor ( n54009 , n54005 , n54008 );
nor ( n54010 , n7841 , n16077 );
xor ( n54011 , n54009 , n54010 );
and ( n54012 , n52809 , n52810 );
and ( n54013 , n52811 , n52814 );
or ( n54014 , n54012 , n54013 );
xor ( n54015 , n54011 , n54014 );
nor ( n54016 , n8281 , n15230 );
xor ( n54017 , n54015 , n54016 );
and ( n54018 , n52815 , n52816 );
and ( n54019 , n52817 , n52820 );
or ( n54020 , n54018 , n54019 );
xor ( n54021 , n54017 , n54020 );
nor ( n54022 , n8737 , n14403 );
xor ( n54023 , n54021 , n54022 );
and ( n54024 , n52821 , n52822 );
and ( n54025 , n52823 , n52826 );
or ( n54026 , n54024 , n54025 );
xor ( n54027 , n54023 , n54026 );
nor ( n54028 , n9420 , n13599 );
xor ( n54029 , n54027 , n54028 );
and ( n54030 , n52827 , n52828 );
and ( n54031 , n52829 , n52832 );
or ( n54032 , n54030 , n54031 );
xor ( n54033 , n54029 , n54032 );
nor ( n54034 , n10312 , n12808 );
xor ( n54035 , n54033 , n54034 );
and ( n54036 , n52833 , n52834 );
and ( n54037 , n52835 , n52838 );
or ( n54038 , n54036 , n54037 );
xor ( n54039 , n54035 , n54038 );
nor ( n54040 , n11041 , n12037 );
xor ( n54041 , n54039 , n54040 );
and ( n54042 , n52839 , n52840 );
and ( n54043 , n52841 , n52844 );
or ( n54044 , n54042 , n54043 );
xor ( n54045 , n54041 , n54044 );
nor ( n54046 , n11790 , n11282 );
xor ( n54047 , n54045 , n54046 );
and ( n54048 , n52845 , n52846 );
and ( n54049 , n52847 , n52850 );
or ( n54050 , n54048 , n54049 );
xor ( n54051 , n54047 , n54050 );
nor ( n54052 , n12555 , n10547 );
xor ( n54053 , n54051 , n54052 );
and ( n54054 , n52851 , n52852 );
and ( n54055 , n52853 , n52856 );
or ( n54056 , n54054 , n54055 );
xor ( n54057 , n54053 , n54056 );
nor ( n54058 , n13340 , n9829 );
xor ( n54059 , n54057 , n54058 );
and ( n54060 , n52857 , n52858 );
and ( n54061 , n52859 , n52862 );
or ( n54062 , n54060 , n54061 );
xor ( n54063 , n54059 , n54062 );
nor ( n54064 , n14138 , n8955 );
xor ( n54065 , n54063 , n54064 );
and ( n54066 , n52863 , n52864 );
and ( n54067 , n52865 , n52868 );
or ( n54068 , n54066 , n54067 );
xor ( n54069 , n54065 , n54068 );
nor ( n54070 , n14959 , n603 );
xor ( n54071 , n54069 , n54070 );
and ( n54072 , n52869 , n52870 );
and ( n54073 , n52871 , n52874 );
or ( n54074 , n54072 , n54073 );
xor ( n54075 , n54071 , n54074 );
nor ( n54076 , n15800 , n652 );
xor ( n54077 , n54075 , n54076 );
and ( n54078 , n52875 , n52876 );
and ( n54079 , n52877 , n52880 );
or ( n54080 , n54078 , n54079 );
xor ( n54081 , n54077 , n54080 );
nor ( n54082 , n16660 , n624 );
xor ( n54083 , n54081 , n54082 );
and ( n54084 , n52881 , n52882 );
and ( n54085 , n52883 , n52886 );
or ( n54086 , n54084 , n54085 );
xor ( n54087 , n54083 , n54086 );
nor ( n54088 , n17539 , n648 );
xor ( n54089 , n54087 , n54088 );
and ( n54090 , n52887 , n52888 );
and ( n54091 , n52889 , n52892 );
or ( n54092 , n54090 , n54091 );
xor ( n54093 , n54089 , n54092 );
nor ( n54094 , n18439 , n686 );
xor ( n54095 , n54093 , n54094 );
and ( n54096 , n52893 , n52894 );
and ( n54097 , n52895 , n52898 );
or ( n54098 , n54096 , n54097 );
xor ( n54099 , n54095 , n54098 );
nor ( n54100 , n19356 , n735 );
xor ( n54101 , n54099 , n54100 );
and ( n54102 , n52899 , n52900 );
and ( n54103 , n52901 , n52904 );
or ( n54104 , n54102 , n54103 );
xor ( n54105 , n54101 , n54104 );
nor ( n54106 , n20294 , n798 );
xor ( n54107 , n54105 , n54106 );
and ( n54108 , n52905 , n52906 );
and ( n54109 , n52907 , n52910 );
or ( n54110 , n54108 , n54109 );
xor ( n54111 , n54107 , n54110 );
nor ( n54112 , n21249 , n870 );
xor ( n54113 , n54111 , n54112 );
and ( n54114 , n52911 , n52912 );
and ( n54115 , n52913 , n52916 );
or ( n54116 , n54114 , n54115 );
xor ( n54117 , n54113 , n54116 );
nor ( n54118 , n22222 , n960 );
xor ( n54119 , n54117 , n54118 );
and ( n54120 , n52917 , n52918 );
and ( n54121 , n52919 , n52922 );
or ( n54122 , n54120 , n54121 );
xor ( n54123 , n54119 , n54122 );
nor ( n54124 , n23216 , n1064 );
xor ( n54125 , n54123 , n54124 );
and ( n54126 , n52923 , n52924 );
and ( n54127 , n52925 , n52928 );
or ( n54128 , n54126 , n54127 );
xor ( n54129 , n54125 , n54128 );
nor ( n54130 , n24233 , n1178 );
xor ( n54131 , n54129 , n54130 );
and ( n54132 , n52929 , n52930 );
and ( n54133 , n52931 , n52934 );
or ( n54134 , n54132 , n54133 );
xor ( n54135 , n54131 , n54134 );
nor ( n54136 , n25263 , n1305 );
xor ( n54137 , n54135 , n54136 );
and ( n54138 , n52935 , n52936 );
and ( n54139 , n52937 , n52940 );
or ( n54140 , n54138 , n54139 );
xor ( n54141 , n54137 , n54140 );
nor ( n54142 , n26317 , n1447 );
xor ( n54143 , n54141 , n54142 );
and ( n54144 , n52941 , n52942 );
and ( n54145 , n52943 , n52946 );
or ( n54146 , n54144 , n54145 );
xor ( n54147 , n54143 , n54146 );
nor ( n54148 , n27388 , n1600 );
xor ( n54149 , n54147 , n54148 );
and ( n54150 , n52947 , n52948 );
and ( n54151 , n52949 , n52952 );
or ( n54152 , n54150 , n54151 );
xor ( n54153 , n54149 , n54152 );
nor ( n54154 , n28478 , n1768 );
xor ( n54155 , n54153 , n54154 );
and ( n54156 , n52953 , n52954 );
and ( n54157 , n52955 , n52958 );
or ( n54158 , n54156 , n54157 );
xor ( n54159 , n54155 , n54158 );
nor ( n54160 , n29587 , n1947 );
xor ( n54161 , n54159 , n54160 );
and ( n54162 , n52959 , n52960 );
and ( n54163 , n52961 , n52964 );
or ( n54164 , n54162 , n54163 );
xor ( n54165 , n54161 , n54164 );
nor ( n54166 , n30716 , n2139 );
xor ( n54167 , n54165 , n54166 );
and ( n54168 , n52965 , n52966 );
and ( n54169 , n52967 , n52970 );
or ( n54170 , n54168 , n54169 );
xor ( n54171 , n54167 , n54170 );
nor ( n54172 , n31858 , n2345 );
xor ( n54173 , n54171 , n54172 );
and ( n54174 , n52971 , n52972 );
and ( n54175 , n52973 , n52976 );
or ( n54176 , n54174 , n54175 );
xor ( n54177 , n54173 , n54176 );
nor ( n54178 , n33024 , n2568 );
xor ( n54179 , n54177 , n54178 );
and ( n54180 , n52977 , n52978 );
and ( n54181 , n52979 , n52982 );
or ( n54182 , n54180 , n54181 );
xor ( n54183 , n54179 , n54182 );
nor ( n54184 , n34215 , n2799 );
xor ( n54185 , n54183 , n54184 );
and ( n54186 , n52983 , n52984 );
and ( n54187 , n52985 , n52988 );
or ( n54188 , n54186 , n54187 );
xor ( n54189 , n54185 , n54188 );
nor ( n54190 , n35410 , n3045 );
xor ( n54191 , n54189 , n54190 );
and ( n54192 , n52989 , n52990 );
and ( n54193 , n52991 , n52994 );
or ( n54194 , n54192 , n54193 );
xor ( n54195 , n54191 , n54194 );
nor ( n54196 , n36611 , n3302 );
xor ( n54197 , n54195 , n54196 );
and ( n54198 , n52995 , n52996 );
and ( n54199 , n52997 , n53000 );
or ( n54200 , n54198 , n54199 );
xor ( n54201 , n54197 , n54200 );
nor ( n54202 , n37816 , n3572 );
xor ( n54203 , n54201 , n54202 );
and ( n54204 , n53001 , n53002 );
and ( n54205 , n53003 , n53006 );
or ( n54206 , n54204 , n54205 );
xor ( n54207 , n54203 , n54206 );
nor ( n54208 , n39018 , n3855 );
xor ( n54209 , n54207 , n54208 );
and ( n54210 , n53007 , n53008 );
and ( n54211 , n53009 , n53012 );
or ( n54212 , n54210 , n54211 );
xor ( n54213 , n54209 , n54212 );
nor ( n54214 , n40223 , n4153 );
xor ( n54215 , n54213 , n54214 );
and ( n54216 , n53013 , n53014 );
and ( n54217 , n53015 , n53018 );
or ( n54218 , n54216 , n54217 );
xor ( n54219 , n54215 , n54218 );
nor ( n54220 , n41428 , n4460 );
xor ( n54221 , n54219 , n54220 );
and ( n54222 , n53019 , n53020 );
and ( n54223 , n53021 , n53024 );
or ( n54224 , n54222 , n54223 );
xor ( n54225 , n54221 , n54224 );
nor ( n54226 , n42632 , n4788 );
xor ( n54227 , n54225 , n54226 );
and ( n54228 , n53025 , n53026 );
and ( n54229 , n53027 , n53030 );
or ( n54230 , n54228 , n54229 );
xor ( n54231 , n54227 , n54230 );
nor ( n54232 , n43834 , n5128 );
xor ( n54233 , n54231 , n54232 );
and ( n54234 , n53031 , n53032 );
and ( n54235 , n53033 , n53036 );
or ( n54236 , n54234 , n54235 );
xor ( n54237 , n54233 , n54236 );
nor ( n54238 , n45038 , n5479 );
xor ( n54239 , n54237 , n54238 );
and ( n54240 , n53037 , n53038 );
and ( n54241 , n53039 , n53042 );
or ( n54242 , n54240 , n54241 );
xor ( n54243 , n54239 , n54242 );
nor ( n54244 , n46239 , n5840 );
xor ( n54245 , n54243 , n54244 );
and ( n54246 , n53043 , n53044 );
and ( n54247 , n53045 , n53048 );
or ( n54248 , n54246 , n54247 );
xor ( n54249 , n54245 , n54248 );
nor ( n54250 , n47440 , n6214 );
xor ( n54251 , n54249 , n54250 );
and ( n54252 , n53049 , n53050 );
and ( n54253 , n53051 , n53054 );
or ( n54254 , n54252 , n54253 );
xor ( n54255 , n54251 , n54254 );
nor ( n54256 , n48641 , n6598 );
xor ( n54257 , n54255 , n54256 );
and ( n54258 , n53055 , n53056 );
and ( n54259 , n53057 , n53060 );
or ( n54260 , n54258 , n54259 );
xor ( n54261 , n54257 , n54260 );
nor ( n54262 , n49841 , n6999 );
xor ( n54263 , n54261 , n54262 );
and ( n54264 , n53061 , n53062 );
and ( n54265 , n53063 , n53066 );
or ( n54266 , n54264 , n54265 );
xor ( n54267 , n54263 , n54266 );
nor ( n54268 , n51040 , n7415 );
xor ( n54269 , n54267 , n54268 );
and ( n54270 , n53067 , n53068 );
and ( n54271 , n53069 , n53072 );
or ( n54272 , n54270 , n54271 );
xor ( n54273 , n54269 , n54272 );
nor ( n54274 , n52238 , n7843 );
xor ( n54275 , n54273 , n54274 );
and ( n54276 , n53073 , n53074 );
and ( n54277 , n53075 , n53078 );
or ( n54278 , n54276 , n54277 );
xor ( n54279 , n54275 , n54278 );
nor ( n54280 , n53432 , n8283 );
xor ( n54281 , n54279 , n54280 );
and ( n54282 , n53079 , n53080 );
and ( n54283 , n53081 , n53084 );
or ( n54284 , n54282 , n54283 );
xor ( n54285 , n54281 , n54284 );
and ( n54286 , n53097 , n53101 );
and ( n54287 , n53101 , n53418 );
and ( n54288 , n53097 , n53418 );
or ( n54289 , n54286 , n54287 , n54288 );
and ( n54290 , n33774 , n2298 );
not ( n54291 , n2298 );
nor ( n54292 , n54290 , n54291 );
xor ( n54293 , n54289 , n54292 );
and ( n54294 , n53110 , n53114 );
and ( n54295 , n53114 , n53182 );
and ( n54296 , n53110 , n53182 );
or ( n54297 , n54294 , n54295 , n54296 );
and ( n54298 , n53106 , n53183 );
and ( n54299 , n53183 , n53417 );
and ( n54300 , n53106 , n53417 );
or ( n54301 , n54298 , n54299 , n54300 );
xor ( n54302 , n54297 , n54301 );
and ( n54303 , n53188 , n53305 );
and ( n54304 , n53305 , n53416 );
and ( n54305 , n53188 , n53416 );
or ( n54306 , n54303 , n54304 , n54305 );
and ( n54307 , n53119 , n53123 );
and ( n54308 , n53123 , n53181 );
and ( n54309 , n53119 , n53181 );
or ( n54310 , n54307 , n54308 , n54309 );
and ( n54311 , n53192 , n53196 );
and ( n54312 , n53196 , n53304 );
and ( n54313 , n53192 , n53304 );
or ( n54314 , n54311 , n54312 , n54313 );
xor ( n54315 , n54310 , n54314 );
and ( n54316 , n53150 , n53154 );
and ( n54317 , n53154 , n53160 );
and ( n54318 , n53150 , n53160 );
or ( n54319 , n54316 , n54317 , n54318 );
and ( n54320 , n53128 , n53132 );
and ( n54321 , n53132 , n53180 );
and ( n54322 , n53128 , n53180 );
or ( n54323 , n54320 , n54321 , n54322 );
xor ( n54324 , n54319 , n54323 );
and ( n54325 , n53205 , n53230 );
and ( n54326 , n53230 , n53268 );
and ( n54327 , n53205 , n53268 );
or ( n54328 , n54325 , n54326 , n54327 );
and ( n54329 , n53137 , n53141 );
and ( n54330 , n53141 , n53179 );
and ( n54331 , n53137 , n53179 );
or ( n54332 , n54329 , n54330 , n54331 );
xor ( n54333 , n54328 , n54332 );
and ( n54334 , n53209 , n53213 );
and ( n54335 , n53213 , n53229 );
and ( n54336 , n53209 , n53229 );
or ( n54337 , n54334 , n54335 , n54336 );
and ( n54338 , n53146 , n53161 );
and ( n54339 , n53161 , n53178 );
and ( n54340 , n53146 , n53178 );
or ( n54341 , n54338 , n54339 , n54340 );
xor ( n54342 , n54337 , n54341 );
and ( n54343 , n53166 , n53171 );
and ( n54344 , n53171 , n53177 );
and ( n54345 , n53166 , n53177 );
or ( n54346 , n54343 , n54344 , n54345 );
and ( n54347 , n53156 , n53157 );
and ( n54348 , n53157 , n53159 );
and ( n54349 , n53156 , n53159 );
or ( n54350 , n54347 , n54348 , n54349 );
and ( n54351 , n53167 , n53168 );
and ( n54352 , n53168 , n53170 );
and ( n54353 , n53167 , n53170 );
or ( n54354 , n54351 , n54352 , n54353 );
xor ( n54355 , n54350 , n54354 );
and ( n54356 , n30695 , n2981 );
and ( n54357 , n31836 , n2739 );
xor ( n54358 , n54356 , n54357 );
and ( n54359 , n32649 , n2544 );
xor ( n54360 , n54358 , n54359 );
xor ( n54361 , n54355 , n54360 );
xor ( n54362 , n54346 , n54361 );
and ( n54363 , n53173 , n53174 );
and ( n54364 , n53174 , n53176 );
and ( n54365 , n53173 , n53176 );
or ( n54366 , n54363 , n54364 , n54365 );
and ( n54367 , n27361 , n3749 );
and ( n54368 , n28456 , n3495 );
xor ( n54369 , n54367 , n54368 );
and ( n54370 , n29559 , n3271 );
xor ( n54371 , n54369 , n54370 );
xor ( n54372 , n54366 , n54371 );
and ( n54373 , n24214 , n4730 );
and ( n54374 , n25243 , n4403 );
xor ( n54375 , n54373 , n54374 );
and ( n54376 , n26296 , n4102 );
xor ( n54377 , n54375 , n54376 );
xor ( n54378 , n54372 , n54377 );
xor ( n54379 , n54362 , n54378 );
xor ( n54380 , n54342 , n54379 );
xor ( n54381 , n54333 , n54380 );
xor ( n54382 , n54324 , n54381 );
xor ( n54383 , n54315 , n54382 );
xor ( n54384 , n54306 , n54383 );
and ( n54385 , n53381 , n53415 );
and ( n54386 , n53201 , n53269 );
and ( n54387 , n53269 , n53303 );
and ( n54388 , n53201 , n53303 );
or ( n54389 , n54386 , n54387 , n54388 );
and ( n54390 , n53310 , n53311 );
and ( n54391 , n53311 , n53380 );
and ( n54392 , n53310 , n53380 );
or ( n54393 , n54390 , n54391 , n54392 );
xor ( n54394 , n54389 , n54393 );
and ( n54395 , n53274 , n53278 );
and ( n54396 , n53278 , n53302 );
and ( n54397 , n53274 , n53302 );
or ( n54398 , n54395 , n54396 , n54397 );
and ( n54399 , n53235 , n53251 );
and ( n54400 , n53251 , n53267 );
and ( n54401 , n53235 , n53267 );
or ( n54402 , n54399 , n54400 , n54401 );
and ( n54403 , n53218 , n53222 );
and ( n54404 , n53222 , n53228 );
and ( n54405 , n53218 , n53228 );
or ( n54406 , n54403 , n54404 , n54405 );
and ( n54407 , n53239 , n53244 );
and ( n54408 , n53244 , n53250 );
and ( n54409 , n53239 , n53250 );
or ( n54410 , n54407 , n54408 , n54409 );
xor ( n54411 , n54406 , n54410 );
and ( n54412 , n53224 , n53225 );
and ( n54413 , n53225 , n53227 );
and ( n54414 , n53224 , n53227 );
or ( n54415 , n54412 , n54413 , n54414 );
and ( n54416 , n53240 , n53241 );
and ( n54417 , n53241 , n53243 );
and ( n54418 , n53240 , n53243 );
or ( n54419 , n54416 , n54417 , n54418 );
xor ( n54420 , n54415 , n54419 );
and ( n54421 , n21216 , n5765 );
and ( n54422 , n22186 , n5408 );
xor ( n54423 , n54421 , n54422 );
and ( n54424 , n22892 , n5103 );
xor ( n54425 , n54423 , n54424 );
xor ( n54426 , n54420 , n54425 );
xor ( n54427 , n54411 , n54426 );
xor ( n54428 , n54402 , n54427 );
and ( n54429 , n53256 , n53260 );
and ( n54430 , n53260 , n53266 );
and ( n54431 , n53256 , n53266 );
or ( n54432 , n54429 , n54430 , n54431 );
and ( n54433 , n53246 , n53247 );
and ( n54434 , n53247 , n53249 );
and ( n54435 , n53246 , n53249 );
or ( n54436 , n54433 , n54434 , n54435 );
and ( n54437 , n18144 , n6971 );
and ( n54438 , n19324 , n6504 );
xor ( n54439 , n54437 , n54438 );
and ( n54440 , n20233 , n6132 );
xor ( n54441 , n54439 , n54440 );
xor ( n54442 , n54436 , n54441 );
and ( n54443 , n15758 , n8243 );
and ( n54444 , n16637 , n7662 );
xor ( n54445 , n54443 , n54444 );
and ( n54446 , n17512 , n7310 );
xor ( n54447 , n54445 , n54446 );
xor ( n54448 , n54442 , n54447 );
xor ( n54449 , n54432 , n54448 );
and ( n54450 , n53262 , n53263 );
and ( n54451 , n53263 , n53265 );
and ( n54452 , n53262 , n53265 );
or ( n54453 , n54450 , n54451 , n54452 );
and ( n54454 , n11015 , n11718 );
and ( n54455 , n11769 , n10977 );
and ( n54456 , n54454 , n54455 );
and ( n54457 , n54455 , n53293 );
and ( n54458 , n54454 , n53293 );
or ( n54459 , n54456 , n54457 , n54458 );
xor ( n54460 , n54453 , n54459 );
and ( n54461 , n13322 , n10239 );
and ( n54462 , n14118 , n9348 );
xor ( n54463 , n54461 , n54462 );
and ( n54464 , n14938 , n8669 );
xor ( n54465 , n54463 , n54464 );
xor ( n54466 , n54460 , n54465 );
xor ( n54467 , n54449 , n54466 );
xor ( n54468 , n54428 , n54467 );
xor ( n54469 , n54398 , n54468 );
and ( n54470 , n53283 , n53287 );
and ( n54471 , n53287 , n53301 );
and ( n54472 , n53283 , n53301 );
or ( n54473 , n54470 , n54471 , n54472 );
and ( n54474 , n53320 , n53335 );
and ( n54475 , n53335 , n53352 );
and ( n54476 , n53320 , n53352 );
or ( n54477 , n54474 , n54475 , n54476 );
xor ( n54478 , n54473 , n54477 );
and ( n54479 , n53292 , n53294 );
and ( n54480 , n53294 , n53300 );
and ( n54481 , n53292 , n53300 );
or ( n54482 , n54479 , n54480 , n54481 );
and ( n54483 , n53324 , n53328 );
and ( n54484 , n53328 , n53334 );
and ( n54485 , n53324 , n53334 );
or ( n54486 , n54483 , n54484 , n54485 );
xor ( n54487 , n54482 , n54486 );
and ( n54488 , n53296 , n53297 );
and ( n54489 , n53297 , n53299 );
and ( n54490 , n53296 , n53299 );
or ( n54491 , n54488 , n54489 , n54490 );
and ( n54492 , n11015 , n12531 );
buf ( n54493 , n11769 );
xor ( n54494 , n54492 , n54493 );
and ( n54495 , n12320 , n10977 );
xor ( n54496 , n54494 , n54495 );
xor ( n54497 , n54491 , n54496 );
and ( n54498 , n8718 , n14838 );
and ( n54499 , n9400 , n14044 );
xor ( n54500 , n54498 , n54499 );
and ( n54501 , n10291 , n13256 );
xor ( n54502 , n54500 , n54501 );
xor ( n54503 , n54497 , n54502 );
xor ( n54504 , n54487 , n54503 );
xor ( n54505 , n54478 , n54504 );
xor ( n54506 , n54469 , n54505 );
xor ( n54507 , n54394 , n54506 );
xor ( n54508 , n54385 , n54507 );
and ( n54509 , n53316 , n53353 );
and ( n54510 , n53353 , n53379 );
and ( n54511 , n53316 , n53379 );
or ( n54512 , n54509 , n54510 , n54511 );
and ( n54513 , n53385 , n53414 );
xor ( n54514 , n54512 , n54513 );
and ( n54515 , n53358 , n53362 );
and ( n54516 , n53362 , n53378 );
and ( n54517 , n53358 , n53378 );
or ( n54518 , n54515 , n54516 , n54517 );
and ( n54519 , n53340 , n53345 );
and ( n54520 , n53345 , n53351 );
and ( n54521 , n53340 , n53351 );
or ( n54522 , n54519 , n54520 , n54521 );
and ( n54523 , n53330 , n53331 );
and ( n54524 , n53331 , n53333 );
and ( n54525 , n53330 , n53333 );
or ( n54526 , n54523 , n54524 , n54525 );
and ( n54527 , n53341 , n53342 );
and ( n54528 , n53342 , n53344 );
and ( n54529 , n53341 , n53344 );
or ( n54530 , n54527 , n54528 , n54529 );
xor ( n54531 , n54526 , n54530 );
and ( n54532 , n7385 , n17422 );
and ( n54533 , n7808 , n16550 );
xor ( n54534 , n54532 , n54533 );
and ( n54535 , n8079 , n15691 );
xor ( n54536 , n54534 , n54535 );
xor ( n54537 , n54531 , n54536 );
xor ( n54538 , n54522 , n54537 );
and ( n54539 , n53347 , n53348 );
and ( n54540 , n53348 , n53350 );
and ( n54541 , n53347 , n53350 );
or ( n54542 , n54539 , n54540 , n54541 );
and ( n54543 , n6187 , n20156 );
and ( n54544 , n6569 , n19222 );
xor ( n54545 , n54543 , n54544 );
and ( n54546 , n6816 , n18407 );
xor ( n54547 , n54545 , n54546 );
xor ( n54548 , n54542 , n54547 );
and ( n54549 , n4959 , n23075 );
and ( n54550 , n5459 , n22065 );
xor ( n54551 , n54549 , n54550 );
and ( n54552 , n5819 , n20976 );
xor ( n54553 , n54551 , n54552 );
xor ( n54554 , n54548 , n54553 );
xor ( n54555 , n54538 , n54554 );
xor ( n54556 , n54518 , n54555 );
and ( n54557 , n53367 , n53371 );
and ( n54558 , n53371 , n53377 );
and ( n54559 , n53367 , n53377 );
or ( n54560 , n54557 , n54558 , n54559 );
and ( n54561 , n53390 , n53395 );
and ( n54562 , n53395 , n53401 );
and ( n54563 , n53390 , n53401 );
or ( n54564 , n54561 , n54562 , n54563 );
xor ( n54565 , n54560 , n54564 );
and ( n54566 , n53397 , n53398 );
and ( n54567 , n53398 , n53400 );
and ( n54568 , n53397 , n53400 );
or ( n54569 , n54566 , n54567 , n54568 );
and ( n54570 , n53373 , n53374 );
and ( n54571 , n53374 , n53376 );
and ( n54572 , n53373 , n53376 );
or ( n54573 , n54570 , n54571 , n54572 );
xor ( n54574 , n54569 , n54573 );
and ( n54575 , n4132 , n26216 );
and ( n54576 , n4438 , n25163 );
xor ( n54577 , n54575 , n54576 );
and ( n54578 , n4766 , n24137 );
xor ( n54579 , n54577 , n54578 );
xor ( n54580 , n54574 , n54579 );
xor ( n54581 , n54565 , n54580 );
xor ( n54582 , n54556 , n54581 );
xor ( n54583 , n54514 , n54582 );
and ( n54584 , n53386 , n53402 );
and ( n54585 , n53402 , n53413 );
and ( n54586 , n53386 , n53413 );
or ( n54587 , n54584 , n54585 , n54586 );
and ( n54588 , n53407 , n53412 );
and ( n54589 , n53391 , n53392 );
and ( n54590 , n53392 , n53394 );
and ( n54591 , n53391 , n53394 );
or ( n54592 , n54589 , n54590 , n54591 );
and ( n54593 , n3182 , n29508 );
and ( n54594 , n3545 , n28406 );
xor ( n54595 , n54593 , n54594 );
and ( n54596 , n3801 , n27296 );
xor ( n54597 , n54595 , n54596 );
xor ( n54598 , n54592 , n54597 );
and ( n54599 , n2462 , n32999 );
and ( n54600 , n2779 , n31761 );
xor ( n54601 , n54599 , n54600 );
and ( n54602 , n3024 , n30629 );
xor ( n54603 , n54601 , n54602 );
xor ( n54604 , n54598 , n54603 );
xor ( n54605 , n54588 , n54604 );
and ( n54606 , n53410 , n53411 );
not ( n54607 , n2324 );
and ( n54608 , n34193 , n2324 );
nor ( n54609 , n54607 , n54608 );
xor ( n54610 , n54606 , n54609 );
xor ( n54611 , n54605 , n54610 );
xor ( n54612 , n54587 , n54611 );
xor ( n54613 , n54583 , n54612 );
xor ( n54614 , n54508 , n54613 );
xor ( n54615 , n54384 , n54614 );
xor ( n54616 , n54302 , n54615 );
xor ( n54617 , n54293 , n54616 );
and ( n54618 , n53089 , n53092 );
and ( n54619 , n53092 , n53419 );
and ( n54620 , n53089 , n53419 );
or ( n54621 , n54618 , n54619 , n54620 );
xor ( n54622 , n54617 , n54621 );
and ( n54623 , n53420 , n53424 );
and ( n54624 , n53425 , n53428 );
or ( n54625 , n54623 , n54624 );
xor ( n54626 , n54622 , n54625 );
buf ( n54627 , n54626 );
buf ( n54628 , n54627 );
not ( n54629 , n54628 );
nor ( n54630 , n54629 , n8739 );
xor ( n54631 , n54285 , n54630 );
and ( n54632 , n53085 , n53433 );
and ( n54633 , n53434 , n53437 );
or ( n54634 , n54632 , n54633 );
xor ( n54635 , n54631 , n54634 );
buf ( n54636 , n54635 );
buf ( n54637 , n54636 );
not ( n54638 , n54637 );
buf ( n54639 , n579 );
not ( n54640 , n54639 );
nor ( n54641 , n54638 , n54640 );
xor ( n54642 , n53911 , n54641 );
xor ( n54643 , n53449 , n53908 );
nor ( n54644 , n53441 , n54640 );
and ( n54645 , n54643 , n54644 );
xor ( n54646 , n54643 , n54644 );
xor ( n54647 , n53453 , n53906 );
nor ( n54648 , n52247 , n54640 );
and ( n54649 , n54647 , n54648 );
xor ( n54650 , n54647 , n54648 );
xor ( n54651 , n53457 , n53904 );
nor ( n54652 , n51049 , n54640 );
and ( n54653 , n54651 , n54652 );
xor ( n54654 , n54651 , n54652 );
xor ( n54655 , n53461 , n53902 );
nor ( n54656 , n49850 , n54640 );
and ( n54657 , n54655 , n54656 );
xor ( n54658 , n54655 , n54656 );
xor ( n54659 , n53465 , n53900 );
nor ( n54660 , n48650 , n54640 );
and ( n54661 , n54659 , n54660 );
xor ( n54662 , n54659 , n54660 );
xor ( n54663 , n53469 , n53898 );
nor ( n54664 , n47449 , n54640 );
and ( n54665 , n54663 , n54664 );
xor ( n54666 , n54663 , n54664 );
xor ( n54667 , n53473 , n53896 );
nor ( n54668 , n46248 , n54640 );
and ( n54669 , n54667 , n54668 );
xor ( n54670 , n54667 , n54668 );
xor ( n54671 , n53477 , n53894 );
nor ( n54672 , n45047 , n54640 );
and ( n54673 , n54671 , n54672 );
xor ( n54674 , n54671 , n54672 );
xor ( n54675 , n53481 , n53892 );
nor ( n54676 , n43843 , n54640 );
and ( n54677 , n54675 , n54676 );
xor ( n54678 , n54675 , n54676 );
xor ( n54679 , n53485 , n53890 );
nor ( n54680 , n42641 , n54640 );
and ( n54681 , n54679 , n54680 );
xor ( n54682 , n54679 , n54680 );
xor ( n54683 , n53489 , n53888 );
nor ( n54684 , n41437 , n54640 );
and ( n54685 , n54683 , n54684 );
xor ( n54686 , n54683 , n54684 );
xor ( n54687 , n53493 , n53886 );
nor ( n54688 , n40232 , n54640 );
and ( n54689 , n54687 , n54688 );
xor ( n54690 , n54687 , n54688 );
xor ( n54691 , n53497 , n53884 );
nor ( n54692 , n39027 , n54640 );
and ( n54693 , n54691 , n54692 );
xor ( n54694 , n54691 , n54692 );
xor ( n54695 , n53501 , n53882 );
nor ( n54696 , n37825 , n54640 );
and ( n54697 , n54695 , n54696 );
xor ( n54698 , n54695 , n54696 );
xor ( n54699 , n53505 , n53880 );
nor ( n54700 , n36620 , n54640 );
and ( n54701 , n54699 , n54700 );
xor ( n54702 , n54699 , n54700 );
xor ( n54703 , n53509 , n53878 );
nor ( n54704 , n35419 , n54640 );
and ( n54705 , n54703 , n54704 );
xor ( n54706 , n54703 , n54704 );
xor ( n54707 , n53513 , n53876 );
nor ( n54708 , n34224 , n54640 );
and ( n54709 , n54707 , n54708 );
xor ( n54710 , n54707 , n54708 );
xor ( n54711 , n53517 , n53874 );
nor ( n54712 , n33033 , n54640 );
and ( n54713 , n54711 , n54712 );
xor ( n54714 , n54711 , n54712 );
xor ( n54715 , n53521 , n53872 );
nor ( n54716 , n31867 , n54640 );
and ( n54717 , n54715 , n54716 );
xor ( n54718 , n54715 , n54716 );
xor ( n54719 , n53525 , n53870 );
nor ( n54720 , n30725 , n54640 );
and ( n54721 , n54719 , n54720 );
xor ( n54722 , n54719 , n54720 );
xor ( n54723 , n53529 , n53868 );
nor ( n54724 , n29596 , n54640 );
and ( n54725 , n54723 , n54724 );
xor ( n54726 , n54723 , n54724 );
xor ( n54727 , n53533 , n53866 );
nor ( n54728 , n28487 , n54640 );
and ( n54729 , n54727 , n54728 );
xor ( n54730 , n54727 , n54728 );
xor ( n54731 , n53537 , n53864 );
nor ( n54732 , n27397 , n54640 );
and ( n54733 , n54731 , n54732 );
xor ( n54734 , n54731 , n54732 );
xor ( n54735 , n53541 , n53862 );
nor ( n54736 , n26326 , n54640 );
and ( n54737 , n54735 , n54736 );
xor ( n54738 , n54735 , n54736 );
xor ( n54739 , n53545 , n53860 );
nor ( n54740 , n25272 , n54640 );
and ( n54741 , n54739 , n54740 );
xor ( n54742 , n54739 , n54740 );
xor ( n54743 , n53549 , n53858 );
nor ( n54744 , n24242 , n54640 );
and ( n54745 , n54743 , n54744 );
xor ( n54746 , n54743 , n54744 );
xor ( n54747 , n53553 , n53856 );
nor ( n54748 , n23225 , n54640 );
and ( n54749 , n54747 , n54748 );
xor ( n54750 , n54747 , n54748 );
xor ( n54751 , n53557 , n53854 );
nor ( n54752 , n22231 , n54640 );
and ( n54753 , n54751 , n54752 );
xor ( n54754 , n54751 , n54752 );
xor ( n54755 , n53561 , n53852 );
nor ( n54756 , n21258 , n54640 );
and ( n54757 , n54755 , n54756 );
xor ( n54758 , n54755 , n54756 );
xor ( n54759 , n53565 , n53850 );
nor ( n54760 , n20303 , n54640 );
and ( n54761 , n54759 , n54760 );
xor ( n54762 , n54759 , n54760 );
xor ( n54763 , n53569 , n53848 );
nor ( n54764 , n19365 , n54640 );
and ( n54765 , n54763 , n54764 );
xor ( n54766 , n54763 , n54764 );
xor ( n54767 , n53573 , n53846 );
nor ( n54768 , n18448 , n54640 );
and ( n54769 , n54767 , n54768 );
xor ( n54770 , n54767 , n54768 );
xor ( n54771 , n53577 , n53844 );
nor ( n54772 , n17548 , n54640 );
and ( n54773 , n54771 , n54772 );
xor ( n54774 , n54771 , n54772 );
xor ( n54775 , n53581 , n53842 );
nor ( n54776 , n16669 , n54640 );
and ( n54777 , n54775 , n54776 );
xor ( n54778 , n54775 , n54776 );
xor ( n54779 , n53585 , n53840 );
nor ( n54780 , n15809 , n54640 );
and ( n54781 , n54779 , n54780 );
xor ( n54782 , n54779 , n54780 );
xor ( n54783 , n53589 , n53838 );
nor ( n54784 , n14968 , n54640 );
and ( n54785 , n54783 , n54784 );
xor ( n54786 , n54783 , n54784 );
xor ( n54787 , n53593 , n53836 );
nor ( n54788 , n14147 , n54640 );
and ( n54789 , n54787 , n54788 );
xor ( n54790 , n54787 , n54788 );
xor ( n54791 , n53597 , n53834 );
nor ( n54792 , n13349 , n54640 );
and ( n54793 , n54791 , n54792 );
xor ( n54794 , n54791 , n54792 );
xor ( n54795 , n53601 , n53832 );
nor ( n54796 , n12564 , n54640 );
and ( n54797 , n54795 , n54796 );
xor ( n54798 , n54795 , n54796 );
xor ( n54799 , n53605 , n53830 );
nor ( n54800 , n11799 , n54640 );
and ( n54801 , n54799 , n54800 );
xor ( n54802 , n54799 , n54800 );
xor ( n54803 , n53609 , n53828 );
nor ( n54804 , n11050 , n54640 );
and ( n54805 , n54803 , n54804 );
xor ( n54806 , n54803 , n54804 );
xor ( n54807 , n53613 , n53826 );
nor ( n54808 , n10321 , n54640 );
and ( n54809 , n54807 , n54808 );
xor ( n54810 , n54807 , n54808 );
xor ( n54811 , n53617 , n53824 );
nor ( n54812 , n9429 , n54640 );
and ( n54813 , n54811 , n54812 );
xor ( n54814 , n54811 , n54812 );
xor ( n54815 , n53621 , n53822 );
nor ( n54816 , n8949 , n54640 );
and ( n54817 , n54815 , n54816 );
xor ( n54818 , n54815 , n54816 );
xor ( n54819 , n53625 , n53820 );
nor ( n54820 , n9437 , n54640 );
and ( n54821 , n54819 , n54820 );
xor ( n54822 , n54819 , n54820 );
xor ( n54823 , n53629 , n53818 );
nor ( n54824 , n9446 , n54640 );
and ( n54825 , n54823 , n54824 );
xor ( n54826 , n54823 , n54824 );
xor ( n54827 , n53633 , n53816 );
nor ( n54828 , n9455 , n54640 );
and ( n54829 , n54827 , n54828 );
xor ( n54830 , n54827 , n54828 );
xor ( n54831 , n53637 , n53814 );
nor ( n54832 , n9464 , n54640 );
and ( n54833 , n54831 , n54832 );
xor ( n54834 , n54831 , n54832 );
xor ( n54835 , n53641 , n53812 );
nor ( n54836 , n9473 , n54640 );
and ( n54837 , n54835 , n54836 );
xor ( n54838 , n54835 , n54836 );
xor ( n54839 , n53645 , n53810 );
nor ( n54840 , n9482 , n54640 );
and ( n54841 , n54839 , n54840 );
xor ( n54842 , n54839 , n54840 );
xor ( n54843 , n53649 , n53808 );
nor ( n54844 , n9491 , n54640 );
and ( n54845 , n54843 , n54844 );
xor ( n54846 , n54843 , n54844 );
xor ( n54847 , n53653 , n53806 );
nor ( n54848 , n9500 , n54640 );
and ( n54849 , n54847 , n54848 );
xor ( n54850 , n54847 , n54848 );
xor ( n54851 , n53657 , n53804 );
nor ( n54852 , n9509 , n54640 );
and ( n54853 , n54851 , n54852 );
xor ( n54854 , n54851 , n54852 );
xor ( n54855 , n53661 , n53802 );
nor ( n54856 , n9518 , n54640 );
and ( n54857 , n54855 , n54856 );
xor ( n54858 , n54855 , n54856 );
xor ( n54859 , n53665 , n53800 );
nor ( n54860 , n9527 , n54640 );
and ( n54861 , n54859 , n54860 );
xor ( n54862 , n54859 , n54860 );
xor ( n54863 , n53669 , n53798 );
nor ( n54864 , n9536 , n54640 );
and ( n54865 , n54863 , n54864 );
xor ( n54866 , n54863 , n54864 );
xor ( n54867 , n53673 , n53796 );
nor ( n54868 , n9545 , n54640 );
and ( n54869 , n54867 , n54868 );
xor ( n54870 , n54867 , n54868 );
xor ( n54871 , n53677 , n53794 );
nor ( n54872 , n9554 , n54640 );
and ( n54873 , n54871 , n54872 );
xor ( n54874 , n54871 , n54872 );
xor ( n54875 , n53681 , n53792 );
nor ( n54876 , n9563 , n54640 );
and ( n54877 , n54875 , n54876 );
xor ( n54878 , n54875 , n54876 );
xor ( n54879 , n53685 , n53790 );
nor ( n54880 , n9572 , n54640 );
and ( n54881 , n54879 , n54880 );
xor ( n54882 , n54879 , n54880 );
xor ( n54883 , n53689 , n53788 );
nor ( n54884 , n9581 , n54640 );
and ( n54885 , n54883 , n54884 );
xor ( n54886 , n54883 , n54884 );
xor ( n54887 , n53693 , n53786 );
nor ( n54888 , n9590 , n54640 );
and ( n54889 , n54887 , n54888 );
xor ( n54890 , n54887 , n54888 );
xor ( n54891 , n53697 , n53784 );
nor ( n54892 , n9599 , n54640 );
and ( n54893 , n54891 , n54892 );
xor ( n54894 , n54891 , n54892 );
xor ( n54895 , n53701 , n53782 );
nor ( n54896 , n9608 , n54640 );
and ( n54897 , n54895 , n54896 );
xor ( n54898 , n54895 , n54896 );
xor ( n54899 , n53705 , n53780 );
nor ( n54900 , n9617 , n54640 );
and ( n54901 , n54899 , n54900 );
xor ( n54902 , n54899 , n54900 );
xor ( n54903 , n53709 , n53778 );
nor ( n54904 , n9626 , n54640 );
and ( n54905 , n54903 , n54904 );
xor ( n54906 , n54903 , n54904 );
xor ( n54907 , n53713 , n53776 );
nor ( n54908 , n9635 , n54640 );
and ( n54909 , n54907 , n54908 );
xor ( n54910 , n54907 , n54908 );
xor ( n54911 , n53717 , n53774 );
nor ( n54912 , n9644 , n54640 );
and ( n54913 , n54911 , n54912 );
xor ( n54914 , n54911 , n54912 );
xor ( n54915 , n53721 , n53772 );
nor ( n54916 , n9653 , n54640 );
and ( n54917 , n54915 , n54916 );
xor ( n54918 , n54915 , n54916 );
xor ( n54919 , n53725 , n53770 );
nor ( n54920 , n9662 , n54640 );
and ( n54921 , n54919 , n54920 );
xor ( n54922 , n54919 , n54920 );
xor ( n54923 , n53729 , n53768 );
nor ( n54924 , n9671 , n54640 );
and ( n54925 , n54923 , n54924 );
xor ( n54926 , n54923 , n54924 );
xor ( n54927 , n53733 , n53766 );
nor ( n54928 , n9680 , n54640 );
and ( n54929 , n54927 , n54928 );
xor ( n54930 , n54927 , n54928 );
xor ( n54931 , n53737 , n53764 );
nor ( n54932 , n9689 , n54640 );
and ( n54933 , n54931 , n54932 );
xor ( n54934 , n54931 , n54932 );
xor ( n54935 , n53741 , n53762 );
nor ( n54936 , n9698 , n54640 );
and ( n54937 , n54935 , n54936 );
xor ( n54938 , n54935 , n54936 );
xor ( n54939 , n53745 , n53760 );
nor ( n54940 , n9707 , n54640 );
and ( n54941 , n54939 , n54940 );
xor ( n54942 , n54939 , n54940 );
xor ( n54943 , n53749 , n53758 );
nor ( n54944 , n9716 , n54640 );
and ( n54945 , n54943 , n54944 );
xor ( n54946 , n54943 , n54944 );
xor ( n54947 , n53753 , n53756 );
nor ( n54948 , n9725 , n54640 );
and ( n54949 , n54947 , n54948 );
xor ( n54950 , n54947 , n54948 );
xor ( n54951 , n53754 , n53755 );
nor ( n54952 , n9734 , n54640 );
and ( n54953 , n54951 , n54952 );
xor ( n54954 , n54951 , n54952 );
nor ( n54955 , n9752 , n53443 );
nor ( n54956 , n9743 , n54640 );
and ( n54957 , n54955 , n54956 );
and ( n54958 , n54954 , n54957 );
or ( n54959 , n54953 , n54958 );
and ( n54960 , n54950 , n54959 );
or ( n54961 , n54949 , n54960 );
and ( n54962 , n54946 , n54961 );
or ( n54963 , n54945 , n54962 );
and ( n54964 , n54942 , n54963 );
or ( n54965 , n54941 , n54964 );
and ( n54966 , n54938 , n54965 );
or ( n54967 , n54937 , n54966 );
and ( n54968 , n54934 , n54967 );
or ( n54969 , n54933 , n54968 );
and ( n54970 , n54930 , n54969 );
or ( n54971 , n54929 , n54970 );
and ( n54972 , n54926 , n54971 );
or ( n54973 , n54925 , n54972 );
and ( n54974 , n54922 , n54973 );
or ( n54975 , n54921 , n54974 );
and ( n54976 , n54918 , n54975 );
or ( n54977 , n54917 , n54976 );
and ( n54978 , n54914 , n54977 );
or ( n54979 , n54913 , n54978 );
and ( n54980 , n54910 , n54979 );
or ( n54981 , n54909 , n54980 );
and ( n54982 , n54906 , n54981 );
or ( n54983 , n54905 , n54982 );
and ( n54984 , n54902 , n54983 );
or ( n54985 , n54901 , n54984 );
and ( n54986 , n54898 , n54985 );
or ( n54987 , n54897 , n54986 );
and ( n54988 , n54894 , n54987 );
or ( n54989 , n54893 , n54988 );
and ( n54990 , n54890 , n54989 );
or ( n54991 , n54889 , n54990 );
and ( n54992 , n54886 , n54991 );
or ( n54993 , n54885 , n54992 );
and ( n54994 , n54882 , n54993 );
or ( n54995 , n54881 , n54994 );
and ( n54996 , n54878 , n54995 );
or ( n54997 , n54877 , n54996 );
and ( n54998 , n54874 , n54997 );
or ( n54999 , n54873 , n54998 );
and ( n55000 , n54870 , n54999 );
or ( n55001 , n54869 , n55000 );
and ( n55002 , n54866 , n55001 );
or ( n55003 , n54865 , n55002 );
and ( n55004 , n54862 , n55003 );
or ( n55005 , n54861 , n55004 );
and ( n55006 , n54858 , n55005 );
or ( n55007 , n54857 , n55006 );
and ( n55008 , n54854 , n55007 );
or ( n55009 , n54853 , n55008 );
and ( n55010 , n54850 , n55009 );
or ( n55011 , n54849 , n55010 );
and ( n55012 , n54846 , n55011 );
or ( n55013 , n54845 , n55012 );
and ( n55014 , n54842 , n55013 );
or ( n55015 , n54841 , n55014 );
and ( n55016 , n54838 , n55015 );
or ( n55017 , n54837 , n55016 );
and ( n55018 , n54834 , n55017 );
or ( n55019 , n54833 , n55018 );
and ( n55020 , n54830 , n55019 );
or ( n55021 , n54829 , n55020 );
and ( n55022 , n54826 , n55021 );
or ( n55023 , n54825 , n55022 );
and ( n55024 , n54822 , n55023 );
or ( n55025 , n54821 , n55024 );
and ( n55026 , n54818 , n55025 );
or ( n55027 , n54817 , n55026 );
and ( n55028 , n54814 , n55027 );
or ( n55029 , n54813 , n55028 );
and ( n55030 , n54810 , n55029 );
or ( n55031 , n54809 , n55030 );
and ( n55032 , n54806 , n55031 );
or ( n55033 , n54805 , n55032 );
and ( n55034 , n54802 , n55033 );
or ( n55035 , n54801 , n55034 );
and ( n55036 , n54798 , n55035 );
or ( n55037 , n54797 , n55036 );
and ( n55038 , n54794 , n55037 );
or ( n55039 , n54793 , n55038 );
and ( n55040 , n54790 , n55039 );
or ( n55041 , n54789 , n55040 );
and ( n55042 , n54786 , n55041 );
or ( n55043 , n54785 , n55042 );
and ( n55044 , n54782 , n55043 );
or ( n55045 , n54781 , n55044 );
and ( n55046 , n54778 , n55045 );
or ( n55047 , n54777 , n55046 );
and ( n55048 , n54774 , n55047 );
or ( n55049 , n54773 , n55048 );
and ( n55050 , n54770 , n55049 );
or ( n55051 , n54769 , n55050 );
and ( n55052 , n54766 , n55051 );
or ( n55053 , n54765 , n55052 );
and ( n55054 , n54762 , n55053 );
or ( n55055 , n54761 , n55054 );
and ( n55056 , n54758 , n55055 );
or ( n55057 , n54757 , n55056 );
and ( n55058 , n54754 , n55057 );
or ( n55059 , n54753 , n55058 );
and ( n55060 , n54750 , n55059 );
or ( n55061 , n54749 , n55060 );
and ( n55062 , n54746 , n55061 );
or ( n55063 , n54745 , n55062 );
and ( n55064 , n54742 , n55063 );
or ( n55065 , n54741 , n55064 );
and ( n55066 , n54738 , n55065 );
or ( n55067 , n54737 , n55066 );
and ( n55068 , n54734 , n55067 );
or ( n55069 , n54733 , n55068 );
and ( n55070 , n54730 , n55069 );
or ( n55071 , n54729 , n55070 );
and ( n55072 , n54726 , n55071 );
or ( n55073 , n54725 , n55072 );
and ( n55074 , n54722 , n55073 );
or ( n55075 , n54721 , n55074 );
and ( n55076 , n54718 , n55075 );
or ( n55077 , n54717 , n55076 );
and ( n55078 , n54714 , n55077 );
or ( n55079 , n54713 , n55078 );
and ( n55080 , n54710 , n55079 );
or ( n55081 , n54709 , n55080 );
and ( n55082 , n54706 , n55081 );
or ( n55083 , n54705 , n55082 );
and ( n55084 , n54702 , n55083 );
or ( n55085 , n54701 , n55084 );
and ( n55086 , n54698 , n55085 );
or ( n55087 , n54697 , n55086 );
and ( n55088 , n54694 , n55087 );
or ( n55089 , n54693 , n55088 );
and ( n55090 , n54690 , n55089 );
or ( n55091 , n54689 , n55090 );
and ( n55092 , n54686 , n55091 );
or ( n55093 , n54685 , n55092 );
and ( n55094 , n54682 , n55093 );
or ( n55095 , n54681 , n55094 );
and ( n55096 , n54678 , n55095 );
or ( n55097 , n54677 , n55096 );
and ( n55098 , n54674 , n55097 );
or ( n55099 , n54673 , n55098 );
and ( n55100 , n54670 , n55099 );
or ( n55101 , n54669 , n55100 );
and ( n55102 , n54666 , n55101 );
or ( n55103 , n54665 , n55102 );
and ( n55104 , n54662 , n55103 );
or ( n55105 , n54661 , n55104 );
and ( n55106 , n54658 , n55105 );
or ( n55107 , n54657 , n55106 );
and ( n55108 , n54654 , n55107 );
or ( n55109 , n54653 , n55108 );
and ( n55110 , n54650 , n55109 );
or ( n55111 , n54649 , n55110 );
and ( n55112 , n54646 , n55111 );
or ( n55113 , n54645 , n55112 );
xor ( n55114 , n54642 , n55113 );
and ( n55115 , n33403 , n2565 );
nor ( n55116 , n2566 , n55115 );
nor ( n55117 , n2797 , n32231 );
xor ( n55118 , n55116 , n55117 );
and ( n55119 , n53913 , n53914 );
and ( n55120 , n53915 , n53918 );
or ( n55121 , n55119 , n55120 );
xor ( n55122 , n55118 , n55121 );
nor ( n55123 , n3043 , n31083 );
xor ( n55124 , n55122 , n55123 );
and ( n55125 , n53919 , n53920 );
and ( n55126 , n53921 , n53924 );
or ( n55127 , n55125 , n55126 );
xor ( n55128 , n55124 , n55127 );
nor ( n55129 , n3300 , n29948 );
xor ( n55130 , n55128 , n55129 );
and ( n55131 , n53925 , n53926 );
and ( n55132 , n53927 , n53930 );
or ( n55133 , n55131 , n55132 );
xor ( n55134 , n55130 , n55133 );
nor ( n55135 , n3570 , n28833 );
xor ( n55136 , n55134 , n55135 );
and ( n55137 , n53931 , n53932 );
and ( n55138 , n53933 , n53936 );
or ( n55139 , n55137 , n55138 );
xor ( n55140 , n55136 , n55139 );
nor ( n55141 , n3853 , n27737 );
xor ( n55142 , n55140 , n55141 );
and ( n55143 , n53937 , n53938 );
and ( n55144 , n53939 , n53942 );
or ( n55145 , n55143 , n55144 );
xor ( n55146 , n55142 , n55145 );
nor ( n55147 , n4151 , n26660 );
xor ( n55148 , n55146 , n55147 );
and ( n55149 , n53943 , n53944 );
and ( n55150 , n53945 , n53948 );
or ( n55151 , n55149 , n55150 );
xor ( n55152 , n55148 , n55151 );
nor ( n55153 , n4458 , n25600 );
xor ( n55154 , n55152 , n55153 );
and ( n55155 , n53949 , n53950 );
and ( n55156 , n53951 , n53954 );
or ( n55157 , n55155 , n55156 );
xor ( n55158 , n55154 , n55157 );
nor ( n55159 , n4786 , n24564 );
xor ( n55160 , n55158 , n55159 );
and ( n55161 , n53955 , n53956 );
and ( n55162 , n53957 , n53960 );
or ( n55163 , n55161 , n55162 );
xor ( n55164 , n55160 , n55163 );
nor ( n55165 , n5126 , n23541 );
xor ( n55166 , n55164 , n55165 );
and ( n55167 , n53961 , n53962 );
and ( n55168 , n53963 , n53966 );
or ( n55169 , n55167 , n55168 );
xor ( n55170 , n55166 , n55169 );
nor ( n55171 , n5477 , n22541 );
xor ( n55172 , n55170 , n55171 );
and ( n55173 , n53967 , n53968 );
and ( n55174 , n53969 , n53972 );
or ( n55175 , n55173 , n55174 );
xor ( n55176 , n55172 , n55175 );
nor ( n55177 , n5838 , n21562 );
xor ( n55178 , n55176 , n55177 );
and ( n55179 , n53973 , n53974 );
and ( n55180 , n53975 , n53978 );
or ( n55181 , n55179 , n55180 );
xor ( n55182 , n55178 , n55181 );
nor ( n55183 , n6212 , n20601 );
xor ( n55184 , n55182 , n55183 );
and ( n55185 , n53979 , n53980 );
and ( n55186 , n53981 , n53984 );
or ( n55187 , n55185 , n55186 );
xor ( n55188 , n55184 , n55187 );
nor ( n55189 , n6596 , n19657 );
xor ( n55190 , n55188 , n55189 );
and ( n55191 , n53985 , n53986 );
and ( n55192 , n53987 , n53990 );
or ( n55193 , n55191 , n55192 );
xor ( n55194 , n55190 , n55193 );
nor ( n55195 , n6997 , n18734 );
xor ( n55196 , n55194 , n55195 );
and ( n55197 , n53991 , n53992 );
and ( n55198 , n53993 , n53996 );
or ( n55199 , n55197 , n55198 );
xor ( n55200 , n55196 , n55199 );
nor ( n55201 , n7413 , n17828 );
xor ( n55202 , n55200 , n55201 );
and ( n55203 , n53997 , n53998 );
and ( n55204 , n53999 , n54002 );
or ( n55205 , n55203 , n55204 );
xor ( n55206 , n55202 , n55205 );
nor ( n55207 , n7841 , n16943 );
xor ( n55208 , n55206 , n55207 );
and ( n55209 , n54003 , n54004 );
and ( n55210 , n54005 , n54008 );
or ( n55211 , n55209 , n55210 );
xor ( n55212 , n55208 , n55211 );
nor ( n55213 , n8281 , n16077 );
xor ( n55214 , n55212 , n55213 );
and ( n55215 , n54009 , n54010 );
and ( n55216 , n54011 , n54014 );
or ( n55217 , n55215 , n55216 );
xor ( n55218 , n55214 , n55217 );
nor ( n55219 , n8737 , n15230 );
xor ( n55220 , n55218 , n55219 );
and ( n55221 , n54015 , n54016 );
and ( n55222 , n54017 , n54020 );
or ( n55223 , n55221 , n55222 );
xor ( n55224 , n55220 , n55223 );
nor ( n55225 , n9420 , n14403 );
xor ( n55226 , n55224 , n55225 );
and ( n55227 , n54021 , n54022 );
and ( n55228 , n54023 , n54026 );
or ( n55229 , n55227 , n55228 );
xor ( n55230 , n55226 , n55229 );
nor ( n55231 , n10312 , n13599 );
xor ( n55232 , n55230 , n55231 );
and ( n55233 , n54027 , n54028 );
and ( n55234 , n54029 , n54032 );
or ( n55235 , n55233 , n55234 );
xor ( n55236 , n55232 , n55235 );
nor ( n55237 , n11041 , n12808 );
xor ( n55238 , n55236 , n55237 );
and ( n55239 , n54033 , n54034 );
and ( n55240 , n54035 , n54038 );
or ( n55241 , n55239 , n55240 );
xor ( n55242 , n55238 , n55241 );
nor ( n55243 , n11790 , n12037 );
xor ( n55244 , n55242 , n55243 );
and ( n55245 , n54039 , n54040 );
and ( n55246 , n54041 , n54044 );
or ( n55247 , n55245 , n55246 );
xor ( n55248 , n55244 , n55247 );
nor ( n55249 , n12555 , n11282 );
xor ( n55250 , n55248 , n55249 );
and ( n55251 , n54045 , n54046 );
and ( n55252 , n54047 , n54050 );
or ( n55253 , n55251 , n55252 );
xor ( n55254 , n55250 , n55253 );
nor ( n55255 , n13340 , n10547 );
xor ( n55256 , n55254 , n55255 );
and ( n55257 , n54051 , n54052 );
and ( n55258 , n54053 , n54056 );
or ( n55259 , n55257 , n55258 );
xor ( n55260 , n55256 , n55259 );
nor ( n55261 , n14138 , n9829 );
xor ( n55262 , n55260 , n55261 );
and ( n55263 , n54057 , n54058 );
and ( n55264 , n54059 , n54062 );
or ( n55265 , n55263 , n55264 );
xor ( n55266 , n55262 , n55265 );
nor ( n55267 , n14959 , n8955 );
xor ( n55268 , n55266 , n55267 );
and ( n55269 , n54063 , n54064 );
and ( n55270 , n54065 , n54068 );
or ( n55271 , n55269 , n55270 );
xor ( n55272 , n55268 , n55271 );
nor ( n55273 , n15800 , n603 );
xor ( n55274 , n55272 , n55273 );
and ( n55275 , n54069 , n54070 );
and ( n55276 , n54071 , n54074 );
or ( n55277 , n55275 , n55276 );
xor ( n55278 , n55274 , n55277 );
nor ( n55279 , n16660 , n652 );
xor ( n55280 , n55278 , n55279 );
and ( n55281 , n54075 , n54076 );
and ( n55282 , n54077 , n54080 );
or ( n55283 , n55281 , n55282 );
xor ( n55284 , n55280 , n55283 );
nor ( n55285 , n17539 , n624 );
xor ( n55286 , n55284 , n55285 );
and ( n55287 , n54081 , n54082 );
and ( n55288 , n54083 , n54086 );
or ( n55289 , n55287 , n55288 );
xor ( n55290 , n55286 , n55289 );
nor ( n55291 , n18439 , n648 );
xor ( n55292 , n55290 , n55291 );
and ( n55293 , n54087 , n54088 );
and ( n55294 , n54089 , n54092 );
or ( n55295 , n55293 , n55294 );
xor ( n55296 , n55292 , n55295 );
nor ( n55297 , n19356 , n686 );
xor ( n55298 , n55296 , n55297 );
and ( n55299 , n54093 , n54094 );
and ( n55300 , n54095 , n54098 );
or ( n55301 , n55299 , n55300 );
xor ( n55302 , n55298 , n55301 );
nor ( n55303 , n20294 , n735 );
xor ( n55304 , n55302 , n55303 );
and ( n55305 , n54099 , n54100 );
and ( n55306 , n54101 , n54104 );
or ( n55307 , n55305 , n55306 );
xor ( n55308 , n55304 , n55307 );
nor ( n55309 , n21249 , n798 );
xor ( n55310 , n55308 , n55309 );
and ( n55311 , n54105 , n54106 );
and ( n55312 , n54107 , n54110 );
or ( n55313 , n55311 , n55312 );
xor ( n55314 , n55310 , n55313 );
nor ( n55315 , n22222 , n870 );
xor ( n55316 , n55314 , n55315 );
and ( n55317 , n54111 , n54112 );
and ( n55318 , n54113 , n54116 );
or ( n55319 , n55317 , n55318 );
xor ( n55320 , n55316 , n55319 );
nor ( n55321 , n23216 , n960 );
xor ( n55322 , n55320 , n55321 );
and ( n55323 , n54117 , n54118 );
and ( n55324 , n54119 , n54122 );
or ( n55325 , n55323 , n55324 );
xor ( n55326 , n55322 , n55325 );
nor ( n55327 , n24233 , n1064 );
xor ( n55328 , n55326 , n55327 );
and ( n55329 , n54123 , n54124 );
and ( n55330 , n54125 , n54128 );
or ( n55331 , n55329 , n55330 );
xor ( n55332 , n55328 , n55331 );
nor ( n55333 , n25263 , n1178 );
xor ( n55334 , n55332 , n55333 );
and ( n55335 , n54129 , n54130 );
and ( n55336 , n54131 , n54134 );
or ( n55337 , n55335 , n55336 );
xor ( n55338 , n55334 , n55337 );
nor ( n55339 , n26317 , n1305 );
xor ( n55340 , n55338 , n55339 );
and ( n55341 , n54135 , n54136 );
and ( n55342 , n54137 , n54140 );
or ( n55343 , n55341 , n55342 );
xor ( n55344 , n55340 , n55343 );
nor ( n55345 , n27388 , n1447 );
xor ( n55346 , n55344 , n55345 );
and ( n55347 , n54141 , n54142 );
and ( n55348 , n54143 , n54146 );
or ( n55349 , n55347 , n55348 );
xor ( n55350 , n55346 , n55349 );
nor ( n55351 , n28478 , n1600 );
xor ( n55352 , n55350 , n55351 );
and ( n55353 , n54147 , n54148 );
and ( n55354 , n54149 , n54152 );
or ( n55355 , n55353 , n55354 );
xor ( n55356 , n55352 , n55355 );
nor ( n55357 , n29587 , n1768 );
xor ( n55358 , n55356 , n55357 );
and ( n55359 , n54153 , n54154 );
and ( n55360 , n54155 , n54158 );
or ( n55361 , n55359 , n55360 );
xor ( n55362 , n55358 , n55361 );
nor ( n55363 , n30716 , n1947 );
xor ( n55364 , n55362 , n55363 );
and ( n55365 , n54159 , n54160 );
and ( n55366 , n54161 , n54164 );
or ( n55367 , n55365 , n55366 );
xor ( n55368 , n55364 , n55367 );
nor ( n55369 , n31858 , n2139 );
xor ( n55370 , n55368 , n55369 );
and ( n55371 , n54165 , n54166 );
and ( n55372 , n54167 , n54170 );
or ( n55373 , n55371 , n55372 );
xor ( n55374 , n55370 , n55373 );
nor ( n55375 , n33024 , n2345 );
xor ( n55376 , n55374 , n55375 );
and ( n55377 , n54171 , n54172 );
and ( n55378 , n54173 , n54176 );
or ( n55379 , n55377 , n55378 );
xor ( n55380 , n55376 , n55379 );
nor ( n55381 , n34215 , n2568 );
xor ( n55382 , n55380 , n55381 );
and ( n55383 , n54177 , n54178 );
and ( n55384 , n54179 , n54182 );
or ( n55385 , n55383 , n55384 );
xor ( n55386 , n55382 , n55385 );
nor ( n55387 , n35410 , n2799 );
xor ( n55388 , n55386 , n55387 );
and ( n55389 , n54183 , n54184 );
and ( n55390 , n54185 , n54188 );
or ( n55391 , n55389 , n55390 );
xor ( n55392 , n55388 , n55391 );
nor ( n55393 , n36611 , n3045 );
xor ( n55394 , n55392 , n55393 );
and ( n55395 , n54189 , n54190 );
and ( n55396 , n54191 , n54194 );
or ( n55397 , n55395 , n55396 );
xor ( n55398 , n55394 , n55397 );
nor ( n55399 , n37816 , n3302 );
xor ( n55400 , n55398 , n55399 );
and ( n55401 , n54195 , n54196 );
and ( n55402 , n54197 , n54200 );
or ( n55403 , n55401 , n55402 );
xor ( n55404 , n55400 , n55403 );
nor ( n55405 , n39018 , n3572 );
xor ( n55406 , n55404 , n55405 );
and ( n55407 , n54201 , n54202 );
and ( n55408 , n54203 , n54206 );
or ( n55409 , n55407 , n55408 );
xor ( n55410 , n55406 , n55409 );
nor ( n55411 , n40223 , n3855 );
xor ( n55412 , n55410 , n55411 );
and ( n55413 , n54207 , n54208 );
and ( n55414 , n54209 , n54212 );
or ( n55415 , n55413 , n55414 );
xor ( n55416 , n55412 , n55415 );
nor ( n55417 , n41428 , n4153 );
xor ( n55418 , n55416 , n55417 );
and ( n55419 , n54213 , n54214 );
and ( n55420 , n54215 , n54218 );
or ( n55421 , n55419 , n55420 );
xor ( n55422 , n55418 , n55421 );
nor ( n55423 , n42632 , n4460 );
xor ( n55424 , n55422 , n55423 );
and ( n55425 , n54219 , n54220 );
and ( n55426 , n54221 , n54224 );
or ( n55427 , n55425 , n55426 );
xor ( n55428 , n55424 , n55427 );
nor ( n55429 , n43834 , n4788 );
xor ( n55430 , n55428 , n55429 );
and ( n55431 , n54225 , n54226 );
and ( n55432 , n54227 , n54230 );
or ( n55433 , n55431 , n55432 );
xor ( n55434 , n55430 , n55433 );
nor ( n55435 , n45038 , n5128 );
xor ( n55436 , n55434 , n55435 );
and ( n55437 , n54231 , n54232 );
and ( n55438 , n54233 , n54236 );
or ( n55439 , n55437 , n55438 );
xor ( n55440 , n55436 , n55439 );
nor ( n55441 , n46239 , n5479 );
xor ( n55442 , n55440 , n55441 );
and ( n55443 , n54237 , n54238 );
and ( n55444 , n54239 , n54242 );
or ( n55445 , n55443 , n55444 );
xor ( n55446 , n55442 , n55445 );
nor ( n55447 , n47440 , n5840 );
xor ( n55448 , n55446 , n55447 );
and ( n55449 , n54243 , n54244 );
and ( n55450 , n54245 , n54248 );
or ( n55451 , n55449 , n55450 );
xor ( n55452 , n55448 , n55451 );
nor ( n55453 , n48641 , n6214 );
xor ( n55454 , n55452 , n55453 );
and ( n55455 , n54249 , n54250 );
and ( n55456 , n54251 , n54254 );
or ( n55457 , n55455 , n55456 );
xor ( n55458 , n55454 , n55457 );
nor ( n55459 , n49841 , n6598 );
xor ( n55460 , n55458 , n55459 );
and ( n55461 , n54255 , n54256 );
and ( n55462 , n54257 , n54260 );
or ( n55463 , n55461 , n55462 );
xor ( n55464 , n55460 , n55463 );
nor ( n55465 , n51040 , n6999 );
xor ( n55466 , n55464 , n55465 );
and ( n55467 , n54261 , n54262 );
and ( n55468 , n54263 , n54266 );
or ( n55469 , n55467 , n55468 );
xor ( n55470 , n55466 , n55469 );
nor ( n55471 , n52238 , n7415 );
xor ( n55472 , n55470 , n55471 );
and ( n55473 , n54267 , n54268 );
and ( n55474 , n54269 , n54272 );
or ( n55475 , n55473 , n55474 );
xor ( n55476 , n55472 , n55475 );
nor ( n55477 , n53432 , n7843 );
xor ( n55478 , n55476 , n55477 );
and ( n55479 , n54273 , n54274 );
and ( n55480 , n54275 , n54278 );
or ( n55481 , n55479 , n55480 );
xor ( n55482 , n55478 , n55481 );
nor ( n55483 , n54629 , n8283 );
xor ( n55484 , n55482 , n55483 );
and ( n55485 , n54279 , n54280 );
and ( n55486 , n54281 , n54284 );
or ( n55487 , n55485 , n55486 );
xor ( n55488 , n55484 , n55487 );
and ( n55489 , n54297 , n54301 );
and ( n55490 , n54301 , n54615 );
and ( n55491 , n54297 , n54615 );
or ( n55492 , n55489 , n55490 , n55491 );
and ( n55493 , n33774 , n2544 );
not ( n55494 , n2544 );
nor ( n55495 , n55493 , n55494 );
xor ( n55496 , n55492 , n55495 );
and ( n55497 , n54310 , n54314 );
and ( n55498 , n54314 , n54382 );
and ( n55499 , n54310 , n54382 );
or ( n55500 , n55497 , n55498 , n55499 );
and ( n55501 , n54306 , n54383 );
and ( n55502 , n54383 , n54614 );
and ( n55503 , n54306 , n54614 );
or ( n55504 , n55501 , n55502 , n55503 );
xor ( n55505 , n55500 , n55504 );
and ( n55506 , n54385 , n54507 );
and ( n55507 , n54507 , n54613 );
and ( n55508 , n54385 , n54613 );
or ( n55509 , n55506 , n55507 , n55508 );
and ( n55510 , n54319 , n54323 );
and ( n55511 , n54323 , n54381 );
and ( n55512 , n54319 , n54381 );
or ( n55513 , n55510 , n55511 , n55512 );
and ( n55514 , n54389 , n54393 );
and ( n55515 , n54393 , n54506 );
and ( n55516 , n54389 , n54506 );
or ( n55517 , n55514 , n55515 , n55516 );
xor ( n55518 , n55513 , n55517 );
and ( n55519 , n54350 , n54354 );
and ( n55520 , n54354 , n54360 );
and ( n55521 , n54350 , n54360 );
or ( n55522 , n55519 , n55520 , n55521 );
and ( n55523 , n54328 , n54332 );
and ( n55524 , n54332 , n54380 );
and ( n55525 , n54328 , n54380 );
or ( n55526 , n55523 , n55524 , n55525 );
xor ( n55527 , n55522 , n55526 );
and ( n55528 , n54337 , n54341 );
and ( n55529 , n54341 , n54379 );
and ( n55530 , n54337 , n54379 );
or ( n55531 , n55528 , n55529 , n55530 );
and ( n55532 , n54402 , n54427 );
and ( n55533 , n54427 , n54467 );
and ( n55534 , n54402 , n54467 );
or ( n55535 , n55532 , n55533 , n55534 );
xor ( n55536 , n55531 , n55535 );
and ( n55537 , n54346 , n54361 );
and ( n55538 , n54361 , n54378 );
and ( n55539 , n54346 , n54378 );
or ( n55540 , n55537 , n55538 , n55539 );
and ( n55541 , n54406 , n54410 );
and ( n55542 , n54410 , n54426 );
and ( n55543 , n54406 , n54426 );
or ( n55544 , n55541 , n55542 , n55543 );
xor ( n55545 , n55540 , n55544 );
and ( n55546 , n54366 , n54371 );
and ( n55547 , n54371 , n54377 );
and ( n55548 , n54366 , n54377 );
or ( n55549 , n55546 , n55547 , n55548 );
and ( n55550 , n54356 , n54357 );
and ( n55551 , n54357 , n54359 );
and ( n55552 , n54356 , n54359 );
or ( n55553 , n55550 , n55551 , n55552 );
and ( n55554 , n54367 , n54368 );
and ( n55555 , n54368 , n54370 );
and ( n55556 , n54367 , n54370 );
or ( n55557 , n55554 , n55555 , n55556 );
xor ( n55558 , n55553 , n55557 );
and ( n55559 , n30695 , n3271 );
and ( n55560 , n31836 , n2981 );
xor ( n55561 , n55559 , n55560 );
and ( n55562 , n32649 , n2739 );
xor ( n55563 , n55561 , n55562 );
xor ( n55564 , n55558 , n55563 );
xor ( n55565 , n55549 , n55564 );
and ( n55566 , n54373 , n54374 );
and ( n55567 , n54374 , n54376 );
and ( n55568 , n54373 , n54376 );
or ( n55569 , n55566 , n55567 , n55568 );
and ( n55570 , n27361 , n4102 );
and ( n55571 , n28456 , n3749 );
xor ( n55572 , n55570 , n55571 );
and ( n55573 , n29559 , n3495 );
xor ( n55574 , n55572 , n55573 );
xor ( n55575 , n55569 , n55574 );
and ( n55576 , n24214 , n5103 );
and ( n55577 , n25243 , n4730 );
xor ( n55578 , n55576 , n55577 );
and ( n55579 , n26296 , n4403 );
xor ( n55580 , n55578 , n55579 );
xor ( n55581 , n55575 , n55580 );
xor ( n55582 , n55565 , n55581 );
xor ( n55583 , n55545 , n55582 );
xor ( n55584 , n55536 , n55583 );
xor ( n55585 , n55527 , n55584 );
xor ( n55586 , n55518 , n55585 );
xor ( n55587 , n55509 , n55586 );
and ( n55588 , n54583 , n54612 );
and ( n55589 , n54512 , n54513 );
and ( n55590 , n54513 , n54582 );
and ( n55591 , n54512 , n54582 );
or ( n55592 , n55589 , n55590 , n55591 );
and ( n55593 , n54398 , n54468 );
and ( n55594 , n54468 , n54505 );
and ( n55595 , n54398 , n54505 );
or ( n55596 , n55593 , n55594 , n55595 );
xor ( n55597 , n55592 , n55596 );
and ( n55598 , n54473 , n54477 );
and ( n55599 , n54477 , n54504 );
and ( n55600 , n54473 , n54504 );
or ( n55601 , n55598 , n55599 , n55600 );
and ( n55602 , n54432 , n54448 );
and ( n55603 , n54448 , n54466 );
and ( n55604 , n54432 , n54466 );
or ( n55605 , n55602 , n55603 , n55604 );
and ( n55606 , n54415 , n54419 );
and ( n55607 , n54419 , n54425 );
and ( n55608 , n54415 , n54425 );
or ( n55609 , n55606 , n55607 , n55608 );
and ( n55610 , n54436 , n54441 );
and ( n55611 , n54441 , n54447 );
and ( n55612 , n54436 , n54447 );
or ( n55613 , n55610 , n55611 , n55612 );
xor ( n55614 , n55609 , n55613 );
and ( n55615 , n54421 , n54422 );
and ( n55616 , n54422 , n54424 );
and ( n55617 , n54421 , n54424 );
or ( n55618 , n55615 , n55616 , n55617 );
and ( n55619 , n54437 , n54438 );
and ( n55620 , n54438 , n54440 );
and ( n55621 , n54437 , n54440 );
or ( n55622 , n55619 , n55620 , n55621 );
xor ( n55623 , n55618 , n55622 );
and ( n55624 , n21216 , n6132 );
and ( n55625 , n22186 , n5765 );
xor ( n55626 , n55624 , n55625 );
and ( n55627 , n22892 , n5408 );
xor ( n55628 , n55626 , n55627 );
xor ( n55629 , n55623 , n55628 );
xor ( n55630 , n55614 , n55629 );
xor ( n55631 , n55605 , n55630 );
and ( n55632 , n54453 , n54459 );
and ( n55633 , n54459 , n54465 );
and ( n55634 , n54453 , n54465 );
or ( n55635 , n55632 , n55633 , n55634 );
and ( n55636 , n54443 , n54444 );
and ( n55637 , n54444 , n54446 );
and ( n55638 , n54443 , n54446 );
or ( n55639 , n55636 , n55637 , n55638 );
and ( n55640 , n18144 , n7310 );
and ( n55641 , n19324 , n6971 );
xor ( n55642 , n55640 , n55641 );
and ( n55643 , n20233 , n6504 );
xor ( n55644 , n55642 , n55643 );
xor ( n55645 , n55639 , n55644 );
and ( n55646 , n15758 , n8669 );
and ( n55647 , n16637 , n8243 );
xor ( n55648 , n55646 , n55647 );
and ( n55649 , n17512 , n7662 );
xor ( n55650 , n55648 , n55649 );
xor ( n55651 , n55645 , n55650 );
xor ( n55652 , n55635 , n55651 );
and ( n55653 , n54461 , n54462 );
and ( n55654 , n54462 , n54464 );
and ( n55655 , n54461 , n54464 );
or ( n55656 , n55653 , n55654 , n55655 );
and ( n55657 , n54492 , n54493 );
and ( n55658 , n54493 , n54495 );
and ( n55659 , n54492 , n54495 );
or ( n55660 , n55657 , n55658 , n55659 );
xor ( n55661 , n55656 , n55660 );
and ( n55662 , n13322 , n10977 );
and ( n55663 , n14118 , n10239 );
xor ( n55664 , n55662 , n55663 );
and ( n55665 , n14938 , n9348 );
xor ( n55666 , n55664 , n55665 );
xor ( n55667 , n55661 , n55666 );
xor ( n55668 , n55652 , n55667 );
xor ( n55669 , n55631 , n55668 );
xor ( n55670 , n55601 , n55669 );
and ( n55671 , n54482 , n54486 );
and ( n55672 , n54486 , n54503 );
and ( n55673 , n54482 , n54503 );
or ( n55674 , n55671 , n55672 , n55673 );
and ( n55675 , n54522 , n54537 );
and ( n55676 , n54537 , n54554 );
and ( n55677 , n54522 , n54554 );
or ( n55678 , n55675 , n55676 , n55677 );
xor ( n55679 , n55674 , n55678 );
and ( n55680 , n54491 , n54496 );
and ( n55681 , n54496 , n54502 );
and ( n55682 , n54491 , n54502 );
or ( n55683 , n55680 , n55681 , n55682 );
and ( n55684 , n54526 , n54530 );
and ( n55685 , n54530 , n54536 );
and ( n55686 , n54526 , n54536 );
or ( n55687 , n55684 , n55685 , n55686 );
xor ( n55688 , n55683 , n55687 );
and ( n55689 , n54498 , n54499 );
and ( n55690 , n54499 , n54501 );
and ( n55691 , n54498 , n54501 );
or ( n55692 , n55689 , n55690 , n55691 );
and ( n55693 , n11015 , n13256 );
and ( n55694 , n11769 , n12531 );
xor ( n55695 , n55693 , n55694 );
and ( n55696 , n12320 , n11718 );
xor ( n55697 , n55695 , n55696 );
xor ( n55698 , n55692 , n55697 );
and ( n55699 , n8718 , n15691 );
and ( n55700 , n9400 , n14838 );
xor ( n55701 , n55699 , n55700 );
and ( n55702 , n10291 , n14044 );
xor ( n55703 , n55701 , n55702 );
xor ( n55704 , n55698 , n55703 );
xor ( n55705 , n55688 , n55704 );
xor ( n55706 , n55679 , n55705 );
xor ( n55707 , n55670 , n55706 );
xor ( n55708 , n55597 , n55707 );
xor ( n55709 , n55588 , n55708 );
and ( n55710 , n54518 , n54555 );
and ( n55711 , n54555 , n54581 );
and ( n55712 , n54518 , n54581 );
or ( n55713 , n55710 , n55711 , n55712 );
and ( n55714 , n54587 , n54611 );
xor ( n55715 , n55713 , n55714 );
and ( n55716 , n54560 , n54564 );
and ( n55717 , n54564 , n54580 );
and ( n55718 , n54560 , n54580 );
or ( n55719 , n55716 , n55717 , n55718 );
and ( n55720 , n54569 , n54573 );
and ( n55721 , n54573 , n54579 );
and ( n55722 , n54569 , n54579 );
or ( n55723 , n55720 , n55721 , n55722 );
and ( n55724 , n54592 , n54597 );
and ( n55725 , n54597 , n54603 );
and ( n55726 , n54592 , n54603 );
or ( n55727 , n55724 , n55725 , n55726 );
xor ( n55728 , n55723 , n55727 );
and ( n55729 , n54575 , n54576 );
and ( n55730 , n54576 , n54578 );
and ( n55731 , n54575 , n54578 );
or ( n55732 , n55729 , n55730 , n55731 );
and ( n55733 , n54593 , n54594 );
and ( n55734 , n54594 , n54596 );
and ( n55735 , n54593 , n54596 );
or ( n55736 , n55733 , n55734 , n55735 );
xor ( n55737 , n55732 , n55736 );
and ( n55738 , n4132 , n27296 );
and ( n55739 , n4438 , n26216 );
xor ( n55740 , n55738 , n55739 );
and ( n55741 , n4766 , n25163 );
xor ( n55742 , n55740 , n55741 );
xor ( n55743 , n55737 , n55742 );
xor ( n55744 , n55728 , n55743 );
xor ( n55745 , n55719 , n55744 );
and ( n55746 , n54542 , n54547 );
and ( n55747 , n54547 , n54553 );
and ( n55748 , n54542 , n54553 );
or ( n55749 , n55746 , n55747 , n55748 );
and ( n55750 , n54532 , n54533 );
and ( n55751 , n54533 , n54535 );
and ( n55752 , n54532 , n54535 );
or ( n55753 , n55750 , n55751 , n55752 );
and ( n55754 , n54543 , n54544 );
and ( n55755 , n54544 , n54546 );
and ( n55756 , n54543 , n54546 );
or ( n55757 , n55754 , n55755 , n55756 );
xor ( n55758 , n55753 , n55757 );
and ( n55759 , n7385 , n18407 );
and ( n55760 , n7808 , n17422 );
xor ( n55761 , n55759 , n55760 );
and ( n55762 , n8079 , n16550 );
xor ( n55763 , n55761 , n55762 );
xor ( n55764 , n55758 , n55763 );
xor ( n55765 , n55749 , n55764 );
and ( n55766 , n54549 , n54550 );
and ( n55767 , n54550 , n54552 );
and ( n55768 , n54549 , n54552 );
or ( n55769 , n55766 , n55767 , n55768 );
and ( n55770 , n6187 , n20976 );
and ( n55771 , n6569 , n20156 );
xor ( n55772 , n55770 , n55771 );
and ( n55773 , n6816 , n19222 );
xor ( n55774 , n55772 , n55773 );
xor ( n55775 , n55769 , n55774 );
and ( n55776 , n4959 , n24137 );
and ( n55777 , n5459 , n23075 );
xor ( n55778 , n55776 , n55777 );
and ( n55779 , n5819 , n22065 );
xor ( n55780 , n55778 , n55779 );
xor ( n55781 , n55775 , n55780 );
xor ( n55782 , n55765 , n55781 );
xor ( n55783 , n55745 , n55782 );
xor ( n55784 , n55715 , n55783 );
and ( n55785 , n54588 , n54604 );
and ( n55786 , n54604 , n54610 );
and ( n55787 , n54588 , n54610 );
or ( n55788 , n55785 , n55786 , n55787 );
and ( n55789 , n54606 , n54609 );
and ( n55790 , n54599 , n54600 );
and ( n55791 , n54600 , n54602 );
and ( n55792 , n54599 , n54602 );
or ( n55793 , n55790 , n55791 , n55792 );
and ( n55794 , n3182 , n30629 );
and ( n55795 , n3545 , n29508 );
xor ( n55796 , n55794 , n55795 );
and ( n55797 , n3801 , n28406 );
xor ( n55798 , n55796 , n55797 );
xor ( n55799 , n55793 , n55798 );
not ( n55800 , n2462 );
and ( n55801 , n34193 , n2462 );
nor ( n55802 , n55800 , n55801 );
and ( n55803 , n2779 , n32999 );
xor ( n55804 , n55802 , n55803 );
and ( n55805 , n3024 , n31761 );
xor ( n55806 , n55804 , n55805 );
xor ( n55807 , n55799 , n55806 );
xor ( n55808 , n55789 , n55807 );
xor ( n55809 , n55788 , n55808 );
xor ( n55810 , n55784 , n55809 );
xor ( n55811 , n55709 , n55810 );
xor ( n55812 , n55587 , n55811 );
xor ( n55813 , n55505 , n55812 );
xor ( n55814 , n55496 , n55813 );
and ( n55815 , n54289 , n54292 );
and ( n55816 , n54292 , n54616 );
and ( n55817 , n54289 , n54616 );
or ( n55818 , n55815 , n55816 , n55817 );
xor ( n55819 , n55814 , n55818 );
and ( n55820 , n54617 , n54621 );
and ( n55821 , n54622 , n54625 );
or ( n55822 , n55820 , n55821 );
xor ( n55823 , n55819 , n55822 );
buf ( n55824 , n55823 );
buf ( n55825 , n55824 );
not ( n55826 , n55825 );
nor ( n55827 , n55826 , n8739 );
xor ( n55828 , n55488 , n55827 );
and ( n55829 , n54285 , n54630 );
and ( n55830 , n54631 , n54634 );
or ( n55831 , n55829 , n55830 );
xor ( n55832 , n55828 , n55831 );
buf ( n55833 , n55832 );
buf ( n55834 , n55833 );
not ( n55835 , n55834 );
buf ( n55836 , n580 );
not ( n55837 , n55836 );
nor ( n55838 , n55835 , n55837 );
xor ( n55839 , n55114 , n55838 );
xor ( n55840 , n54646 , n55111 );
nor ( n55841 , n54638 , n55837 );
and ( n55842 , n55840 , n55841 );
xor ( n55843 , n55840 , n55841 );
xor ( n55844 , n54650 , n55109 );
nor ( n55845 , n53441 , n55837 );
and ( n55846 , n55844 , n55845 );
xor ( n55847 , n55844 , n55845 );
xor ( n55848 , n54654 , n55107 );
nor ( n55849 , n52247 , n55837 );
and ( n55850 , n55848 , n55849 );
xor ( n55851 , n55848 , n55849 );
xor ( n55852 , n54658 , n55105 );
nor ( n55853 , n51049 , n55837 );
and ( n55854 , n55852 , n55853 );
xor ( n55855 , n55852 , n55853 );
xor ( n55856 , n54662 , n55103 );
nor ( n55857 , n49850 , n55837 );
and ( n55858 , n55856 , n55857 );
xor ( n55859 , n55856 , n55857 );
xor ( n55860 , n54666 , n55101 );
nor ( n55861 , n48650 , n55837 );
and ( n55862 , n55860 , n55861 );
xor ( n55863 , n55860 , n55861 );
xor ( n55864 , n54670 , n55099 );
nor ( n55865 , n47449 , n55837 );
and ( n55866 , n55864 , n55865 );
xor ( n55867 , n55864 , n55865 );
xor ( n55868 , n54674 , n55097 );
nor ( n55869 , n46248 , n55837 );
and ( n55870 , n55868 , n55869 );
xor ( n55871 , n55868 , n55869 );
xor ( n55872 , n54678 , n55095 );
nor ( n55873 , n45047 , n55837 );
and ( n55874 , n55872 , n55873 );
xor ( n55875 , n55872 , n55873 );
xor ( n55876 , n54682 , n55093 );
nor ( n55877 , n43843 , n55837 );
and ( n55878 , n55876 , n55877 );
xor ( n55879 , n55876 , n55877 );
xor ( n55880 , n54686 , n55091 );
nor ( n55881 , n42641 , n55837 );
and ( n55882 , n55880 , n55881 );
xor ( n55883 , n55880 , n55881 );
xor ( n55884 , n54690 , n55089 );
nor ( n55885 , n41437 , n55837 );
and ( n55886 , n55884 , n55885 );
xor ( n55887 , n55884 , n55885 );
xor ( n55888 , n54694 , n55087 );
nor ( n55889 , n40232 , n55837 );
and ( n55890 , n55888 , n55889 );
xor ( n55891 , n55888 , n55889 );
xor ( n55892 , n54698 , n55085 );
nor ( n55893 , n39027 , n55837 );
and ( n55894 , n55892 , n55893 );
xor ( n55895 , n55892 , n55893 );
xor ( n55896 , n54702 , n55083 );
nor ( n55897 , n37825 , n55837 );
and ( n55898 , n55896 , n55897 );
xor ( n55899 , n55896 , n55897 );
xor ( n55900 , n54706 , n55081 );
nor ( n55901 , n36620 , n55837 );
and ( n55902 , n55900 , n55901 );
xor ( n55903 , n55900 , n55901 );
xor ( n55904 , n54710 , n55079 );
nor ( n55905 , n35419 , n55837 );
and ( n55906 , n55904 , n55905 );
xor ( n55907 , n55904 , n55905 );
xor ( n55908 , n54714 , n55077 );
nor ( n55909 , n34224 , n55837 );
and ( n55910 , n55908 , n55909 );
xor ( n55911 , n55908 , n55909 );
xor ( n55912 , n54718 , n55075 );
nor ( n55913 , n33033 , n55837 );
and ( n55914 , n55912 , n55913 );
xor ( n55915 , n55912 , n55913 );
xor ( n55916 , n54722 , n55073 );
nor ( n55917 , n31867 , n55837 );
and ( n55918 , n55916 , n55917 );
xor ( n55919 , n55916 , n55917 );
xor ( n55920 , n54726 , n55071 );
nor ( n55921 , n30725 , n55837 );
and ( n55922 , n55920 , n55921 );
xor ( n55923 , n55920 , n55921 );
xor ( n55924 , n54730 , n55069 );
nor ( n55925 , n29596 , n55837 );
and ( n55926 , n55924 , n55925 );
xor ( n55927 , n55924 , n55925 );
xor ( n55928 , n54734 , n55067 );
nor ( n55929 , n28487 , n55837 );
and ( n55930 , n55928 , n55929 );
xor ( n55931 , n55928 , n55929 );
xor ( n55932 , n54738 , n55065 );
nor ( n55933 , n27397 , n55837 );
and ( n55934 , n55932 , n55933 );
xor ( n55935 , n55932 , n55933 );
xor ( n55936 , n54742 , n55063 );
nor ( n55937 , n26326 , n55837 );
and ( n55938 , n55936 , n55937 );
xor ( n55939 , n55936 , n55937 );
xor ( n55940 , n54746 , n55061 );
nor ( n55941 , n25272 , n55837 );
and ( n55942 , n55940 , n55941 );
xor ( n55943 , n55940 , n55941 );
xor ( n55944 , n54750 , n55059 );
nor ( n55945 , n24242 , n55837 );
and ( n55946 , n55944 , n55945 );
xor ( n55947 , n55944 , n55945 );
xor ( n55948 , n54754 , n55057 );
nor ( n55949 , n23225 , n55837 );
and ( n55950 , n55948 , n55949 );
xor ( n55951 , n55948 , n55949 );
xor ( n55952 , n54758 , n55055 );
nor ( n55953 , n22231 , n55837 );
and ( n55954 , n55952 , n55953 );
xor ( n55955 , n55952 , n55953 );
xor ( n55956 , n54762 , n55053 );
nor ( n55957 , n21258 , n55837 );
and ( n55958 , n55956 , n55957 );
xor ( n55959 , n55956 , n55957 );
xor ( n55960 , n54766 , n55051 );
nor ( n55961 , n20303 , n55837 );
and ( n55962 , n55960 , n55961 );
xor ( n55963 , n55960 , n55961 );
xor ( n55964 , n54770 , n55049 );
nor ( n55965 , n19365 , n55837 );
and ( n55966 , n55964 , n55965 );
xor ( n55967 , n55964 , n55965 );
xor ( n55968 , n54774 , n55047 );
nor ( n55969 , n18448 , n55837 );
and ( n55970 , n55968 , n55969 );
xor ( n55971 , n55968 , n55969 );
xor ( n55972 , n54778 , n55045 );
nor ( n55973 , n17548 , n55837 );
and ( n55974 , n55972 , n55973 );
xor ( n55975 , n55972 , n55973 );
xor ( n55976 , n54782 , n55043 );
nor ( n55977 , n16669 , n55837 );
and ( n55978 , n55976 , n55977 );
xor ( n55979 , n55976 , n55977 );
xor ( n55980 , n54786 , n55041 );
nor ( n55981 , n15809 , n55837 );
and ( n55982 , n55980 , n55981 );
xor ( n55983 , n55980 , n55981 );
xor ( n55984 , n54790 , n55039 );
nor ( n55985 , n14968 , n55837 );
and ( n55986 , n55984 , n55985 );
xor ( n55987 , n55984 , n55985 );
xor ( n55988 , n54794 , n55037 );
nor ( n55989 , n14147 , n55837 );
and ( n55990 , n55988 , n55989 );
xor ( n55991 , n55988 , n55989 );
xor ( n55992 , n54798 , n55035 );
nor ( n55993 , n13349 , n55837 );
and ( n55994 , n55992 , n55993 );
xor ( n55995 , n55992 , n55993 );
xor ( n55996 , n54802 , n55033 );
nor ( n55997 , n12564 , n55837 );
and ( n55998 , n55996 , n55997 );
xor ( n55999 , n55996 , n55997 );
xor ( n56000 , n54806 , n55031 );
nor ( n56001 , n11799 , n55837 );
and ( n56002 , n56000 , n56001 );
xor ( n56003 , n56000 , n56001 );
xor ( n56004 , n54810 , n55029 );
nor ( n56005 , n11050 , n55837 );
and ( n56006 , n56004 , n56005 );
xor ( n56007 , n56004 , n56005 );
xor ( n56008 , n54814 , n55027 );
nor ( n56009 , n10321 , n55837 );
and ( n56010 , n56008 , n56009 );
xor ( n56011 , n56008 , n56009 );
xor ( n56012 , n54818 , n55025 );
nor ( n56013 , n9429 , n55837 );
and ( n56014 , n56012 , n56013 );
xor ( n56015 , n56012 , n56013 );
xor ( n56016 , n54822 , n55023 );
nor ( n56017 , n8949 , n55837 );
and ( n56018 , n56016 , n56017 );
xor ( n56019 , n56016 , n56017 );
xor ( n56020 , n54826 , n55021 );
nor ( n56021 , n9437 , n55837 );
and ( n56022 , n56020 , n56021 );
xor ( n56023 , n56020 , n56021 );
xor ( n56024 , n54830 , n55019 );
nor ( n56025 , n9446 , n55837 );
and ( n56026 , n56024 , n56025 );
xor ( n56027 , n56024 , n56025 );
xor ( n56028 , n54834 , n55017 );
nor ( n56029 , n9455 , n55837 );
and ( n56030 , n56028 , n56029 );
xor ( n56031 , n56028 , n56029 );
xor ( n56032 , n54838 , n55015 );
nor ( n56033 , n9464 , n55837 );
and ( n56034 , n56032 , n56033 );
xor ( n56035 , n56032 , n56033 );
xor ( n56036 , n54842 , n55013 );
nor ( n56037 , n9473 , n55837 );
and ( n56038 , n56036 , n56037 );
xor ( n56039 , n56036 , n56037 );
xor ( n56040 , n54846 , n55011 );
nor ( n56041 , n9482 , n55837 );
and ( n56042 , n56040 , n56041 );
xor ( n56043 , n56040 , n56041 );
xor ( n56044 , n54850 , n55009 );
nor ( n56045 , n9491 , n55837 );
and ( n56046 , n56044 , n56045 );
xor ( n56047 , n56044 , n56045 );
xor ( n56048 , n54854 , n55007 );
nor ( n56049 , n9500 , n55837 );
and ( n56050 , n56048 , n56049 );
xor ( n56051 , n56048 , n56049 );
xor ( n56052 , n54858 , n55005 );
nor ( n56053 , n9509 , n55837 );
and ( n56054 , n56052 , n56053 );
xor ( n56055 , n56052 , n56053 );
xor ( n56056 , n54862 , n55003 );
nor ( n56057 , n9518 , n55837 );
and ( n56058 , n56056 , n56057 );
xor ( n56059 , n56056 , n56057 );
xor ( n56060 , n54866 , n55001 );
nor ( n56061 , n9527 , n55837 );
and ( n56062 , n56060 , n56061 );
xor ( n56063 , n56060 , n56061 );
xor ( n56064 , n54870 , n54999 );
nor ( n56065 , n9536 , n55837 );
and ( n56066 , n56064 , n56065 );
xor ( n56067 , n56064 , n56065 );
xor ( n56068 , n54874 , n54997 );
nor ( n56069 , n9545 , n55837 );
and ( n56070 , n56068 , n56069 );
xor ( n56071 , n56068 , n56069 );
xor ( n56072 , n54878 , n54995 );
nor ( n56073 , n9554 , n55837 );
and ( n56074 , n56072 , n56073 );
xor ( n56075 , n56072 , n56073 );
xor ( n56076 , n54882 , n54993 );
nor ( n56077 , n9563 , n55837 );
and ( n56078 , n56076 , n56077 );
xor ( n56079 , n56076 , n56077 );
xor ( n56080 , n54886 , n54991 );
nor ( n56081 , n9572 , n55837 );
and ( n56082 , n56080 , n56081 );
xor ( n56083 , n56080 , n56081 );
xor ( n56084 , n54890 , n54989 );
nor ( n56085 , n9581 , n55837 );
and ( n56086 , n56084 , n56085 );
xor ( n56087 , n56084 , n56085 );
xor ( n56088 , n54894 , n54987 );
nor ( n56089 , n9590 , n55837 );
and ( n56090 , n56088 , n56089 );
xor ( n56091 , n56088 , n56089 );
xor ( n56092 , n54898 , n54985 );
nor ( n56093 , n9599 , n55837 );
and ( n56094 , n56092 , n56093 );
xor ( n56095 , n56092 , n56093 );
xor ( n56096 , n54902 , n54983 );
nor ( n56097 , n9608 , n55837 );
and ( n56098 , n56096 , n56097 );
xor ( n56099 , n56096 , n56097 );
xor ( n56100 , n54906 , n54981 );
nor ( n56101 , n9617 , n55837 );
and ( n56102 , n56100 , n56101 );
xor ( n56103 , n56100 , n56101 );
xor ( n56104 , n54910 , n54979 );
nor ( n56105 , n9626 , n55837 );
and ( n56106 , n56104 , n56105 );
xor ( n56107 , n56104 , n56105 );
xor ( n56108 , n54914 , n54977 );
nor ( n56109 , n9635 , n55837 );
and ( n56110 , n56108 , n56109 );
xor ( n56111 , n56108 , n56109 );
xor ( n56112 , n54918 , n54975 );
nor ( n56113 , n9644 , n55837 );
and ( n56114 , n56112 , n56113 );
xor ( n56115 , n56112 , n56113 );
xor ( n56116 , n54922 , n54973 );
nor ( n56117 , n9653 , n55837 );
and ( n56118 , n56116 , n56117 );
xor ( n56119 , n56116 , n56117 );
xor ( n56120 , n54926 , n54971 );
nor ( n56121 , n9662 , n55837 );
and ( n56122 , n56120 , n56121 );
xor ( n56123 , n56120 , n56121 );
xor ( n56124 , n54930 , n54969 );
nor ( n56125 , n9671 , n55837 );
and ( n56126 , n56124 , n56125 );
xor ( n56127 , n56124 , n56125 );
xor ( n56128 , n54934 , n54967 );
nor ( n56129 , n9680 , n55837 );
and ( n56130 , n56128 , n56129 );
xor ( n56131 , n56128 , n56129 );
xor ( n56132 , n54938 , n54965 );
nor ( n56133 , n9689 , n55837 );
and ( n56134 , n56132 , n56133 );
xor ( n56135 , n56132 , n56133 );
xor ( n56136 , n54942 , n54963 );
nor ( n56137 , n9698 , n55837 );
and ( n56138 , n56136 , n56137 );
xor ( n56139 , n56136 , n56137 );
xor ( n56140 , n54946 , n54961 );
nor ( n56141 , n9707 , n55837 );
and ( n56142 , n56140 , n56141 );
xor ( n56143 , n56140 , n56141 );
xor ( n56144 , n54950 , n54959 );
nor ( n56145 , n9716 , n55837 );
and ( n56146 , n56144 , n56145 );
xor ( n56147 , n56144 , n56145 );
xor ( n56148 , n54954 , n54957 );
nor ( n56149 , n9725 , n55837 );
and ( n56150 , n56148 , n56149 );
xor ( n56151 , n56148 , n56149 );
xor ( n56152 , n54955 , n54956 );
nor ( n56153 , n9734 , n55837 );
and ( n56154 , n56152 , n56153 );
xor ( n56155 , n56152 , n56153 );
nor ( n56156 , n9752 , n54640 );
nor ( n56157 , n9743 , n55837 );
and ( n56158 , n56156 , n56157 );
and ( n56159 , n56155 , n56158 );
or ( n56160 , n56154 , n56159 );
and ( n56161 , n56151 , n56160 );
or ( n56162 , n56150 , n56161 );
and ( n56163 , n56147 , n56162 );
or ( n56164 , n56146 , n56163 );
and ( n56165 , n56143 , n56164 );
or ( n56166 , n56142 , n56165 );
and ( n56167 , n56139 , n56166 );
or ( n56168 , n56138 , n56167 );
and ( n56169 , n56135 , n56168 );
or ( n56170 , n56134 , n56169 );
and ( n56171 , n56131 , n56170 );
or ( n56172 , n56130 , n56171 );
and ( n56173 , n56127 , n56172 );
or ( n56174 , n56126 , n56173 );
and ( n56175 , n56123 , n56174 );
or ( n56176 , n56122 , n56175 );
and ( n56177 , n56119 , n56176 );
or ( n56178 , n56118 , n56177 );
and ( n56179 , n56115 , n56178 );
or ( n56180 , n56114 , n56179 );
and ( n56181 , n56111 , n56180 );
or ( n56182 , n56110 , n56181 );
and ( n56183 , n56107 , n56182 );
or ( n56184 , n56106 , n56183 );
and ( n56185 , n56103 , n56184 );
or ( n56186 , n56102 , n56185 );
and ( n56187 , n56099 , n56186 );
or ( n56188 , n56098 , n56187 );
and ( n56189 , n56095 , n56188 );
or ( n56190 , n56094 , n56189 );
and ( n56191 , n56091 , n56190 );
or ( n56192 , n56090 , n56191 );
and ( n56193 , n56087 , n56192 );
or ( n56194 , n56086 , n56193 );
and ( n56195 , n56083 , n56194 );
or ( n56196 , n56082 , n56195 );
and ( n56197 , n56079 , n56196 );
or ( n56198 , n56078 , n56197 );
and ( n56199 , n56075 , n56198 );
or ( n56200 , n56074 , n56199 );
and ( n56201 , n56071 , n56200 );
or ( n56202 , n56070 , n56201 );
and ( n56203 , n56067 , n56202 );
or ( n56204 , n56066 , n56203 );
and ( n56205 , n56063 , n56204 );
or ( n56206 , n56062 , n56205 );
and ( n56207 , n56059 , n56206 );
or ( n56208 , n56058 , n56207 );
and ( n56209 , n56055 , n56208 );
or ( n56210 , n56054 , n56209 );
and ( n56211 , n56051 , n56210 );
or ( n56212 , n56050 , n56211 );
and ( n56213 , n56047 , n56212 );
or ( n56214 , n56046 , n56213 );
and ( n56215 , n56043 , n56214 );
or ( n56216 , n56042 , n56215 );
and ( n56217 , n56039 , n56216 );
or ( n56218 , n56038 , n56217 );
and ( n56219 , n56035 , n56218 );
or ( n56220 , n56034 , n56219 );
and ( n56221 , n56031 , n56220 );
or ( n56222 , n56030 , n56221 );
and ( n56223 , n56027 , n56222 );
or ( n56224 , n56026 , n56223 );
and ( n56225 , n56023 , n56224 );
or ( n56226 , n56022 , n56225 );
and ( n56227 , n56019 , n56226 );
or ( n56228 , n56018 , n56227 );
and ( n56229 , n56015 , n56228 );
or ( n56230 , n56014 , n56229 );
and ( n56231 , n56011 , n56230 );
or ( n56232 , n56010 , n56231 );
and ( n56233 , n56007 , n56232 );
or ( n56234 , n56006 , n56233 );
and ( n56235 , n56003 , n56234 );
or ( n56236 , n56002 , n56235 );
and ( n56237 , n55999 , n56236 );
or ( n56238 , n55998 , n56237 );
and ( n56239 , n55995 , n56238 );
or ( n56240 , n55994 , n56239 );
and ( n56241 , n55991 , n56240 );
or ( n56242 , n55990 , n56241 );
and ( n56243 , n55987 , n56242 );
or ( n56244 , n55986 , n56243 );
and ( n56245 , n55983 , n56244 );
or ( n56246 , n55982 , n56245 );
and ( n56247 , n55979 , n56246 );
or ( n56248 , n55978 , n56247 );
and ( n56249 , n55975 , n56248 );
or ( n56250 , n55974 , n56249 );
and ( n56251 , n55971 , n56250 );
or ( n56252 , n55970 , n56251 );
and ( n56253 , n55967 , n56252 );
or ( n56254 , n55966 , n56253 );
and ( n56255 , n55963 , n56254 );
or ( n56256 , n55962 , n56255 );
and ( n56257 , n55959 , n56256 );
or ( n56258 , n55958 , n56257 );
and ( n56259 , n55955 , n56258 );
or ( n56260 , n55954 , n56259 );
and ( n56261 , n55951 , n56260 );
or ( n56262 , n55950 , n56261 );
and ( n56263 , n55947 , n56262 );
or ( n56264 , n55946 , n56263 );
and ( n56265 , n55943 , n56264 );
or ( n56266 , n55942 , n56265 );
and ( n56267 , n55939 , n56266 );
or ( n56268 , n55938 , n56267 );
and ( n56269 , n55935 , n56268 );
or ( n56270 , n55934 , n56269 );
and ( n56271 , n55931 , n56270 );
or ( n56272 , n55930 , n56271 );
and ( n56273 , n55927 , n56272 );
or ( n56274 , n55926 , n56273 );
and ( n56275 , n55923 , n56274 );
or ( n56276 , n55922 , n56275 );
and ( n56277 , n55919 , n56276 );
or ( n56278 , n55918 , n56277 );
and ( n56279 , n55915 , n56278 );
or ( n56280 , n55914 , n56279 );
and ( n56281 , n55911 , n56280 );
or ( n56282 , n55910 , n56281 );
and ( n56283 , n55907 , n56282 );
or ( n56284 , n55906 , n56283 );
and ( n56285 , n55903 , n56284 );
or ( n56286 , n55902 , n56285 );
and ( n56287 , n55899 , n56286 );
or ( n56288 , n55898 , n56287 );
and ( n56289 , n55895 , n56288 );
or ( n56290 , n55894 , n56289 );
and ( n56291 , n55891 , n56290 );
or ( n56292 , n55890 , n56291 );
and ( n56293 , n55887 , n56292 );
or ( n56294 , n55886 , n56293 );
and ( n56295 , n55883 , n56294 );
or ( n56296 , n55882 , n56295 );
and ( n56297 , n55879 , n56296 );
or ( n56298 , n55878 , n56297 );
and ( n56299 , n55875 , n56298 );
or ( n56300 , n55874 , n56299 );
and ( n56301 , n55871 , n56300 );
or ( n56302 , n55870 , n56301 );
and ( n56303 , n55867 , n56302 );
or ( n56304 , n55866 , n56303 );
and ( n56305 , n55863 , n56304 );
or ( n56306 , n55862 , n56305 );
and ( n56307 , n55859 , n56306 );
or ( n56308 , n55858 , n56307 );
and ( n56309 , n55855 , n56308 );
or ( n56310 , n55854 , n56309 );
and ( n56311 , n55851 , n56310 );
or ( n56312 , n55850 , n56311 );
and ( n56313 , n55847 , n56312 );
or ( n56314 , n55846 , n56313 );
and ( n56315 , n55843 , n56314 );
or ( n56316 , n55842 , n56315 );
xor ( n56317 , n55839 , n56316 );
and ( n56318 , n33403 , n2796 );
nor ( n56319 , n2797 , n56318 );
nor ( n56320 , n3043 , n32231 );
xor ( n56321 , n56319 , n56320 );
and ( n56322 , n55116 , n55117 );
and ( n56323 , n55118 , n55121 );
or ( n56324 , n56322 , n56323 );
xor ( n56325 , n56321 , n56324 );
nor ( n56326 , n3300 , n31083 );
xor ( n56327 , n56325 , n56326 );
and ( n56328 , n55122 , n55123 );
and ( n56329 , n55124 , n55127 );
or ( n56330 , n56328 , n56329 );
xor ( n56331 , n56327 , n56330 );
nor ( n56332 , n3570 , n29948 );
xor ( n56333 , n56331 , n56332 );
and ( n56334 , n55128 , n55129 );
and ( n56335 , n55130 , n55133 );
or ( n56336 , n56334 , n56335 );
xor ( n56337 , n56333 , n56336 );
nor ( n56338 , n3853 , n28833 );
xor ( n56339 , n56337 , n56338 );
and ( n56340 , n55134 , n55135 );
and ( n56341 , n55136 , n55139 );
or ( n56342 , n56340 , n56341 );
xor ( n56343 , n56339 , n56342 );
nor ( n56344 , n4151 , n27737 );
xor ( n56345 , n56343 , n56344 );
and ( n56346 , n55140 , n55141 );
and ( n56347 , n55142 , n55145 );
or ( n56348 , n56346 , n56347 );
xor ( n56349 , n56345 , n56348 );
nor ( n56350 , n4458 , n26660 );
xor ( n56351 , n56349 , n56350 );
and ( n56352 , n55146 , n55147 );
and ( n56353 , n55148 , n55151 );
or ( n56354 , n56352 , n56353 );
xor ( n56355 , n56351 , n56354 );
nor ( n56356 , n4786 , n25600 );
xor ( n56357 , n56355 , n56356 );
and ( n56358 , n55152 , n55153 );
and ( n56359 , n55154 , n55157 );
or ( n56360 , n56358 , n56359 );
xor ( n56361 , n56357 , n56360 );
nor ( n56362 , n5126 , n24564 );
xor ( n56363 , n56361 , n56362 );
and ( n56364 , n55158 , n55159 );
and ( n56365 , n55160 , n55163 );
or ( n56366 , n56364 , n56365 );
xor ( n56367 , n56363 , n56366 );
nor ( n56368 , n5477 , n23541 );
xor ( n56369 , n56367 , n56368 );
and ( n56370 , n55164 , n55165 );
and ( n56371 , n55166 , n55169 );
or ( n56372 , n56370 , n56371 );
xor ( n56373 , n56369 , n56372 );
nor ( n56374 , n5838 , n22541 );
xor ( n56375 , n56373 , n56374 );
and ( n56376 , n55170 , n55171 );
and ( n56377 , n55172 , n55175 );
or ( n56378 , n56376 , n56377 );
xor ( n56379 , n56375 , n56378 );
nor ( n56380 , n6212 , n21562 );
xor ( n56381 , n56379 , n56380 );
and ( n56382 , n55176 , n55177 );
and ( n56383 , n55178 , n55181 );
or ( n56384 , n56382 , n56383 );
xor ( n56385 , n56381 , n56384 );
nor ( n56386 , n6596 , n20601 );
xor ( n56387 , n56385 , n56386 );
and ( n56388 , n55182 , n55183 );
and ( n56389 , n55184 , n55187 );
or ( n56390 , n56388 , n56389 );
xor ( n56391 , n56387 , n56390 );
nor ( n56392 , n6997 , n19657 );
xor ( n56393 , n56391 , n56392 );
and ( n56394 , n55188 , n55189 );
and ( n56395 , n55190 , n55193 );
or ( n56396 , n56394 , n56395 );
xor ( n56397 , n56393 , n56396 );
nor ( n56398 , n7413 , n18734 );
xor ( n56399 , n56397 , n56398 );
and ( n56400 , n55194 , n55195 );
and ( n56401 , n55196 , n55199 );
or ( n56402 , n56400 , n56401 );
xor ( n56403 , n56399 , n56402 );
nor ( n56404 , n7841 , n17828 );
xor ( n56405 , n56403 , n56404 );
and ( n56406 , n55200 , n55201 );
and ( n56407 , n55202 , n55205 );
or ( n56408 , n56406 , n56407 );
xor ( n56409 , n56405 , n56408 );
nor ( n56410 , n8281 , n16943 );
xor ( n56411 , n56409 , n56410 );
and ( n56412 , n55206 , n55207 );
and ( n56413 , n55208 , n55211 );
or ( n56414 , n56412 , n56413 );
xor ( n56415 , n56411 , n56414 );
nor ( n56416 , n8737 , n16077 );
xor ( n56417 , n56415 , n56416 );
and ( n56418 , n55212 , n55213 );
and ( n56419 , n55214 , n55217 );
or ( n56420 , n56418 , n56419 );
xor ( n56421 , n56417 , n56420 );
nor ( n56422 , n9420 , n15230 );
xor ( n56423 , n56421 , n56422 );
and ( n56424 , n55218 , n55219 );
and ( n56425 , n55220 , n55223 );
or ( n56426 , n56424 , n56425 );
xor ( n56427 , n56423 , n56426 );
nor ( n56428 , n10312 , n14403 );
xor ( n56429 , n56427 , n56428 );
and ( n56430 , n55224 , n55225 );
and ( n56431 , n55226 , n55229 );
or ( n56432 , n56430 , n56431 );
xor ( n56433 , n56429 , n56432 );
nor ( n56434 , n11041 , n13599 );
xor ( n56435 , n56433 , n56434 );
and ( n56436 , n55230 , n55231 );
and ( n56437 , n55232 , n55235 );
or ( n56438 , n56436 , n56437 );
xor ( n56439 , n56435 , n56438 );
nor ( n56440 , n11790 , n12808 );
xor ( n56441 , n56439 , n56440 );
and ( n56442 , n55236 , n55237 );
and ( n56443 , n55238 , n55241 );
or ( n56444 , n56442 , n56443 );
xor ( n56445 , n56441 , n56444 );
nor ( n56446 , n12555 , n12037 );
xor ( n56447 , n56445 , n56446 );
and ( n56448 , n55242 , n55243 );
and ( n56449 , n55244 , n55247 );
or ( n56450 , n56448 , n56449 );
xor ( n56451 , n56447 , n56450 );
nor ( n56452 , n13340 , n11282 );
xor ( n56453 , n56451 , n56452 );
and ( n56454 , n55248 , n55249 );
and ( n56455 , n55250 , n55253 );
or ( n56456 , n56454 , n56455 );
xor ( n56457 , n56453 , n56456 );
nor ( n56458 , n14138 , n10547 );
xor ( n56459 , n56457 , n56458 );
and ( n56460 , n55254 , n55255 );
and ( n56461 , n55256 , n55259 );
or ( n56462 , n56460 , n56461 );
xor ( n56463 , n56459 , n56462 );
nor ( n56464 , n14959 , n9829 );
xor ( n56465 , n56463 , n56464 );
and ( n56466 , n55260 , n55261 );
and ( n56467 , n55262 , n55265 );
or ( n56468 , n56466 , n56467 );
xor ( n56469 , n56465 , n56468 );
nor ( n56470 , n15800 , n8955 );
xor ( n56471 , n56469 , n56470 );
and ( n56472 , n55266 , n55267 );
and ( n56473 , n55268 , n55271 );
or ( n56474 , n56472 , n56473 );
xor ( n56475 , n56471 , n56474 );
nor ( n56476 , n16660 , n603 );
xor ( n56477 , n56475 , n56476 );
and ( n56478 , n55272 , n55273 );
and ( n56479 , n55274 , n55277 );
or ( n56480 , n56478 , n56479 );
xor ( n56481 , n56477 , n56480 );
nor ( n56482 , n17539 , n652 );
xor ( n56483 , n56481 , n56482 );
and ( n56484 , n55278 , n55279 );
and ( n56485 , n55280 , n55283 );
or ( n56486 , n56484 , n56485 );
xor ( n56487 , n56483 , n56486 );
nor ( n56488 , n18439 , n624 );
xor ( n56489 , n56487 , n56488 );
and ( n56490 , n55284 , n55285 );
and ( n56491 , n55286 , n55289 );
or ( n56492 , n56490 , n56491 );
xor ( n56493 , n56489 , n56492 );
nor ( n56494 , n19356 , n648 );
xor ( n56495 , n56493 , n56494 );
and ( n56496 , n55290 , n55291 );
and ( n56497 , n55292 , n55295 );
or ( n56498 , n56496 , n56497 );
xor ( n56499 , n56495 , n56498 );
nor ( n56500 , n20294 , n686 );
xor ( n56501 , n56499 , n56500 );
and ( n56502 , n55296 , n55297 );
and ( n56503 , n55298 , n55301 );
or ( n56504 , n56502 , n56503 );
xor ( n56505 , n56501 , n56504 );
nor ( n56506 , n21249 , n735 );
xor ( n56507 , n56505 , n56506 );
and ( n56508 , n55302 , n55303 );
and ( n56509 , n55304 , n55307 );
or ( n56510 , n56508 , n56509 );
xor ( n56511 , n56507 , n56510 );
nor ( n56512 , n22222 , n798 );
xor ( n56513 , n56511 , n56512 );
and ( n56514 , n55308 , n55309 );
and ( n56515 , n55310 , n55313 );
or ( n56516 , n56514 , n56515 );
xor ( n56517 , n56513 , n56516 );
nor ( n56518 , n23216 , n870 );
xor ( n56519 , n56517 , n56518 );
and ( n56520 , n55314 , n55315 );
and ( n56521 , n55316 , n55319 );
or ( n56522 , n56520 , n56521 );
xor ( n56523 , n56519 , n56522 );
nor ( n56524 , n24233 , n960 );
xor ( n56525 , n56523 , n56524 );
and ( n56526 , n55320 , n55321 );
and ( n56527 , n55322 , n55325 );
or ( n56528 , n56526 , n56527 );
xor ( n56529 , n56525 , n56528 );
nor ( n56530 , n25263 , n1064 );
xor ( n56531 , n56529 , n56530 );
and ( n56532 , n55326 , n55327 );
and ( n56533 , n55328 , n55331 );
or ( n56534 , n56532 , n56533 );
xor ( n56535 , n56531 , n56534 );
nor ( n56536 , n26317 , n1178 );
xor ( n56537 , n56535 , n56536 );
and ( n56538 , n55332 , n55333 );
and ( n56539 , n55334 , n55337 );
or ( n56540 , n56538 , n56539 );
xor ( n56541 , n56537 , n56540 );
nor ( n56542 , n27388 , n1305 );
xor ( n56543 , n56541 , n56542 );
and ( n56544 , n55338 , n55339 );
and ( n56545 , n55340 , n55343 );
or ( n56546 , n56544 , n56545 );
xor ( n56547 , n56543 , n56546 );
nor ( n56548 , n28478 , n1447 );
xor ( n56549 , n56547 , n56548 );
and ( n56550 , n55344 , n55345 );
and ( n56551 , n55346 , n55349 );
or ( n56552 , n56550 , n56551 );
xor ( n56553 , n56549 , n56552 );
nor ( n56554 , n29587 , n1600 );
xor ( n56555 , n56553 , n56554 );
and ( n56556 , n55350 , n55351 );
and ( n56557 , n55352 , n55355 );
or ( n56558 , n56556 , n56557 );
xor ( n56559 , n56555 , n56558 );
nor ( n56560 , n30716 , n1768 );
xor ( n56561 , n56559 , n56560 );
and ( n56562 , n55356 , n55357 );
and ( n56563 , n55358 , n55361 );
or ( n56564 , n56562 , n56563 );
xor ( n56565 , n56561 , n56564 );
nor ( n56566 , n31858 , n1947 );
xor ( n56567 , n56565 , n56566 );
and ( n56568 , n55362 , n55363 );
and ( n56569 , n55364 , n55367 );
or ( n56570 , n56568 , n56569 );
xor ( n56571 , n56567 , n56570 );
nor ( n56572 , n33024 , n2139 );
xor ( n56573 , n56571 , n56572 );
and ( n56574 , n55368 , n55369 );
and ( n56575 , n55370 , n55373 );
or ( n56576 , n56574 , n56575 );
xor ( n56577 , n56573 , n56576 );
nor ( n56578 , n34215 , n2345 );
xor ( n56579 , n56577 , n56578 );
and ( n56580 , n55374 , n55375 );
and ( n56581 , n55376 , n55379 );
or ( n56582 , n56580 , n56581 );
xor ( n56583 , n56579 , n56582 );
nor ( n56584 , n35410 , n2568 );
xor ( n56585 , n56583 , n56584 );
and ( n56586 , n55380 , n55381 );
and ( n56587 , n55382 , n55385 );
or ( n56588 , n56586 , n56587 );
xor ( n56589 , n56585 , n56588 );
nor ( n56590 , n36611 , n2799 );
xor ( n56591 , n56589 , n56590 );
and ( n56592 , n55386 , n55387 );
and ( n56593 , n55388 , n55391 );
or ( n56594 , n56592 , n56593 );
xor ( n56595 , n56591 , n56594 );
nor ( n56596 , n37816 , n3045 );
xor ( n56597 , n56595 , n56596 );
and ( n56598 , n55392 , n55393 );
and ( n56599 , n55394 , n55397 );
or ( n56600 , n56598 , n56599 );
xor ( n56601 , n56597 , n56600 );
nor ( n56602 , n39018 , n3302 );
xor ( n56603 , n56601 , n56602 );
and ( n56604 , n55398 , n55399 );
and ( n56605 , n55400 , n55403 );
or ( n56606 , n56604 , n56605 );
xor ( n56607 , n56603 , n56606 );
nor ( n56608 , n40223 , n3572 );
xor ( n56609 , n56607 , n56608 );
and ( n56610 , n55404 , n55405 );
and ( n56611 , n55406 , n55409 );
or ( n56612 , n56610 , n56611 );
xor ( n56613 , n56609 , n56612 );
nor ( n56614 , n41428 , n3855 );
xor ( n56615 , n56613 , n56614 );
and ( n56616 , n55410 , n55411 );
and ( n56617 , n55412 , n55415 );
or ( n56618 , n56616 , n56617 );
xor ( n56619 , n56615 , n56618 );
nor ( n56620 , n42632 , n4153 );
xor ( n56621 , n56619 , n56620 );
and ( n56622 , n55416 , n55417 );
and ( n56623 , n55418 , n55421 );
or ( n56624 , n56622 , n56623 );
xor ( n56625 , n56621 , n56624 );
nor ( n56626 , n43834 , n4460 );
xor ( n56627 , n56625 , n56626 );
and ( n56628 , n55422 , n55423 );
and ( n56629 , n55424 , n55427 );
or ( n56630 , n56628 , n56629 );
xor ( n56631 , n56627 , n56630 );
nor ( n56632 , n45038 , n4788 );
xor ( n56633 , n56631 , n56632 );
and ( n56634 , n55428 , n55429 );
and ( n56635 , n55430 , n55433 );
or ( n56636 , n56634 , n56635 );
xor ( n56637 , n56633 , n56636 );
nor ( n56638 , n46239 , n5128 );
xor ( n56639 , n56637 , n56638 );
and ( n56640 , n55434 , n55435 );
and ( n56641 , n55436 , n55439 );
or ( n56642 , n56640 , n56641 );
xor ( n56643 , n56639 , n56642 );
nor ( n56644 , n47440 , n5479 );
xor ( n56645 , n56643 , n56644 );
and ( n56646 , n55440 , n55441 );
and ( n56647 , n55442 , n55445 );
or ( n56648 , n56646 , n56647 );
xor ( n56649 , n56645 , n56648 );
nor ( n56650 , n48641 , n5840 );
xor ( n56651 , n56649 , n56650 );
and ( n56652 , n55446 , n55447 );
and ( n56653 , n55448 , n55451 );
or ( n56654 , n56652 , n56653 );
xor ( n56655 , n56651 , n56654 );
nor ( n56656 , n49841 , n6214 );
xor ( n56657 , n56655 , n56656 );
and ( n56658 , n55452 , n55453 );
and ( n56659 , n55454 , n55457 );
or ( n56660 , n56658 , n56659 );
xor ( n56661 , n56657 , n56660 );
nor ( n56662 , n51040 , n6598 );
xor ( n56663 , n56661 , n56662 );
and ( n56664 , n55458 , n55459 );
and ( n56665 , n55460 , n55463 );
or ( n56666 , n56664 , n56665 );
xor ( n56667 , n56663 , n56666 );
nor ( n56668 , n52238 , n6999 );
xor ( n56669 , n56667 , n56668 );
and ( n56670 , n55464 , n55465 );
and ( n56671 , n55466 , n55469 );
or ( n56672 , n56670 , n56671 );
xor ( n56673 , n56669 , n56672 );
nor ( n56674 , n53432 , n7415 );
xor ( n56675 , n56673 , n56674 );
and ( n56676 , n55470 , n55471 );
and ( n56677 , n55472 , n55475 );
or ( n56678 , n56676 , n56677 );
xor ( n56679 , n56675 , n56678 );
nor ( n56680 , n54629 , n7843 );
xor ( n56681 , n56679 , n56680 );
and ( n56682 , n55476 , n55477 );
and ( n56683 , n55478 , n55481 );
or ( n56684 , n56682 , n56683 );
xor ( n56685 , n56681 , n56684 );
nor ( n56686 , n55826 , n8283 );
xor ( n56687 , n56685 , n56686 );
and ( n56688 , n55482 , n55483 );
and ( n56689 , n55484 , n55487 );
or ( n56690 , n56688 , n56689 );
xor ( n56691 , n56687 , n56690 );
and ( n56692 , n55500 , n55504 );
and ( n56693 , n55504 , n55812 );
and ( n56694 , n55500 , n55812 );
or ( n56695 , n56692 , n56693 , n56694 );
and ( n56696 , n33774 , n2739 );
not ( n56697 , n2739 );
nor ( n56698 , n56696 , n56697 );
xor ( n56699 , n56695 , n56698 );
and ( n56700 , n55513 , n55517 );
and ( n56701 , n55517 , n55585 );
and ( n56702 , n55513 , n55585 );
or ( n56703 , n56700 , n56701 , n56702 );
and ( n56704 , n55509 , n55586 );
and ( n56705 , n55586 , n55811 );
and ( n56706 , n55509 , n55811 );
or ( n56707 , n56704 , n56705 , n56706 );
xor ( n56708 , n56703 , n56707 );
and ( n56709 , n55588 , n55708 );
and ( n56710 , n55708 , n55810 );
and ( n56711 , n55588 , n55810 );
or ( n56712 , n56709 , n56710 , n56711 );
and ( n56713 , n55522 , n55526 );
and ( n56714 , n55526 , n55584 );
and ( n56715 , n55522 , n55584 );
or ( n56716 , n56713 , n56714 , n56715 );
and ( n56717 , n55592 , n55596 );
and ( n56718 , n55596 , n55707 );
and ( n56719 , n55592 , n55707 );
or ( n56720 , n56717 , n56718 , n56719 );
xor ( n56721 , n56716 , n56720 );
and ( n56722 , n55553 , n55557 );
and ( n56723 , n55557 , n55563 );
and ( n56724 , n55553 , n55563 );
or ( n56725 , n56722 , n56723 , n56724 );
and ( n56726 , n55531 , n55535 );
and ( n56727 , n55535 , n55583 );
and ( n56728 , n55531 , n55583 );
or ( n56729 , n56726 , n56727 , n56728 );
xor ( n56730 , n56725 , n56729 );
and ( n56731 , n55540 , n55544 );
and ( n56732 , n55544 , n55582 );
and ( n56733 , n55540 , n55582 );
or ( n56734 , n56731 , n56732 , n56733 );
and ( n56735 , n55605 , n55630 );
and ( n56736 , n55630 , n55668 );
and ( n56737 , n55605 , n55668 );
or ( n56738 , n56735 , n56736 , n56737 );
xor ( n56739 , n56734 , n56738 );
and ( n56740 , n55549 , n55564 );
and ( n56741 , n55564 , n55581 );
and ( n56742 , n55549 , n55581 );
or ( n56743 , n56740 , n56741 , n56742 );
and ( n56744 , n55609 , n55613 );
and ( n56745 , n55613 , n55629 );
and ( n56746 , n55609 , n55629 );
or ( n56747 , n56744 , n56745 , n56746 );
xor ( n56748 , n56743 , n56747 );
and ( n56749 , n55569 , n55574 );
and ( n56750 , n55574 , n55580 );
and ( n56751 , n55569 , n55580 );
or ( n56752 , n56749 , n56750 , n56751 );
and ( n56753 , n55559 , n55560 );
and ( n56754 , n55560 , n55562 );
and ( n56755 , n55559 , n55562 );
or ( n56756 , n56753 , n56754 , n56755 );
and ( n56757 , n55570 , n55571 );
and ( n56758 , n55571 , n55573 );
and ( n56759 , n55570 , n55573 );
or ( n56760 , n56757 , n56758 , n56759 );
xor ( n56761 , n56756 , n56760 );
and ( n56762 , n30695 , n3495 );
and ( n56763 , n31836 , n3271 );
xor ( n56764 , n56762 , n56763 );
and ( n56765 , n32649 , n2981 );
xor ( n56766 , n56764 , n56765 );
xor ( n56767 , n56761 , n56766 );
xor ( n56768 , n56752 , n56767 );
and ( n56769 , n55576 , n55577 );
and ( n56770 , n55577 , n55579 );
and ( n56771 , n55576 , n55579 );
or ( n56772 , n56769 , n56770 , n56771 );
and ( n56773 , n27361 , n4403 );
and ( n56774 , n28456 , n4102 );
xor ( n56775 , n56773 , n56774 );
and ( n56776 , n29559 , n3749 );
xor ( n56777 , n56775 , n56776 );
xor ( n56778 , n56772 , n56777 );
and ( n56779 , n24214 , n5408 );
and ( n56780 , n25243 , n5103 );
xor ( n56781 , n56779 , n56780 );
and ( n56782 , n26296 , n4730 );
xor ( n56783 , n56781 , n56782 );
xor ( n56784 , n56778 , n56783 );
xor ( n56785 , n56768 , n56784 );
xor ( n56786 , n56748 , n56785 );
xor ( n56787 , n56739 , n56786 );
xor ( n56788 , n56730 , n56787 );
xor ( n56789 , n56721 , n56788 );
xor ( n56790 , n56712 , n56789 );
and ( n56791 , n55784 , n55809 );
and ( n56792 , n55713 , n55714 );
and ( n56793 , n55714 , n55783 );
and ( n56794 , n55713 , n55783 );
or ( n56795 , n56792 , n56793 , n56794 );
and ( n56796 , n55601 , n55669 );
and ( n56797 , n55669 , n55706 );
and ( n56798 , n55601 , n55706 );
or ( n56799 , n56796 , n56797 , n56798 );
xor ( n56800 , n56795 , n56799 );
and ( n56801 , n55674 , n55678 );
and ( n56802 , n55678 , n55705 );
and ( n56803 , n55674 , n55705 );
or ( n56804 , n56801 , n56802 , n56803 );
and ( n56805 , n55635 , n55651 );
and ( n56806 , n55651 , n55667 );
and ( n56807 , n55635 , n55667 );
or ( n56808 , n56805 , n56806 , n56807 );
and ( n56809 , n55618 , n55622 );
and ( n56810 , n55622 , n55628 );
and ( n56811 , n55618 , n55628 );
or ( n56812 , n56809 , n56810 , n56811 );
and ( n56813 , n55639 , n55644 );
and ( n56814 , n55644 , n55650 );
and ( n56815 , n55639 , n55650 );
or ( n56816 , n56813 , n56814 , n56815 );
xor ( n56817 , n56812 , n56816 );
and ( n56818 , n55624 , n55625 );
and ( n56819 , n55625 , n55627 );
and ( n56820 , n55624 , n55627 );
or ( n56821 , n56818 , n56819 , n56820 );
and ( n56822 , n55640 , n55641 );
and ( n56823 , n55641 , n55643 );
and ( n56824 , n55640 , n55643 );
or ( n56825 , n56822 , n56823 , n56824 );
xor ( n56826 , n56821 , n56825 );
and ( n56827 , n21216 , n6504 );
and ( n56828 , n22186 , n6132 );
xor ( n56829 , n56827 , n56828 );
and ( n56830 , n22892 , n5765 );
xor ( n56831 , n56829 , n56830 );
xor ( n56832 , n56826 , n56831 );
xor ( n56833 , n56817 , n56832 );
xor ( n56834 , n56808 , n56833 );
and ( n56835 , n55656 , n55660 );
and ( n56836 , n55660 , n55666 );
and ( n56837 , n55656 , n55666 );
or ( n56838 , n56835 , n56836 , n56837 );
and ( n56839 , n55646 , n55647 );
and ( n56840 , n55647 , n55649 );
and ( n56841 , n55646 , n55649 );
or ( n56842 , n56839 , n56840 , n56841 );
and ( n56843 , n18144 , n7662 );
and ( n56844 , n19324 , n7310 );
xor ( n56845 , n56843 , n56844 );
and ( n56846 , n20233 , n6971 );
xor ( n56847 , n56845 , n56846 );
xor ( n56848 , n56842 , n56847 );
and ( n56849 , n15758 , n9348 );
and ( n56850 , n16637 , n8669 );
xor ( n56851 , n56849 , n56850 );
and ( n56852 , n17512 , n8243 );
xor ( n56853 , n56851 , n56852 );
xor ( n56854 , n56848 , n56853 );
xor ( n56855 , n56838 , n56854 );
and ( n56856 , n55662 , n55663 );
and ( n56857 , n55663 , n55665 );
and ( n56858 , n55662 , n55665 );
or ( n56859 , n56856 , n56857 , n56858 );
and ( n56860 , n55693 , n55694 );
and ( n56861 , n55694 , n55696 );
and ( n56862 , n55693 , n55696 );
or ( n56863 , n56860 , n56861 , n56862 );
xor ( n56864 , n56859 , n56863 );
and ( n56865 , n13322 , n11718 );
and ( n56866 , n14118 , n10977 );
xor ( n56867 , n56865 , n56866 );
and ( n56868 , n14938 , n10239 );
xor ( n56869 , n56867 , n56868 );
xor ( n56870 , n56864 , n56869 );
xor ( n56871 , n56855 , n56870 );
xor ( n56872 , n56834 , n56871 );
xor ( n56873 , n56804 , n56872 );
and ( n56874 , n55683 , n55687 );
and ( n56875 , n55687 , n55704 );
and ( n56876 , n55683 , n55704 );
or ( n56877 , n56874 , n56875 , n56876 );
and ( n56878 , n55749 , n55764 );
and ( n56879 , n55764 , n55781 );
and ( n56880 , n55749 , n55781 );
or ( n56881 , n56878 , n56879 , n56880 );
xor ( n56882 , n56877 , n56881 );
and ( n56883 , n55692 , n55697 );
and ( n56884 , n55697 , n55703 );
and ( n56885 , n55692 , n55703 );
or ( n56886 , n56883 , n56884 , n56885 );
and ( n56887 , n55753 , n55757 );
and ( n56888 , n55757 , n55763 );
and ( n56889 , n55753 , n55763 );
or ( n56890 , n56887 , n56888 , n56889 );
xor ( n56891 , n56886 , n56890 );
and ( n56892 , n55699 , n55700 );
and ( n56893 , n55700 , n55702 );
and ( n56894 , n55699 , n55702 );
or ( n56895 , n56892 , n56893 , n56894 );
and ( n56896 , n11015 , n14044 );
and ( n56897 , n11769 , n13256 );
xor ( n56898 , n56896 , n56897 );
buf ( n56899 , n12320 );
xor ( n56900 , n56898 , n56899 );
xor ( n56901 , n56895 , n56900 );
and ( n56902 , n8718 , n16550 );
and ( n56903 , n9400 , n15691 );
xor ( n56904 , n56902 , n56903 );
and ( n56905 , n10291 , n14838 );
xor ( n56906 , n56904 , n56905 );
xor ( n56907 , n56901 , n56906 );
xor ( n56908 , n56891 , n56907 );
xor ( n56909 , n56882 , n56908 );
xor ( n56910 , n56873 , n56909 );
xor ( n56911 , n56800 , n56910 );
xor ( n56912 , n56791 , n56911 );
and ( n56913 , n55719 , n55744 );
and ( n56914 , n55744 , n55782 );
and ( n56915 , n55719 , n55782 );
or ( n56916 , n56913 , n56914 , n56915 );
and ( n56917 , n55788 , n55808 );
xor ( n56918 , n56916 , n56917 );
and ( n56919 , n55723 , n55727 );
and ( n56920 , n55727 , n55743 );
and ( n56921 , n55723 , n55743 );
or ( n56922 , n56919 , n56920 , n56921 );
and ( n56923 , n55769 , n55774 );
and ( n56924 , n55774 , n55780 );
and ( n56925 , n55769 , n55780 );
or ( n56926 , n56923 , n56924 , n56925 );
and ( n56927 , n55759 , n55760 );
and ( n56928 , n55760 , n55762 );
and ( n56929 , n55759 , n55762 );
or ( n56930 , n56927 , n56928 , n56929 );
and ( n56931 , n55770 , n55771 );
and ( n56932 , n55771 , n55773 );
and ( n56933 , n55770 , n55773 );
or ( n56934 , n56931 , n56932 , n56933 );
xor ( n56935 , n56930 , n56934 );
and ( n56936 , n7385 , n19222 );
and ( n56937 , n7808 , n18407 );
xor ( n56938 , n56936 , n56937 );
and ( n56939 , n8079 , n17422 );
xor ( n56940 , n56938 , n56939 );
xor ( n56941 , n56935 , n56940 );
xor ( n56942 , n56926 , n56941 );
and ( n56943 , n55776 , n55777 );
and ( n56944 , n55777 , n55779 );
and ( n56945 , n55776 , n55779 );
or ( n56946 , n56943 , n56944 , n56945 );
and ( n56947 , n6187 , n22065 );
and ( n56948 , n6569 , n20976 );
xor ( n56949 , n56947 , n56948 );
and ( n56950 , n6816 , n20156 );
xor ( n56951 , n56949 , n56950 );
xor ( n56952 , n56946 , n56951 );
and ( n56953 , n4959 , n25163 );
and ( n56954 , n5459 , n24137 );
xor ( n56955 , n56953 , n56954 );
and ( n56956 , n5819 , n23075 );
xor ( n56957 , n56955 , n56956 );
xor ( n56958 , n56952 , n56957 );
xor ( n56959 , n56942 , n56958 );
xor ( n56960 , n56922 , n56959 );
and ( n56961 , n55793 , n55798 );
and ( n56962 , n55798 , n55806 );
and ( n56963 , n55793 , n55806 );
or ( n56964 , n56961 , n56962 , n56963 );
and ( n56965 , n55732 , n55736 );
and ( n56966 , n55736 , n55742 );
and ( n56967 , n55732 , n55742 );
or ( n56968 , n56965 , n56966 , n56967 );
xor ( n56969 , n56964 , n56968 );
and ( n56970 , n55738 , n55739 );
and ( n56971 , n55739 , n55741 );
and ( n56972 , n55738 , n55741 );
or ( n56973 , n56970 , n56971 , n56972 );
and ( n56974 , n55794 , n55795 );
and ( n56975 , n55795 , n55797 );
and ( n56976 , n55794 , n55797 );
or ( n56977 , n56974 , n56975 , n56976 );
xor ( n56978 , n56973 , n56977 );
and ( n56979 , n4132 , n28406 );
and ( n56980 , n4438 , n27296 );
xor ( n56981 , n56979 , n56980 );
and ( n56982 , n4766 , n26216 );
xor ( n56983 , n56981 , n56982 );
xor ( n56984 , n56978 , n56983 );
xor ( n56985 , n56969 , n56984 );
xor ( n56986 , n56960 , n56985 );
xor ( n56987 , n56918 , n56986 );
and ( n56988 , n55789 , n55807 );
and ( n56989 , n55802 , n55803 );
and ( n56990 , n55803 , n55805 );
and ( n56991 , n55802 , n55805 );
or ( n56992 , n56989 , n56990 , n56991 );
and ( n56993 , n3182 , n31761 );
and ( n56994 , n3545 , n30629 );
xor ( n56995 , n56993 , n56994 );
and ( n56996 , n3801 , n29508 );
xor ( n56997 , n56995 , n56996 );
xor ( n56998 , n56992 , n56997 );
not ( n56999 , n2779 );
and ( n57000 , n34193 , n2779 );
nor ( n57001 , n56999 , n57000 );
and ( n57002 , n3024 , n32999 );
xor ( n57003 , n57001 , n57002 );
xor ( n57004 , n56998 , n57003 );
xor ( n57005 , n56988 , n57004 );
xor ( n57006 , n56987 , n57005 );
xor ( n57007 , n56912 , n57006 );
xor ( n57008 , n56790 , n57007 );
xor ( n57009 , n56708 , n57008 );
xor ( n57010 , n56699 , n57009 );
and ( n57011 , n55492 , n55495 );
and ( n57012 , n55495 , n55813 );
and ( n57013 , n55492 , n55813 );
or ( n57014 , n57011 , n57012 , n57013 );
xor ( n57015 , n57010 , n57014 );
and ( n57016 , n55814 , n55818 );
and ( n57017 , n55819 , n55822 );
or ( n57018 , n57016 , n57017 );
xor ( n57019 , n57015 , n57018 );
buf ( n57020 , n57019 );
buf ( n57021 , n57020 );
not ( n57022 , n57021 );
nor ( n57023 , n57022 , n8739 );
xor ( n57024 , n56691 , n57023 );
and ( n57025 , n55488 , n55827 );
and ( n57026 , n55828 , n55831 );
or ( n57027 , n57025 , n57026 );
xor ( n57028 , n57024 , n57027 );
buf ( n57029 , n57028 );
buf ( n57030 , n57029 );
not ( n57031 , n57030 );
buf ( n57032 , n581 );
not ( n57033 , n57032 );
nor ( n57034 , n57031 , n57033 );
xor ( n57035 , n56317 , n57034 );
xor ( n57036 , n55843 , n56314 );
nor ( n57037 , n55835 , n57033 );
and ( n57038 , n57036 , n57037 );
xor ( n57039 , n57036 , n57037 );
xor ( n57040 , n55847 , n56312 );
nor ( n57041 , n54638 , n57033 );
and ( n57042 , n57040 , n57041 );
xor ( n57043 , n57040 , n57041 );
xor ( n57044 , n55851 , n56310 );
nor ( n57045 , n53441 , n57033 );
and ( n57046 , n57044 , n57045 );
xor ( n57047 , n57044 , n57045 );
xor ( n57048 , n55855 , n56308 );
nor ( n57049 , n52247 , n57033 );
and ( n57050 , n57048 , n57049 );
xor ( n57051 , n57048 , n57049 );
xor ( n57052 , n55859 , n56306 );
nor ( n57053 , n51049 , n57033 );
and ( n57054 , n57052 , n57053 );
xor ( n57055 , n57052 , n57053 );
xor ( n57056 , n55863 , n56304 );
nor ( n57057 , n49850 , n57033 );
and ( n57058 , n57056 , n57057 );
xor ( n57059 , n57056 , n57057 );
xor ( n57060 , n55867 , n56302 );
nor ( n57061 , n48650 , n57033 );
and ( n57062 , n57060 , n57061 );
xor ( n57063 , n57060 , n57061 );
xor ( n57064 , n55871 , n56300 );
nor ( n57065 , n47449 , n57033 );
and ( n57066 , n57064 , n57065 );
xor ( n57067 , n57064 , n57065 );
xor ( n57068 , n55875 , n56298 );
nor ( n57069 , n46248 , n57033 );
and ( n57070 , n57068 , n57069 );
xor ( n57071 , n57068 , n57069 );
xor ( n57072 , n55879 , n56296 );
nor ( n57073 , n45047 , n57033 );
and ( n57074 , n57072 , n57073 );
xor ( n57075 , n57072 , n57073 );
xor ( n57076 , n55883 , n56294 );
nor ( n57077 , n43843 , n57033 );
and ( n57078 , n57076 , n57077 );
xor ( n57079 , n57076 , n57077 );
xor ( n57080 , n55887 , n56292 );
nor ( n57081 , n42641 , n57033 );
and ( n57082 , n57080 , n57081 );
xor ( n57083 , n57080 , n57081 );
xor ( n57084 , n55891 , n56290 );
nor ( n57085 , n41437 , n57033 );
and ( n57086 , n57084 , n57085 );
xor ( n57087 , n57084 , n57085 );
xor ( n57088 , n55895 , n56288 );
nor ( n57089 , n40232 , n57033 );
and ( n57090 , n57088 , n57089 );
xor ( n57091 , n57088 , n57089 );
xor ( n57092 , n55899 , n56286 );
nor ( n57093 , n39027 , n57033 );
and ( n57094 , n57092 , n57093 );
xor ( n57095 , n57092 , n57093 );
xor ( n57096 , n55903 , n56284 );
nor ( n57097 , n37825 , n57033 );
and ( n57098 , n57096 , n57097 );
xor ( n57099 , n57096 , n57097 );
xor ( n57100 , n55907 , n56282 );
nor ( n57101 , n36620 , n57033 );
and ( n57102 , n57100 , n57101 );
xor ( n57103 , n57100 , n57101 );
xor ( n57104 , n55911 , n56280 );
nor ( n57105 , n35419 , n57033 );
and ( n57106 , n57104 , n57105 );
xor ( n57107 , n57104 , n57105 );
xor ( n57108 , n55915 , n56278 );
nor ( n57109 , n34224 , n57033 );
and ( n57110 , n57108 , n57109 );
xor ( n57111 , n57108 , n57109 );
xor ( n57112 , n55919 , n56276 );
nor ( n57113 , n33033 , n57033 );
and ( n57114 , n57112 , n57113 );
xor ( n57115 , n57112 , n57113 );
xor ( n57116 , n55923 , n56274 );
nor ( n57117 , n31867 , n57033 );
and ( n57118 , n57116 , n57117 );
xor ( n57119 , n57116 , n57117 );
xor ( n57120 , n55927 , n56272 );
nor ( n57121 , n30725 , n57033 );
and ( n57122 , n57120 , n57121 );
xor ( n57123 , n57120 , n57121 );
xor ( n57124 , n55931 , n56270 );
nor ( n57125 , n29596 , n57033 );
and ( n57126 , n57124 , n57125 );
xor ( n57127 , n57124 , n57125 );
xor ( n57128 , n55935 , n56268 );
nor ( n57129 , n28487 , n57033 );
and ( n57130 , n57128 , n57129 );
xor ( n57131 , n57128 , n57129 );
xor ( n57132 , n55939 , n56266 );
nor ( n57133 , n27397 , n57033 );
and ( n57134 , n57132 , n57133 );
xor ( n57135 , n57132 , n57133 );
xor ( n57136 , n55943 , n56264 );
nor ( n57137 , n26326 , n57033 );
and ( n57138 , n57136 , n57137 );
xor ( n57139 , n57136 , n57137 );
xor ( n57140 , n55947 , n56262 );
nor ( n57141 , n25272 , n57033 );
and ( n57142 , n57140 , n57141 );
xor ( n57143 , n57140 , n57141 );
xor ( n57144 , n55951 , n56260 );
nor ( n57145 , n24242 , n57033 );
and ( n57146 , n57144 , n57145 );
xor ( n57147 , n57144 , n57145 );
xor ( n57148 , n55955 , n56258 );
nor ( n57149 , n23225 , n57033 );
and ( n57150 , n57148 , n57149 );
xor ( n57151 , n57148 , n57149 );
xor ( n57152 , n55959 , n56256 );
nor ( n57153 , n22231 , n57033 );
and ( n57154 , n57152 , n57153 );
xor ( n57155 , n57152 , n57153 );
xor ( n57156 , n55963 , n56254 );
nor ( n57157 , n21258 , n57033 );
and ( n57158 , n57156 , n57157 );
xor ( n57159 , n57156 , n57157 );
xor ( n57160 , n55967 , n56252 );
nor ( n57161 , n20303 , n57033 );
and ( n57162 , n57160 , n57161 );
xor ( n57163 , n57160 , n57161 );
xor ( n57164 , n55971 , n56250 );
nor ( n57165 , n19365 , n57033 );
and ( n57166 , n57164 , n57165 );
xor ( n57167 , n57164 , n57165 );
xor ( n57168 , n55975 , n56248 );
nor ( n57169 , n18448 , n57033 );
and ( n57170 , n57168 , n57169 );
xor ( n57171 , n57168 , n57169 );
xor ( n57172 , n55979 , n56246 );
nor ( n57173 , n17548 , n57033 );
and ( n57174 , n57172 , n57173 );
xor ( n57175 , n57172 , n57173 );
xor ( n57176 , n55983 , n56244 );
nor ( n57177 , n16669 , n57033 );
and ( n57178 , n57176 , n57177 );
xor ( n57179 , n57176 , n57177 );
xor ( n57180 , n55987 , n56242 );
nor ( n57181 , n15809 , n57033 );
and ( n57182 , n57180 , n57181 );
xor ( n57183 , n57180 , n57181 );
xor ( n57184 , n55991 , n56240 );
nor ( n57185 , n14968 , n57033 );
and ( n57186 , n57184 , n57185 );
xor ( n57187 , n57184 , n57185 );
xor ( n57188 , n55995 , n56238 );
nor ( n57189 , n14147 , n57033 );
and ( n57190 , n57188 , n57189 );
xor ( n57191 , n57188 , n57189 );
xor ( n57192 , n55999 , n56236 );
nor ( n57193 , n13349 , n57033 );
and ( n57194 , n57192 , n57193 );
xor ( n57195 , n57192 , n57193 );
xor ( n57196 , n56003 , n56234 );
nor ( n57197 , n12564 , n57033 );
and ( n57198 , n57196 , n57197 );
xor ( n57199 , n57196 , n57197 );
xor ( n57200 , n56007 , n56232 );
nor ( n57201 , n11799 , n57033 );
and ( n57202 , n57200 , n57201 );
xor ( n57203 , n57200 , n57201 );
xor ( n57204 , n56011 , n56230 );
nor ( n57205 , n11050 , n57033 );
and ( n57206 , n57204 , n57205 );
xor ( n57207 , n57204 , n57205 );
xor ( n57208 , n56015 , n56228 );
nor ( n57209 , n10321 , n57033 );
and ( n57210 , n57208 , n57209 );
xor ( n57211 , n57208 , n57209 );
xor ( n57212 , n56019 , n56226 );
nor ( n57213 , n9429 , n57033 );
and ( n57214 , n57212 , n57213 );
xor ( n57215 , n57212 , n57213 );
xor ( n57216 , n56023 , n56224 );
nor ( n57217 , n8949 , n57033 );
and ( n57218 , n57216 , n57217 );
xor ( n57219 , n57216 , n57217 );
xor ( n57220 , n56027 , n56222 );
nor ( n57221 , n9437 , n57033 );
and ( n57222 , n57220 , n57221 );
xor ( n57223 , n57220 , n57221 );
xor ( n57224 , n56031 , n56220 );
nor ( n57225 , n9446 , n57033 );
and ( n57226 , n57224 , n57225 );
xor ( n57227 , n57224 , n57225 );
xor ( n57228 , n56035 , n56218 );
nor ( n57229 , n9455 , n57033 );
and ( n57230 , n57228 , n57229 );
xor ( n57231 , n57228 , n57229 );
xor ( n57232 , n56039 , n56216 );
nor ( n57233 , n9464 , n57033 );
and ( n57234 , n57232 , n57233 );
xor ( n57235 , n57232 , n57233 );
xor ( n57236 , n56043 , n56214 );
nor ( n57237 , n9473 , n57033 );
and ( n57238 , n57236 , n57237 );
xor ( n57239 , n57236 , n57237 );
xor ( n57240 , n56047 , n56212 );
nor ( n57241 , n9482 , n57033 );
and ( n57242 , n57240 , n57241 );
xor ( n57243 , n57240 , n57241 );
xor ( n57244 , n56051 , n56210 );
nor ( n57245 , n9491 , n57033 );
and ( n57246 , n57244 , n57245 );
xor ( n57247 , n57244 , n57245 );
xor ( n57248 , n56055 , n56208 );
nor ( n57249 , n9500 , n57033 );
and ( n57250 , n57248 , n57249 );
xor ( n57251 , n57248 , n57249 );
xor ( n57252 , n56059 , n56206 );
nor ( n57253 , n9509 , n57033 );
and ( n57254 , n57252 , n57253 );
xor ( n57255 , n57252 , n57253 );
xor ( n57256 , n56063 , n56204 );
nor ( n57257 , n9518 , n57033 );
and ( n57258 , n57256 , n57257 );
xor ( n57259 , n57256 , n57257 );
xor ( n57260 , n56067 , n56202 );
nor ( n57261 , n9527 , n57033 );
and ( n57262 , n57260 , n57261 );
xor ( n57263 , n57260 , n57261 );
xor ( n57264 , n56071 , n56200 );
nor ( n57265 , n9536 , n57033 );
and ( n57266 , n57264 , n57265 );
xor ( n57267 , n57264 , n57265 );
xor ( n57268 , n56075 , n56198 );
nor ( n57269 , n9545 , n57033 );
and ( n57270 , n57268 , n57269 );
xor ( n57271 , n57268 , n57269 );
xor ( n57272 , n56079 , n56196 );
nor ( n57273 , n9554 , n57033 );
and ( n57274 , n57272 , n57273 );
xor ( n57275 , n57272 , n57273 );
xor ( n57276 , n56083 , n56194 );
nor ( n57277 , n9563 , n57033 );
and ( n57278 , n57276 , n57277 );
xor ( n57279 , n57276 , n57277 );
xor ( n57280 , n56087 , n56192 );
nor ( n57281 , n9572 , n57033 );
and ( n57282 , n57280 , n57281 );
xor ( n57283 , n57280 , n57281 );
xor ( n57284 , n56091 , n56190 );
nor ( n57285 , n9581 , n57033 );
and ( n57286 , n57284 , n57285 );
xor ( n57287 , n57284 , n57285 );
xor ( n57288 , n56095 , n56188 );
nor ( n57289 , n9590 , n57033 );
and ( n57290 , n57288 , n57289 );
xor ( n57291 , n57288 , n57289 );
xor ( n57292 , n56099 , n56186 );
nor ( n57293 , n9599 , n57033 );
and ( n57294 , n57292 , n57293 );
xor ( n57295 , n57292 , n57293 );
xor ( n57296 , n56103 , n56184 );
nor ( n57297 , n9608 , n57033 );
and ( n57298 , n57296 , n57297 );
xor ( n57299 , n57296 , n57297 );
xor ( n57300 , n56107 , n56182 );
nor ( n57301 , n9617 , n57033 );
and ( n57302 , n57300 , n57301 );
xor ( n57303 , n57300 , n57301 );
xor ( n57304 , n56111 , n56180 );
nor ( n57305 , n9626 , n57033 );
and ( n57306 , n57304 , n57305 );
xor ( n57307 , n57304 , n57305 );
xor ( n57308 , n56115 , n56178 );
nor ( n57309 , n9635 , n57033 );
and ( n57310 , n57308 , n57309 );
xor ( n57311 , n57308 , n57309 );
xor ( n57312 , n56119 , n56176 );
nor ( n57313 , n9644 , n57033 );
and ( n57314 , n57312 , n57313 );
xor ( n57315 , n57312 , n57313 );
xor ( n57316 , n56123 , n56174 );
nor ( n57317 , n9653 , n57033 );
and ( n57318 , n57316 , n57317 );
xor ( n57319 , n57316 , n57317 );
xor ( n57320 , n56127 , n56172 );
nor ( n57321 , n9662 , n57033 );
and ( n57322 , n57320 , n57321 );
xor ( n57323 , n57320 , n57321 );
xor ( n57324 , n56131 , n56170 );
nor ( n57325 , n9671 , n57033 );
and ( n57326 , n57324 , n57325 );
xor ( n57327 , n57324 , n57325 );
xor ( n57328 , n56135 , n56168 );
nor ( n57329 , n9680 , n57033 );
and ( n57330 , n57328 , n57329 );
xor ( n57331 , n57328 , n57329 );
xor ( n57332 , n56139 , n56166 );
nor ( n57333 , n9689 , n57033 );
and ( n57334 , n57332 , n57333 );
xor ( n57335 , n57332 , n57333 );
xor ( n57336 , n56143 , n56164 );
nor ( n57337 , n9698 , n57033 );
and ( n57338 , n57336 , n57337 );
xor ( n57339 , n57336 , n57337 );
xor ( n57340 , n56147 , n56162 );
nor ( n57341 , n9707 , n57033 );
and ( n57342 , n57340 , n57341 );
xor ( n57343 , n57340 , n57341 );
xor ( n57344 , n56151 , n56160 );
nor ( n57345 , n9716 , n57033 );
and ( n57346 , n57344 , n57345 );
xor ( n57347 , n57344 , n57345 );
xor ( n57348 , n56155 , n56158 );
nor ( n57349 , n9725 , n57033 );
and ( n57350 , n57348 , n57349 );
xor ( n57351 , n57348 , n57349 );
xor ( n57352 , n56156 , n56157 );
nor ( n57353 , n9734 , n57033 );
and ( n57354 , n57352 , n57353 );
xor ( n57355 , n57352 , n57353 );
nor ( n57356 , n9752 , n55837 );
nor ( n57357 , n9743 , n57033 );
and ( n57358 , n57356 , n57357 );
and ( n57359 , n57355 , n57358 );
or ( n57360 , n57354 , n57359 );
and ( n57361 , n57351 , n57360 );
or ( n57362 , n57350 , n57361 );
and ( n57363 , n57347 , n57362 );
or ( n57364 , n57346 , n57363 );
and ( n57365 , n57343 , n57364 );
or ( n57366 , n57342 , n57365 );
and ( n57367 , n57339 , n57366 );
or ( n57368 , n57338 , n57367 );
and ( n57369 , n57335 , n57368 );
or ( n57370 , n57334 , n57369 );
and ( n57371 , n57331 , n57370 );
or ( n57372 , n57330 , n57371 );
and ( n57373 , n57327 , n57372 );
or ( n57374 , n57326 , n57373 );
and ( n57375 , n57323 , n57374 );
or ( n57376 , n57322 , n57375 );
and ( n57377 , n57319 , n57376 );
or ( n57378 , n57318 , n57377 );
and ( n57379 , n57315 , n57378 );
or ( n57380 , n57314 , n57379 );
and ( n57381 , n57311 , n57380 );
or ( n57382 , n57310 , n57381 );
and ( n57383 , n57307 , n57382 );
or ( n57384 , n57306 , n57383 );
and ( n57385 , n57303 , n57384 );
or ( n57386 , n57302 , n57385 );
and ( n57387 , n57299 , n57386 );
or ( n57388 , n57298 , n57387 );
and ( n57389 , n57295 , n57388 );
or ( n57390 , n57294 , n57389 );
and ( n57391 , n57291 , n57390 );
or ( n57392 , n57290 , n57391 );
and ( n57393 , n57287 , n57392 );
or ( n57394 , n57286 , n57393 );
and ( n57395 , n57283 , n57394 );
or ( n57396 , n57282 , n57395 );
and ( n57397 , n57279 , n57396 );
or ( n57398 , n57278 , n57397 );
and ( n57399 , n57275 , n57398 );
or ( n57400 , n57274 , n57399 );
and ( n57401 , n57271 , n57400 );
or ( n57402 , n57270 , n57401 );
and ( n57403 , n57267 , n57402 );
or ( n57404 , n57266 , n57403 );
and ( n57405 , n57263 , n57404 );
or ( n57406 , n57262 , n57405 );
and ( n57407 , n57259 , n57406 );
or ( n57408 , n57258 , n57407 );
and ( n57409 , n57255 , n57408 );
or ( n57410 , n57254 , n57409 );
and ( n57411 , n57251 , n57410 );
or ( n57412 , n57250 , n57411 );
and ( n57413 , n57247 , n57412 );
or ( n57414 , n57246 , n57413 );
and ( n57415 , n57243 , n57414 );
or ( n57416 , n57242 , n57415 );
and ( n57417 , n57239 , n57416 );
or ( n57418 , n57238 , n57417 );
and ( n57419 , n57235 , n57418 );
or ( n57420 , n57234 , n57419 );
and ( n57421 , n57231 , n57420 );
or ( n57422 , n57230 , n57421 );
and ( n57423 , n57227 , n57422 );
or ( n57424 , n57226 , n57423 );
and ( n57425 , n57223 , n57424 );
or ( n57426 , n57222 , n57425 );
and ( n57427 , n57219 , n57426 );
or ( n57428 , n57218 , n57427 );
and ( n57429 , n57215 , n57428 );
or ( n57430 , n57214 , n57429 );
and ( n57431 , n57211 , n57430 );
or ( n57432 , n57210 , n57431 );
and ( n57433 , n57207 , n57432 );
or ( n57434 , n57206 , n57433 );
and ( n57435 , n57203 , n57434 );
or ( n57436 , n57202 , n57435 );
and ( n57437 , n57199 , n57436 );
or ( n57438 , n57198 , n57437 );
and ( n57439 , n57195 , n57438 );
or ( n57440 , n57194 , n57439 );
and ( n57441 , n57191 , n57440 );
or ( n57442 , n57190 , n57441 );
and ( n57443 , n57187 , n57442 );
or ( n57444 , n57186 , n57443 );
and ( n57445 , n57183 , n57444 );
or ( n57446 , n57182 , n57445 );
and ( n57447 , n57179 , n57446 );
or ( n57448 , n57178 , n57447 );
and ( n57449 , n57175 , n57448 );
or ( n57450 , n57174 , n57449 );
and ( n57451 , n57171 , n57450 );
or ( n57452 , n57170 , n57451 );
and ( n57453 , n57167 , n57452 );
or ( n57454 , n57166 , n57453 );
and ( n57455 , n57163 , n57454 );
or ( n57456 , n57162 , n57455 );
and ( n57457 , n57159 , n57456 );
or ( n57458 , n57158 , n57457 );
and ( n57459 , n57155 , n57458 );
or ( n57460 , n57154 , n57459 );
and ( n57461 , n57151 , n57460 );
or ( n57462 , n57150 , n57461 );
and ( n57463 , n57147 , n57462 );
or ( n57464 , n57146 , n57463 );
and ( n57465 , n57143 , n57464 );
or ( n57466 , n57142 , n57465 );
and ( n57467 , n57139 , n57466 );
or ( n57468 , n57138 , n57467 );
and ( n57469 , n57135 , n57468 );
or ( n57470 , n57134 , n57469 );
and ( n57471 , n57131 , n57470 );
or ( n57472 , n57130 , n57471 );
and ( n57473 , n57127 , n57472 );
or ( n57474 , n57126 , n57473 );
and ( n57475 , n57123 , n57474 );
or ( n57476 , n57122 , n57475 );
and ( n57477 , n57119 , n57476 );
or ( n57478 , n57118 , n57477 );
and ( n57479 , n57115 , n57478 );
or ( n57480 , n57114 , n57479 );
and ( n57481 , n57111 , n57480 );
or ( n57482 , n57110 , n57481 );
and ( n57483 , n57107 , n57482 );
or ( n57484 , n57106 , n57483 );
and ( n57485 , n57103 , n57484 );
or ( n57486 , n57102 , n57485 );
and ( n57487 , n57099 , n57486 );
or ( n57488 , n57098 , n57487 );
and ( n57489 , n57095 , n57488 );
or ( n57490 , n57094 , n57489 );
and ( n57491 , n57091 , n57490 );
or ( n57492 , n57090 , n57491 );
and ( n57493 , n57087 , n57492 );
or ( n57494 , n57086 , n57493 );
and ( n57495 , n57083 , n57494 );
or ( n57496 , n57082 , n57495 );
and ( n57497 , n57079 , n57496 );
or ( n57498 , n57078 , n57497 );
and ( n57499 , n57075 , n57498 );
or ( n57500 , n57074 , n57499 );
and ( n57501 , n57071 , n57500 );
or ( n57502 , n57070 , n57501 );
and ( n57503 , n57067 , n57502 );
or ( n57504 , n57066 , n57503 );
and ( n57505 , n57063 , n57504 );
or ( n57506 , n57062 , n57505 );
and ( n57507 , n57059 , n57506 );
or ( n57508 , n57058 , n57507 );
and ( n57509 , n57055 , n57508 );
or ( n57510 , n57054 , n57509 );
and ( n57511 , n57051 , n57510 );
or ( n57512 , n57050 , n57511 );
and ( n57513 , n57047 , n57512 );
or ( n57514 , n57046 , n57513 );
and ( n57515 , n57043 , n57514 );
or ( n57516 , n57042 , n57515 );
and ( n57517 , n57039 , n57516 );
or ( n57518 , n57038 , n57517 );
xor ( n57519 , n57035 , n57518 );
and ( n57520 , n33403 , n3042 );
nor ( n57521 , n3043 , n57520 );
nor ( n57522 , n3300 , n32231 );
xor ( n57523 , n57521 , n57522 );
and ( n57524 , n56319 , n56320 );
and ( n57525 , n56321 , n56324 );
or ( n57526 , n57524 , n57525 );
xor ( n57527 , n57523 , n57526 );
nor ( n57528 , n3570 , n31083 );
xor ( n57529 , n57527 , n57528 );
and ( n57530 , n56325 , n56326 );
and ( n57531 , n56327 , n56330 );
or ( n57532 , n57530 , n57531 );
xor ( n57533 , n57529 , n57532 );
nor ( n57534 , n3853 , n29948 );
xor ( n57535 , n57533 , n57534 );
and ( n57536 , n56331 , n56332 );
and ( n57537 , n56333 , n56336 );
or ( n57538 , n57536 , n57537 );
xor ( n57539 , n57535 , n57538 );
nor ( n57540 , n4151 , n28833 );
xor ( n57541 , n57539 , n57540 );
and ( n57542 , n56337 , n56338 );
and ( n57543 , n56339 , n56342 );
or ( n57544 , n57542 , n57543 );
xor ( n57545 , n57541 , n57544 );
nor ( n57546 , n4458 , n27737 );
xor ( n57547 , n57545 , n57546 );
and ( n57548 , n56343 , n56344 );
and ( n57549 , n56345 , n56348 );
or ( n57550 , n57548 , n57549 );
xor ( n57551 , n57547 , n57550 );
nor ( n57552 , n4786 , n26660 );
xor ( n57553 , n57551 , n57552 );
and ( n57554 , n56349 , n56350 );
and ( n57555 , n56351 , n56354 );
or ( n57556 , n57554 , n57555 );
xor ( n57557 , n57553 , n57556 );
nor ( n57558 , n5126 , n25600 );
xor ( n57559 , n57557 , n57558 );
and ( n57560 , n56355 , n56356 );
and ( n57561 , n56357 , n56360 );
or ( n57562 , n57560 , n57561 );
xor ( n57563 , n57559 , n57562 );
nor ( n57564 , n5477 , n24564 );
xor ( n57565 , n57563 , n57564 );
and ( n57566 , n56361 , n56362 );
and ( n57567 , n56363 , n56366 );
or ( n57568 , n57566 , n57567 );
xor ( n57569 , n57565 , n57568 );
nor ( n57570 , n5838 , n23541 );
xor ( n57571 , n57569 , n57570 );
and ( n57572 , n56367 , n56368 );
and ( n57573 , n56369 , n56372 );
or ( n57574 , n57572 , n57573 );
xor ( n57575 , n57571 , n57574 );
nor ( n57576 , n6212 , n22541 );
xor ( n57577 , n57575 , n57576 );
and ( n57578 , n56373 , n56374 );
and ( n57579 , n56375 , n56378 );
or ( n57580 , n57578 , n57579 );
xor ( n57581 , n57577 , n57580 );
nor ( n57582 , n6596 , n21562 );
xor ( n57583 , n57581 , n57582 );
and ( n57584 , n56379 , n56380 );
and ( n57585 , n56381 , n56384 );
or ( n57586 , n57584 , n57585 );
xor ( n57587 , n57583 , n57586 );
nor ( n57588 , n6997 , n20601 );
xor ( n57589 , n57587 , n57588 );
and ( n57590 , n56385 , n56386 );
and ( n57591 , n56387 , n56390 );
or ( n57592 , n57590 , n57591 );
xor ( n57593 , n57589 , n57592 );
nor ( n57594 , n7413 , n19657 );
xor ( n57595 , n57593 , n57594 );
and ( n57596 , n56391 , n56392 );
and ( n57597 , n56393 , n56396 );
or ( n57598 , n57596 , n57597 );
xor ( n57599 , n57595 , n57598 );
nor ( n57600 , n7841 , n18734 );
xor ( n57601 , n57599 , n57600 );
and ( n57602 , n56397 , n56398 );
and ( n57603 , n56399 , n56402 );
or ( n57604 , n57602 , n57603 );
xor ( n57605 , n57601 , n57604 );
nor ( n57606 , n8281 , n17828 );
xor ( n57607 , n57605 , n57606 );
and ( n57608 , n56403 , n56404 );
and ( n57609 , n56405 , n56408 );
or ( n57610 , n57608 , n57609 );
xor ( n57611 , n57607 , n57610 );
nor ( n57612 , n8737 , n16943 );
xor ( n57613 , n57611 , n57612 );
and ( n57614 , n56409 , n56410 );
and ( n57615 , n56411 , n56414 );
or ( n57616 , n57614 , n57615 );
xor ( n57617 , n57613 , n57616 );
nor ( n57618 , n9420 , n16077 );
xor ( n57619 , n57617 , n57618 );
and ( n57620 , n56415 , n56416 );
and ( n57621 , n56417 , n56420 );
or ( n57622 , n57620 , n57621 );
xor ( n57623 , n57619 , n57622 );
nor ( n57624 , n10312 , n15230 );
xor ( n57625 , n57623 , n57624 );
and ( n57626 , n56421 , n56422 );
and ( n57627 , n56423 , n56426 );
or ( n57628 , n57626 , n57627 );
xor ( n57629 , n57625 , n57628 );
nor ( n57630 , n11041 , n14403 );
xor ( n57631 , n57629 , n57630 );
and ( n57632 , n56427 , n56428 );
and ( n57633 , n56429 , n56432 );
or ( n57634 , n57632 , n57633 );
xor ( n57635 , n57631 , n57634 );
nor ( n57636 , n11790 , n13599 );
xor ( n57637 , n57635 , n57636 );
and ( n57638 , n56433 , n56434 );
and ( n57639 , n56435 , n56438 );
or ( n57640 , n57638 , n57639 );
xor ( n57641 , n57637 , n57640 );
nor ( n57642 , n12555 , n12808 );
xor ( n57643 , n57641 , n57642 );
and ( n57644 , n56439 , n56440 );
and ( n57645 , n56441 , n56444 );
or ( n57646 , n57644 , n57645 );
xor ( n57647 , n57643 , n57646 );
nor ( n57648 , n13340 , n12037 );
xor ( n57649 , n57647 , n57648 );
and ( n57650 , n56445 , n56446 );
and ( n57651 , n56447 , n56450 );
or ( n57652 , n57650 , n57651 );
xor ( n57653 , n57649 , n57652 );
nor ( n57654 , n14138 , n11282 );
xor ( n57655 , n57653 , n57654 );
and ( n57656 , n56451 , n56452 );
and ( n57657 , n56453 , n56456 );
or ( n57658 , n57656 , n57657 );
xor ( n57659 , n57655 , n57658 );
nor ( n57660 , n14959 , n10547 );
xor ( n57661 , n57659 , n57660 );
and ( n57662 , n56457 , n56458 );
and ( n57663 , n56459 , n56462 );
or ( n57664 , n57662 , n57663 );
xor ( n57665 , n57661 , n57664 );
nor ( n57666 , n15800 , n9829 );
xor ( n57667 , n57665 , n57666 );
and ( n57668 , n56463 , n56464 );
and ( n57669 , n56465 , n56468 );
or ( n57670 , n57668 , n57669 );
xor ( n57671 , n57667 , n57670 );
nor ( n57672 , n16660 , n8955 );
xor ( n57673 , n57671 , n57672 );
and ( n57674 , n56469 , n56470 );
and ( n57675 , n56471 , n56474 );
or ( n57676 , n57674 , n57675 );
xor ( n57677 , n57673 , n57676 );
nor ( n57678 , n17539 , n603 );
xor ( n57679 , n57677 , n57678 );
and ( n57680 , n56475 , n56476 );
and ( n57681 , n56477 , n56480 );
or ( n57682 , n57680 , n57681 );
xor ( n57683 , n57679 , n57682 );
nor ( n57684 , n18439 , n652 );
xor ( n57685 , n57683 , n57684 );
and ( n57686 , n56481 , n56482 );
and ( n57687 , n56483 , n56486 );
or ( n57688 , n57686 , n57687 );
xor ( n57689 , n57685 , n57688 );
nor ( n57690 , n19356 , n624 );
xor ( n57691 , n57689 , n57690 );
and ( n57692 , n56487 , n56488 );
and ( n57693 , n56489 , n56492 );
or ( n57694 , n57692 , n57693 );
xor ( n57695 , n57691 , n57694 );
nor ( n57696 , n20294 , n648 );
xor ( n57697 , n57695 , n57696 );
and ( n57698 , n56493 , n56494 );
and ( n57699 , n56495 , n56498 );
or ( n57700 , n57698 , n57699 );
xor ( n57701 , n57697 , n57700 );
nor ( n57702 , n21249 , n686 );
xor ( n57703 , n57701 , n57702 );
and ( n57704 , n56499 , n56500 );
and ( n57705 , n56501 , n56504 );
or ( n57706 , n57704 , n57705 );
xor ( n57707 , n57703 , n57706 );
nor ( n57708 , n22222 , n735 );
xor ( n57709 , n57707 , n57708 );
and ( n57710 , n56505 , n56506 );
and ( n57711 , n56507 , n56510 );
or ( n57712 , n57710 , n57711 );
xor ( n57713 , n57709 , n57712 );
nor ( n57714 , n23216 , n798 );
xor ( n57715 , n57713 , n57714 );
and ( n57716 , n56511 , n56512 );
and ( n57717 , n56513 , n56516 );
or ( n57718 , n57716 , n57717 );
xor ( n57719 , n57715 , n57718 );
nor ( n57720 , n24233 , n870 );
xor ( n57721 , n57719 , n57720 );
and ( n57722 , n56517 , n56518 );
and ( n57723 , n56519 , n56522 );
or ( n57724 , n57722 , n57723 );
xor ( n57725 , n57721 , n57724 );
nor ( n57726 , n25263 , n960 );
xor ( n57727 , n57725 , n57726 );
and ( n57728 , n56523 , n56524 );
and ( n57729 , n56525 , n56528 );
or ( n57730 , n57728 , n57729 );
xor ( n57731 , n57727 , n57730 );
nor ( n57732 , n26317 , n1064 );
xor ( n57733 , n57731 , n57732 );
and ( n57734 , n56529 , n56530 );
and ( n57735 , n56531 , n56534 );
or ( n57736 , n57734 , n57735 );
xor ( n57737 , n57733 , n57736 );
nor ( n57738 , n27388 , n1178 );
xor ( n57739 , n57737 , n57738 );
and ( n57740 , n56535 , n56536 );
and ( n57741 , n56537 , n56540 );
or ( n57742 , n57740 , n57741 );
xor ( n57743 , n57739 , n57742 );
nor ( n57744 , n28478 , n1305 );
xor ( n57745 , n57743 , n57744 );
and ( n57746 , n56541 , n56542 );
and ( n57747 , n56543 , n56546 );
or ( n57748 , n57746 , n57747 );
xor ( n57749 , n57745 , n57748 );
nor ( n57750 , n29587 , n1447 );
xor ( n57751 , n57749 , n57750 );
and ( n57752 , n56547 , n56548 );
and ( n57753 , n56549 , n56552 );
or ( n57754 , n57752 , n57753 );
xor ( n57755 , n57751 , n57754 );
nor ( n57756 , n30716 , n1600 );
xor ( n57757 , n57755 , n57756 );
and ( n57758 , n56553 , n56554 );
and ( n57759 , n56555 , n56558 );
or ( n57760 , n57758 , n57759 );
xor ( n57761 , n57757 , n57760 );
nor ( n57762 , n31858 , n1768 );
xor ( n57763 , n57761 , n57762 );
and ( n57764 , n56559 , n56560 );
and ( n57765 , n56561 , n56564 );
or ( n57766 , n57764 , n57765 );
xor ( n57767 , n57763 , n57766 );
nor ( n57768 , n33024 , n1947 );
xor ( n57769 , n57767 , n57768 );
and ( n57770 , n56565 , n56566 );
and ( n57771 , n56567 , n56570 );
or ( n57772 , n57770 , n57771 );
xor ( n57773 , n57769 , n57772 );
nor ( n57774 , n34215 , n2139 );
xor ( n57775 , n57773 , n57774 );
and ( n57776 , n56571 , n56572 );
and ( n57777 , n56573 , n56576 );
or ( n57778 , n57776 , n57777 );
xor ( n57779 , n57775 , n57778 );
nor ( n57780 , n35410 , n2345 );
xor ( n57781 , n57779 , n57780 );
and ( n57782 , n56577 , n56578 );
and ( n57783 , n56579 , n56582 );
or ( n57784 , n57782 , n57783 );
xor ( n57785 , n57781 , n57784 );
nor ( n57786 , n36611 , n2568 );
xor ( n57787 , n57785 , n57786 );
and ( n57788 , n56583 , n56584 );
and ( n57789 , n56585 , n56588 );
or ( n57790 , n57788 , n57789 );
xor ( n57791 , n57787 , n57790 );
nor ( n57792 , n37816 , n2799 );
xor ( n57793 , n57791 , n57792 );
and ( n57794 , n56589 , n56590 );
and ( n57795 , n56591 , n56594 );
or ( n57796 , n57794 , n57795 );
xor ( n57797 , n57793 , n57796 );
nor ( n57798 , n39018 , n3045 );
xor ( n57799 , n57797 , n57798 );
and ( n57800 , n56595 , n56596 );
and ( n57801 , n56597 , n56600 );
or ( n57802 , n57800 , n57801 );
xor ( n57803 , n57799 , n57802 );
nor ( n57804 , n40223 , n3302 );
xor ( n57805 , n57803 , n57804 );
and ( n57806 , n56601 , n56602 );
and ( n57807 , n56603 , n56606 );
or ( n57808 , n57806 , n57807 );
xor ( n57809 , n57805 , n57808 );
nor ( n57810 , n41428 , n3572 );
xor ( n57811 , n57809 , n57810 );
and ( n57812 , n56607 , n56608 );
and ( n57813 , n56609 , n56612 );
or ( n57814 , n57812 , n57813 );
xor ( n57815 , n57811 , n57814 );
nor ( n57816 , n42632 , n3855 );
xor ( n57817 , n57815 , n57816 );
and ( n57818 , n56613 , n56614 );
and ( n57819 , n56615 , n56618 );
or ( n57820 , n57818 , n57819 );
xor ( n57821 , n57817 , n57820 );
nor ( n57822 , n43834 , n4153 );
xor ( n57823 , n57821 , n57822 );
and ( n57824 , n56619 , n56620 );
and ( n57825 , n56621 , n56624 );
or ( n57826 , n57824 , n57825 );
xor ( n57827 , n57823 , n57826 );
nor ( n57828 , n45038 , n4460 );
xor ( n57829 , n57827 , n57828 );
and ( n57830 , n56625 , n56626 );
and ( n57831 , n56627 , n56630 );
or ( n57832 , n57830 , n57831 );
xor ( n57833 , n57829 , n57832 );
nor ( n57834 , n46239 , n4788 );
xor ( n57835 , n57833 , n57834 );
and ( n57836 , n56631 , n56632 );
and ( n57837 , n56633 , n56636 );
or ( n57838 , n57836 , n57837 );
xor ( n57839 , n57835 , n57838 );
nor ( n57840 , n47440 , n5128 );
xor ( n57841 , n57839 , n57840 );
and ( n57842 , n56637 , n56638 );
and ( n57843 , n56639 , n56642 );
or ( n57844 , n57842 , n57843 );
xor ( n57845 , n57841 , n57844 );
nor ( n57846 , n48641 , n5479 );
xor ( n57847 , n57845 , n57846 );
and ( n57848 , n56643 , n56644 );
and ( n57849 , n56645 , n56648 );
or ( n57850 , n57848 , n57849 );
xor ( n57851 , n57847 , n57850 );
nor ( n57852 , n49841 , n5840 );
xor ( n57853 , n57851 , n57852 );
and ( n57854 , n56649 , n56650 );
and ( n57855 , n56651 , n56654 );
or ( n57856 , n57854 , n57855 );
xor ( n57857 , n57853 , n57856 );
nor ( n57858 , n51040 , n6214 );
xor ( n57859 , n57857 , n57858 );
and ( n57860 , n56655 , n56656 );
and ( n57861 , n56657 , n56660 );
or ( n57862 , n57860 , n57861 );
xor ( n57863 , n57859 , n57862 );
nor ( n57864 , n52238 , n6598 );
xor ( n57865 , n57863 , n57864 );
and ( n57866 , n56661 , n56662 );
and ( n57867 , n56663 , n56666 );
or ( n57868 , n57866 , n57867 );
xor ( n57869 , n57865 , n57868 );
nor ( n57870 , n53432 , n6999 );
xor ( n57871 , n57869 , n57870 );
and ( n57872 , n56667 , n56668 );
and ( n57873 , n56669 , n56672 );
or ( n57874 , n57872 , n57873 );
xor ( n57875 , n57871 , n57874 );
nor ( n57876 , n54629 , n7415 );
xor ( n57877 , n57875 , n57876 );
and ( n57878 , n56673 , n56674 );
and ( n57879 , n56675 , n56678 );
or ( n57880 , n57878 , n57879 );
xor ( n57881 , n57877 , n57880 );
nor ( n57882 , n55826 , n7843 );
xor ( n57883 , n57881 , n57882 );
and ( n57884 , n56679 , n56680 );
and ( n57885 , n56681 , n56684 );
or ( n57886 , n57884 , n57885 );
xor ( n57887 , n57883 , n57886 );
nor ( n57888 , n57022 , n8283 );
xor ( n57889 , n57887 , n57888 );
and ( n57890 , n56685 , n56686 );
and ( n57891 , n56687 , n56690 );
or ( n57892 , n57890 , n57891 );
xor ( n57893 , n57889 , n57892 );
and ( n57894 , n56703 , n56707 );
and ( n57895 , n56707 , n57008 );
and ( n57896 , n56703 , n57008 );
or ( n57897 , n57894 , n57895 , n57896 );
and ( n57898 , n33774 , n2981 );
not ( n57899 , n2981 );
nor ( n57900 , n57898 , n57899 );
xor ( n57901 , n57897 , n57900 );
and ( n57902 , n56716 , n56720 );
and ( n57903 , n56720 , n56788 );
and ( n57904 , n56716 , n56788 );
or ( n57905 , n57902 , n57903 , n57904 );
and ( n57906 , n56712 , n56789 );
and ( n57907 , n56789 , n57007 );
and ( n57908 , n56712 , n57007 );
or ( n57909 , n57906 , n57907 , n57908 );
xor ( n57910 , n57905 , n57909 );
and ( n57911 , n56791 , n56911 );
and ( n57912 , n56911 , n57006 );
and ( n57913 , n56791 , n57006 );
or ( n57914 , n57911 , n57912 , n57913 );
and ( n57915 , n56725 , n56729 );
and ( n57916 , n56729 , n56787 );
and ( n57917 , n56725 , n56787 );
or ( n57918 , n57915 , n57916 , n57917 );
and ( n57919 , n56795 , n56799 );
and ( n57920 , n56799 , n56910 );
and ( n57921 , n56795 , n56910 );
or ( n57922 , n57919 , n57920 , n57921 );
xor ( n57923 , n57918 , n57922 );
and ( n57924 , n56756 , n56760 );
and ( n57925 , n56760 , n56766 );
and ( n57926 , n56756 , n56766 );
or ( n57927 , n57924 , n57925 , n57926 );
and ( n57928 , n56734 , n56738 );
and ( n57929 , n56738 , n56786 );
and ( n57930 , n56734 , n56786 );
or ( n57931 , n57928 , n57929 , n57930 );
xor ( n57932 , n57927 , n57931 );
and ( n57933 , n56743 , n56747 );
and ( n57934 , n56747 , n56785 );
and ( n57935 , n56743 , n56785 );
or ( n57936 , n57933 , n57934 , n57935 );
and ( n57937 , n56808 , n56833 );
and ( n57938 , n56833 , n56871 );
and ( n57939 , n56808 , n56871 );
or ( n57940 , n57937 , n57938 , n57939 );
xor ( n57941 , n57936 , n57940 );
and ( n57942 , n56752 , n56767 );
and ( n57943 , n56767 , n56784 );
and ( n57944 , n56752 , n56784 );
or ( n57945 , n57942 , n57943 , n57944 );
and ( n57946 , n56812 , n56816 );
and ( n57947 , n56816 , n56832 );
and ( n57948 , n56812 , n56832 );
or ( n57949 , n57946 , n57947 , n57948 );
xor ( n57950 , n57945 , n57949 );
and ( n57951 , n56772 , n56777 );
and ( n57952 , n56777 , n56783 );
and ( n57953 , n56772 , n56783 );
or ( n57954 , n57951 , n57952 , n57953 );
and ( n57955 , n56762 , n56763 );
and ( n57956 , n56763 , n56765 );
and ( n57957 , n56762 , n56765 );
or ( n57958 , n57955 , n57956 , n57957 );
and ( n57959 , n56773 , n56774 );
and ( n57960 , n56774 , n56776 );
and ( n57961 , n56773 , n56776 );
or ( n57962 , n57959 , n57960 , n57961 );
xor ( n57963 , n57958 , n57962 );
and ( n57964 , n30695 , n3749 );
and ( n57965 , n31836 , n3495 );
xor ( n57966 , n57964 , n57965 );
and ( n57967 , n32649 , n3271 );
xor ( n57968 , n57966 , n57967 );
xor ( n57969 , n57963 , n57968 );
xor ( n57970 , n57954 , n57969 );
and ( n57971 , n56779 , n56780 );
and ( n57972 , n56780 , n56782 );
and ( n57973 , n56779 , n56782 );
or ( n57974 , n57971 , n57972 , n57973 );
and ( n57975 , n27361 , n4730 );
and ( n57976 , n28456 , n4403 );
xor ( n57977 , n57975 , n57976 );
and ( n57978 , n29559 , n4102 );
xor ( n57979 , n57977 , n57978 );
xor ( n57980 , n57974 , n57979 );
and ( n57981 , n24214 , n5765 );
and ( n57982 , n25243 , n5408 );
xor ( n57983 , n57981 , n57982 );
and ( n57984 , n26296 , n5103 );
xor ( n57985 , n57983 , n57984 );
xor ( n57986 , n57980 , n57985 );
xor ( n57987 , n57970 , n57986 );
xor ( n57988 , n57950 , n57987 );
xor ( n57989 , n57941 , n57988 );
xor ( n57990 , n57932 , n57989 );
xor ( n57991 , n57923 , n57990 );
xor ( n57992 , n57914 , n57991 );
and ( n57993 , n56987 , n57005 );
and ( n57994 , n56916 , n56917 );
and ( n57995 , n56917 , n56986 );
and ( n57996 , n56916 , n56986 );
or ( n57997 , n57994 , n57995 , n57996 );
and ( n57998 , n56804 , n56872 );
and ( n57999 , n56872 , n56909 );
and ( n58000 , n56804 , n56909 );
or ( n58001 , n57998 , n57999 , n58000 );
xor ( n58002 , n57997 , n58001 );
and ( n58003 , n56877 , n56881 );
and ( n58004 , n56881 , n56908 );
and ( n58005 , n56877 , n56908 );
or ( n58006 , n58003 , n58004 , n58005 );
and ( n58007 , n56838 , n56854 );
and ( n58008 , n56854 , n56870 );
and ( n58009 , n56838 , n56870 );
or ( n58010 , n58007 , n58008 , n58009 );
and ( n58011 , n56821 , n56825 );
and ( n58012 , n56825 , n56831 );
and ( n58013 , n56821 , n56831 );
or ( n58014 , n58011 , n58012 , n58013 );
and ( n58015 , n56842 , n56847 );
and ( n58016 , n56847 , n56853 );
and ( n58017 , n56842 , n56853 );
or ( n58018 , n58015 , n58016 , n58017 );
xor ( n58019 , n58014 , n58018 );
and ( n58020 , n56827 , n56828 );
and ( n58021 , n56828 , n56830 );
and ( n58022 , n56827 , n56830 );
or ( n58023 , n58020 , n58021 , n58022 );
and ( n58024 , n56843 , n56844 );
and ( n58025 , n56844 , n56846 );
and ( n58026 , n56843 , n56846 );
or ( n58027 , n58024 , n58025 , n58026 );
xor ( n58028 , n58023 , n58027 );
and ( n58029 , n21216 , n6971 );
and ( n58030 , n22186 , n6504 );
xor ( n58031 , n58029 , n58030 );
and ( n58032 , n22892 , n6132 );
xor ( n58033 , n58031 , n58032 );
xor ( n58034 , n58028 , n58033 );
xor ( n58035 , n58019 , n58034 );
xor ( n58036 , n58010 , n58035 );
and ( n58037 , n56859 , n56863 );
and ( n58038 , n56863 , n56869 );
and ( n58039 , n56859 , n56869 );
or ( n58040 , n58037 , n58038 , n58039 );
and ( n58041 , n56849 , n56850 );
and ( n58042 , n56850 , n56852 );
and ( n58043 , n56849 , n56852 );
or ( n58044 , n58041 , n58042 , n58043 );
and ( n58045 , n18144 , n8243 );
and ( n58046 , n19324 , n7662 );
xor ( n58047 , n58045 , n58046 );
and ( n58048 , n20233 , n7310 );
xor ( n58049 , n58047 , n58048 );
xor ( n58050 , n58044 , n58049 );
and ( n58051 , n15758 , n10239 );
and ( n58052 , n16637 , n9348 );
xor ( n58053 , n58051 , n58052 );
and ( n58054 , n17512 , n8669 );
xor ( n58055 , n58053 , n58054 );
xor ( n58056 , n58050 , n58055 );
xor ( n58057 , n58040 , n58056 );
and ( n58058 , n56865 , n56866 );
and ( n58059 , n56866 , n56868 );
and ( n58060 , n56865 , n56868 );
or ( n58061 , n58058 , n58059 , n58060 );
and ( n58062 , n56896 , n56897 );
and ( n58063 , n56897 , n56899 );
and ( n58064 , n56896 , n56899 );
or ( n58065 , n58062 , n58063 , n58064 );
xor ( n58066 , n58061 , n58065 );
and ( n58067 , n13322 , n12531 );
and ( n58068 , n14118 , n11718 );
xor ( n58069 , n58067 , n58068 );
and ( n58070 , n14938 , n10977 );
xor ( n58071 , n58069 , n58070 );
xor ( n58072 , n58066 , n58071 );
xor ( n58073 , n58057 , n58072 );
xor ( n58074 , n58036 , n58073 );
xor ( n58075 , n58006 , n58074 );
and ( n58076 , n56886 , n56890 );
and ( n58077 , n56890 , n56907 );
and ( n58078 , n56886 , n56907 );
or ( n58079 , n58076 , n58077 , n58078 );
and ( n58080 , n56926 , n56941 );
and ( n58081 , n56941 , n56958 );
and ( n58082 , n56926 , n56958 );
or ( n58083 , n58080 , n58081 , n58082 );
xor ( n58084 , n58079 , n58083 );
and ( n58085 , n56895 , n56900 );
and ( n58086 , n56900 , n56906 );
and ( n58087 , n56895 , n56906 );
or ( n58088 , n58085 , n58086 , n58087 );
and ( n58089 , n56930 , n56934 );
and ( n58090 , n56934 , n56940 );
and ( n58091 , n56930 , n56940 );
or ( n58092 , n58089 , n58090 , n58091 );
xor ( n58093 , n58088 , n58092 );
and ( n58094 , n56902 , n56903 );
and ( n58095 , n56903 , n56905 );
and ( n58096 , n56902 , n56905 );
or ( n58097 , n58094 , n58095 , n58096 );
and ( n58098 , n11015 , n14838 );
and ( n58099 , n11769 , n14044 );
xor ( n58100 , n58098 , n58099 );
and ( n58101 , n12320 , n13256 );
xor ( n58102 , n58100 , n58101 );
xor ( n58103 , n58097 , n58102 );
and ( n58104 , n8718 , n17422 );
and ( n58105 , n9400 , n16550 );
xor ( n58106 , n58104 , n58105 );
and ( n58107 , n10291 , n15691 );
xor ( n58108 , n58106 , n58107 );
xor ( n58109 , n58103 , n58108 );
xor ( n58110 , n58093 , n58109 );
xor ( n58111 , n58084 , n58110 );
xor ( n58112 , n58075 , n58111 );
xor ( n58113 , n58002 , n58112 );
xor ( n58114 , n57993 , n58113 );
and ( n58115 , n57001 , n57002 );
not ( n58116 , n3024 );
and ( n58117 , n34193 , n3024 );
nor ( n58118 , n58116 , n58117 );
xor ( n58119 , n58115 , n58118 );
and ( n58120 , n3182 , n32999 );
and ( n58121 , n3545 , n31761 );
xor ( n58122 , n58120 , n58121 );
and ( n58123 , n3801 , n30629 );
xor ( n58124 , n58122 , n58123 );
xor ( n58125 , n58119 , n58124 );
and ( n58126 , n56922 , n56959 );
and ( n58127 , n56959 , n56985 );
and ( n58128 , n56922 , n56985 );
or ( n58129 , n58126 , n58127 , n58128 );
and ( n58130 , n56988 , n57004 );
xor ( n58131 , n58129 , n58130 );
and ( n58132 , n56964 , n56968 );
and ( n58133 , n56968 , n56984 );
and ( n58134 , n56964 , n56984 );
or ( n58135 , n58132 , n58133 , n58134 );
and ( n58136 , n56946 , n56951 );
and ( n58137 , n56951 , n56957 );
and ( n58138 , n56946 , n56957 );
or ( n58139 , n58136 , n58137 , n58138 );
and ( n58140 , n56936 , n56937 );
and ( n58141 , n56937 , n56939 );
and ( n58142 , n56936 , n56939 );
or ( n58143 , n58140 , n58141 , n58142 );
and ( n58144 , n56947 , n56948 );
and ( n58145 , n56948 , n56950 );
and ( n58146 , n56947 , n56950 );
or ( n58147 , n58144 , n58145 , n58146 );
xor ( n58148 , n58143 , n58147 );
and ( n58149 , n7385 , n20156 );
and ( n58150 , n7808 , n19222 );
xor ( n58151 , n58149 , n58150 );
and ( n58152 , n8079 , n18407 );
xor ( n58153 , n58151 , n58152 );
xor ( n58154 , n58148 , n58153 );
xor ( n58155 , n58139 , n58154 );
and ( n58156 , n56953 , n56954 );
and ( n58157 , n56954 , n56956 );
and ( n58158 , n56953 , n56956 );
or ( n58159 , n58156 , n58157 , n58158 );
and ( n58160 , n6187 , n23075 );
and ( n58161 , n6569 , n22065 );
xor ( n58162 , n58160 , n58161 );
and ( n58163 , n6816 , n20976 );
xor ( n58164 , n58162 , n58163 );
xor ( n58165 , n58159 , n58164 );
and ( n58166 , n4959 , n26216 );
and ( n58167 , n5459 , n25163 );
xor ( n58168 , n58166 , n58167 );
and ( n58169 , n5819 , n24137 );
xor ( n58170 , n58168 , n58169 );
xor ( n58171 , n58165 , n58170 );
xor ( n58172 , n58155 , n58171 );
xor ( n58173 , n58135 , n58172 );
and ( n58174 , n56973 , n56977 );
and ( n58175 , n56977 , n56983 );
and ( n58176 , n56973 , n56983 );
or ( n58177 , n58174 , n58175 , n58176 );
and ( n58178 , n56992 , n56997 );
and ( n58179 , n56997 , n57003 );
and ( n58180 , n56992 , n57003 );
or ( n58181 , n58178 , n58179 , n58180 );
xor ( n58182 , n58177 , n58181 );
and ( n58183 , n56979 , n56980 );
and ( n58184 , n56980 , n56982 );
and ( n58185 , n56979 , n56982 );
or ( n58186 , n58183 , n58184 , n58185 );
and ( n58187 , n56993 , n56994 );
and ( n58188 , n56994 , n56996 );
and ( n58189 , n56993 , n56996 );
or ( n58190 , n58187 , n58188 , n58189 );
xor ( n58191 , n58186 , n58190 );
and ( n58192 , n4132 , n29508 );
and ( n58193 , n4438 , n28406 );
xor ( n58194 , n58192 , n58193 );
and ( n58195 , n4766 , n27296 );
xor ( n58196 , n58194 , n58195 );
xor ( n58197 , n58191 , n58196 );
xor ( n58198 , n58182 , n58197 );
xor ( n58199 , n58173 , n58198 );
xor ( n58200 , n58131 , n58199 );
xor ( n58201 , n58125 , n58200 );
xor ( n58202 , n58114 , n58201 );
xor ( n58203 , n57992 , n58202 );
xor ( n58204 , n57910 , n58203 );
xor ( n58205 , n57901 , n58204 );
and ( n58206 , n56695 , n56698 );
and ( n58207 , n56698 , n57009 );
and ( n58208 , n56695 , n57009 );
or ( n58209 , n58206 , n58207 , n58208 );
xor ( n58210 , n58205 , n58209 );
and ( n58211 , n57010 , n57014 );
and ( n58212 , n57015 , n57018 );
or ( n58213 , n58211 , n58212 );
xor ( n58214 , n58210 , n58213 );
buf ( n58215 , n58214 );
buf ( n58216 , n58215 );
not ( n58217 , n58216 );
nor ( n58218 , n58217 , n8739 );
xor ( n58219 , n57893 , n58218 );
and ( n58220 , n56691 , n57023 );
and ( n58221 , n57024 , n57027 );
or ( n58222 , n58220 , n58221 );
xor ( n58223 , n58219 , n58222 );
buf ( n58224 , n58223 );
buf ( n58225 , n58224 );
not ( n58226 , n58225 );
buf ( n58227 , n582 );
not ( n58228 , n58227 );
nor ( n58229 , n58226 , n58228 );
xor ( n58230 , n57519 , n58229 );
xor ( n58231 , n57039 , n57516 );
nor ( n58232 , n57031 , n58228 );
and ( n58233 , n58231 , n58232 );
xor ( n58234 , n58231 , n58232 );
xor ( n58235 , n57043 , n57514 );
nor ( n58236 , n55835 , n58228 );
and ( n58237 , n58235 , n58236 );
xor ( n58238 , n58235 , n58236 );
xor ( n58239 , n57047 , n57512 );
nor ( n58240 , n54638 , n58228 );
and ( n58241 , n58239 , n58240 );
xor ( n58242 , n58239 , n58240 );
xor ( n58243 , n57051 , n57510 );
nor ( n58244 , n53441 , n58228 );
and ( n58245 , n58243 , n58244 );
xor ( n58246 , n58243 , n58244 );
xor ( n58247 , n57055 , n57508 );
nor ( n58248 , n52247 , n58228 );
and ( n58249 , n58247 , n58248 );
xor ( n58250 , n58247 , n58248 );
xor ( n58251 , n57059 , n57506 );
nor ( n58252 , n51049 , n58228 );
and ( n58253 , n58251 , n58252 );
xor ( n58254 , n58251 , n58252 );
xor ( n58255 , n57063 , n57504 );
nor ( n58256 , n49850 , n58228 );
and ( n58257 , n58255 , n58256 );
xor ( n58258 , n58255 , n58256 );
xor ( n58259 , n57067 , n57502 );
nor ( n58260 , n48650 , n58228 );
and ( n58261 , n58259 , n58260 );
xor ( n58262 , n58259 , n58260 );
xor ( n58263 , n57071 , n57500 );
nor ( n58264 , n47449 , n58228 );
and ( n58265 , n58263 , n58264 );
xor ( n58266 , n58263 , n58264 );
xor ( n58267 , n57075 , n57498 );
nor ( n58268 , n46248 , n58228 );
and ( n58269 , n58267 , n58268 );
xor ( n58270 , n58267 , n58268 );
xor ( n58271 , n57079 , n57496 );
nor ( n58272 , n45047 , n58228 );
and ( n58273 , n58271 , n58272 );
xor ( n58274 , n58271 , n58272 );
xor ( n58275 , n57083 , n57494 );
nor ( n58276 , n43843 , n58228 );
and ( n58277 , n58275 , n58276 );
xor ( n58278 , n58275 , n58276 );
xor ( n58279 , n57087 , n57492 );
nor ( n58280 , n42641 , n58228 );
and ( n58281 , n58279 , n58280 );
xor ( n58282 , n58279 , n58280 );
xor ( n58283 , n57091 , n57490 );
nor ( n58284 , n41437 , n58228 );
and ( n58285 , n58283 , n58284 );
xor ( n58286 , n58283 , n58284 );
xor ( n58287 , n57095 , n57488 );
nor ( n58288 , n40232 , n58228 );
and ( n58289 , n58287 , n58288 );
xor ( n58290 , n58287 , n58288 );
xor ( n58291 , n57099 , n57486 );
nor ( n58292 , n39027 , n58228 );
and ( n58293 , n58291 , n58292 );
xor ( n58294 , n58291 , n58292 );
xor ( n58295 , n57103 , n57484 );
nor ( n58296 , n37825 , n58228 );
and ( n58297 , n58295 , n58296 );
xor ( n58298 , n58295 , n58296 );
xor ( n58299 , n57107 , n57482 );
nor ( n58300 , n36620 , n58228 );
and ( n58301 , n58299 , n58300 );
xor ( n58302 , n58299 , n58300 );
xor ( n58303 , n57111 , n57480 );
nor ( n58304 , n35419 , n58228 );
and ( n58305 , n58303 , n58304 );
xor ( n58306 , n58303 , n58304 );
xor ( n58307 , n57115 , n57478 );
nor ( n58308 , n34224 , n58228 );
and ( n58309 , n58307 , n58308 );
xor ( n58310 , n58307 , n58308 );
xor ( n58311 , n57119 , n57476 );
nor ( n58312 , n33033 , n58228 );
and ( n58313 , n58311 , n58312 );
xor ( n58314 , n58311 , n58312 );
xor ( n58315 , n57123 , n57474 );
nor ( n58316 , n31867 , n58228 );
and ( n58317 , n58315 , n58316 );
xor ( n58318 , n58315 , n58316 );
xor ( n58319 , n57127 , n57472 );
nor ( n58320 , n30725 , n58228 );
and ( n58321 , n58319 , n58320 );
xor ( n58322 , n58319 , n58320 );
xor ( n58323 , n57131 , n57470 );
nor ( n58324 , n29596 , n58228 );
and ( n58325 , n58323 , n58324 );
xor ( n58326 , n58323 , n58324 );
xor ( n58327 , n57135 , n57468 );
nor ( n58328 , n28487 , n58228 );
and ( n58329 , n58327 , n58328 );
xor ( n58330 , n58327 , n58328 );
xor ( n58331 , n57139 , n57466 );
nor ( n58332 , n27397 , n58228 );
and ( n58333 , n58331 , n58332 );
xor ( n58334 , n58331 , n58332 );
xor ( n58335 , n57143 , n57464 );
nor ( n58336 , n26326 , n58228 );
and ( n58337 , n58335 , n58336 );
xor ( n58338 , n58335 , n58336 );
xor ( n58339 , n57147 , n57462 );
nor ( n58340 , n25272 , n58228 );
and ( n58341 , n58339 , n58340 );
xor ( n58342 , n58339 , n58340 );
xor ( n58343 , n57151 , n57460 );
nor ( n58344 , n24242 , n58228 );
and ( n58345 , n58343 , n58344 );
xor ( n58346 , n58343 , n58344 );
xor ( n58347 , n57155 , n57458 );
nor ( n58348 , n23225 , n58228 );
and ( n58349 , n58347 , n58348 );
xor ( n58350 , n58347 , n58348 );
xor ( n58351 , n57159 , n57456 );
nor ( n58352 , n22231 , n58228 );
and ( n58353 , n58351 , n58352 );
xor ( n58354 , n58351 , n58352 );
xor ( n58355 , n57163 , n57454 );
nor ( n58356 , n21258 , n58228 );
and ( n58357 , n58355 , n58356 );
xor ( n58358 , n58355 , n58356 );
xor ( n58359 , n57167 , n57452 );
nor ( n58360 , n20303 , n58228 );
and ( n58361 , n58359 , n58360 );
xor ( n58362 , n58359 , n58360 );
xor ( n58363 , n57171 , n57450 );
nor ( n58364 , n19365 , n58228 );
and ( n58365 , n58363 , n58364 );
xor ( n58366 , n58363 , n58364 );
xor ( n58367 , n57175 , n57448 );
nor ( n58368 , n18448 , n58228 );
and ( n58369 , n58367 , n58368 );
xor ( n58370 , n58367 , n58368 );
xor ( n58371 , n57179 , n57446 );
nor ( n58372 , n17548 , n58228 );
and ( n58373 , n58371 , n58372 );
xor ( n58374 , n58371 , n58372 );
xor ( n58375 , n57183 , n57444 );
nor ( n58376 , n16669 , n58228 );
and ( n58377 , n58375 , n58376 );
xor ( n58378 , n58375 , n58376 );
xor ( n58379 , n57187 , n57442 );
nor ( n58380 , n15809 , n58228 );
and ( n58381 , n58379 , n58380 );
xor ( n58382 , n58379 , n58380 );
xor ( n58383 , n57191 , n57440 );
nor ( n58384 , n14968 , n58228 );
and ( n58385 , n58383 , n58384 );
xor ( n58386 , n58383 , n58384 );
xor ( n58387 , n57195 , n57438 );
nor ( n58388 , n14147 , n58228 );
and ( n58389 , n58387 , n58388 );
xor ( n58390 , n58387 , n58388 );
xor ( n58391 , n57199 , n57436 );
nor ( n58392 , n13349 , n58228 );
and ( n58393 , n58391 , n58392 );
xor ( n58394 , n58391 , n58392 );
xor ( n58395 , n57203 , n57434 );
nor ( n58396 , n12564 , n58228 );
and ( n58397 , n58395 , n58396 );
xor ( n58398 , n58395 , n58396 );
xor ( n58399 , n57207 , n57432 );
nor ( n58400 , n11799 , n58228 );
and ( n58401 , n58399 , n58400 );
xor ( n58402 , n58399 , n58400 );
xor ( n58403 , n57211 , n57430 );
nor ( n58404 , n11050 , n58228 );
and ( n58405 , n58403 , n58404 );
xor ( n58406 , n58403 , n58404 );
xor ( n58407 , n57215 , n57428 );
nor ( n58408 , n10321 , n58228 );
and ( n58409 , n58407 , n58408 );
xor ( n58410 , n58407 , n58408 );
xor ( n58411 , n57219 , n57426 );
nor ( n58412 , n9429 , n58228 );
and ( n58413 , n58411 , n58412 );
xor ( n58414 , n58411 , n58412 );
xor ( n58415 , n57223 , n57424 );
nor ( n58416 , n8949 , n58228 );
and ( n58417 , n58415 , n58416 );
xor ( n58418 , n58415 , n58416 );
xor ( n58419 , n57227 , n57422 );
nor ( n58420 , n9437 , n58228 );
and ( n58421 , n58419 , n58420 );
xor ( n58422 , n58419 , n58420 );
xor ( n58423 , n57231 , n57420 );
nor ( n58424 , n9446 , n58228 );
and ( n58425 , n58423 , n58424 );
xor ( n58426 , n58423 , n58424 );
xor ( n58427 , n57235 , n57418 );
nor ( n58428 , n9455 , n58228 );
and ( n58429 , n58427 , n58428 );
xor ( n58430 , n58427 , n58428 );
xor ( n58431 , n57239 , n57416 );
nor ( n58432 , n9464 , n58228 );
and ( n58433 , n58431 , n58432 );
xor ( n58434 , n58431 , n58432 );
xor ( n58435 , n57243 , n57414 );
nor ( n58436 , n9473 , n58228 );
and ( n58437 , n58435 , n58436 );
xor ( n58438 , n58435 , n58436 );
xor ( n58439 , n57247 , n57412 );
nor ( n58440 , n9482 , n58228 );
and ( n58441 , n58439 , n58440 );
xor ( n58442 , n58439 , n58440 );
xor ( n58443 , n57251 , n57410 );
nor ( n58444 , n9491 , n58228 );
and ( n58445 , n58443 , n58444 );
xor ( n58446 , n58443 , n58444 );
xor ( n58447 , n57255 , n57408 );
nor ( n58448 , n9500 , n58228 );
and ( n58449 , n58447 , n58448 );
xor ( n58450 , n58447 , n58448 );
xor ( n58451 , n57259 , n57406 );
nor ( n58452 , n9509 , n58228 );
and ( n58453 , n58451 , n58452 );
xor ( n58454 , n58451 , n58452 );
xor ( n58455 , n57263 , n57404 );
nor ( n58456 , n9518 , n58228 );
and ( n58457 , n58455 , n58456 );
xor ( n58458 , n58455 , n58456 );
xor ( n58459 , n57267 , n57402 );
nor ( n58460 , n9527 , n58228 );
and ( n58461 , n58459 , n58460 );
xor ( n58462 , n58459 , n58460 );
xor ( n58463 , n57271 , n57400 );
nor ( n58464 , n9536 , n58228 );
and ( n58465 , n58463 , n58464 );
xor ( n58466 , n58463 , n58464 );
xor ( n58467 , n57275 , n57398 );
nor ( n58468 , n9545 , n58228 );
and ( n58469 , n58467 , n58468 );
xor ( n58470 , n58467 , n58468 );
xor ( n58471 , n57279 , n57396 );
nor ( n58472 , n9554 , n58228 );
and ( n58473 , n58471 , n58472 );
xor ( n58474 , n58471 , n58472 );
xor ( n58475 , n57283 , n57394 );
nor ( n58476 , n9563 , n58228 );
and ( n58477 , n58475 , n58476 );
xor ( n58478 , n58475 , n58476 );
xor ( n58479 , n57287 , n57392 );
nor ( n58480 , n9572 , n58228 );
and ( n58481 , n58479 , n58480 );
xor ( n58482 , n58479 , n58480 );
xor ( n58483 , n57291 , n57390 );
nor ( n58484 , n9581 , n58228 );
and ( n58485 , n58483 , n58484 );
xor ( n58486 , n58483 , n58484 );
xor ( n58487 , n57295 , n57388 );
nor ( n58488 , n9590 , n58228 );
and ( n58489 , n58487 , n58488 );
xor ( n58490 , n58487 , n58488 );
xor ( n58491 , n57299 , n57386 );
nor ( n58492 , n9599 , n58228 );
and ( n58493 , n58491 , n58492 );
xor ( n58494 , n58491 , n58492 );
xor ( n58495 , n57303 , n57384 );
nor ( n58496 , n9608 , n58228 );
and ( n58497 , n58495 , n58496 );
xor ( n58498 , n58495 , n58496 );
xor ( n58499 , n57307 , n57382 );
nor ( n58500 , n9617 , n58228 );
and ( n58501 , n58499 , n58500 );
xor ( n58502 , n58499 , n58500 );
xor ( n58503 , n57311 , n57380 );
nor ( n58504 , n9626 , n58228 );
and ( n58505 , n58503 , n58504 );
xor ( n58506 , n58503 , n58504 );
xor ( n58507 , n57315 , n57378 );
nor ( n58508 , n9635 , n58228 );
and ( n58509 , n58507 , n58508 );
xor ( n58510 , n58507 , n58508 );
xor ( n58511 , n57319 , n57376 );
nor ( n58512 , n9644 , n58228 );
and ( n58513 , n58511 , n58512 );
xor ( n58514 , n58511 , n58512 );
xor ( n58515 , n57323 , n57374 );
nor ( n58516 , n9653 , n58228 );
and ( n58517 , n58515 , n58516 );
xor ( n58518 , n58515 , n58516 );
xor ( n58519 , n57327 , n57372 );
nor ( n58520 , n9662 , n58228 );
and ( n58521 , n58519 , n58520 );
xor ( n58522 , n58519 , n58520 );
xor ( n58523 , n57331 , n57370 );
nor ( n58524 , n9671 , n58228 );
and ( n58525 , n58523 , n58524 );
xor ( n58526 , n58523 , n58524 );
xor ( n58527 , n57335 , n57368 );
nor ( n58528 , n9680 , n58228 );
and ( n58529 , n58527 , n58528 );
xor ( n58530 , n58527 , n58528 );
xor ( n58531 , n57339 , n57366 );
nor ( n58532 , n9689 , n58228 );
and ( n58533 , n58531 , n58532 );
xor ( n58534 , n58531 , n58532 );
xor ( n58535 , n57343 , n57364 );
nor ( n58536 , n9698 , n58228 );
and ( n58537 , n58535 , n58536 );
xor ( n58538 , n58535 , n58536 );
xor ( n58539 , n57347 , n57362 );
nor ( n58540 , n9707 , n58228 );
and ( n58541 , n58539 , n58540 );
xor ( n58542 , n58539 , n58540 );
xor ( n58543 , n57351 , n57360 );
nor ( n58544 , n9716 , n58228 );
and ( n58545 , n58543 , n58544 );
xor ( n58546 , n58543 , n58544 );
xor ( n58547 , n57355 , n57358 );
nor ( n58548 , n9725 , n58228 );
and ( n58549 , n58547 , n58548 );
xor ( n58550 , n58547 , n58548 );
xor ( n58551 , n57356 , n57357 );
nor ( n58552 , n9734 , n58228 );
and ( n58553 , n58551 , n58552 );
xor ( n58554 , n58551 , n58552 );
nor ( n58555 , n9752 , n57033 );
nor ( n58556 , n9743 , n58228 );
and ( n58557 , n58555 , n58556 );
and ( n58558 , n58554 , n58557 );
or ( n58559 , n58553 , n58558 );
and ( n58560 , n58550 , n58559 );
or ( n58561 , n58549 , n58560 );
and ( n58562 , n58546 , n58561 );
or ( n58563 , n58545 , n58562 );
and ( n58564 , n58542 , n58563 );
or ( n58565 , n58541 , n58564 );
and ( n58566 , n58538 , n58565 );
or ( n58567 , n58537 , n58566 );
and ( n58568 , n58534 , n58567 );
or ( n58569 , n58533 , n58568 );
and ( n58570 , n58530 , n58569 );
or ( n58571 , n58529 , n58570 );
and ( n58572 , n58526 , n58571 );
or ( n58573 , n58525 , n58572 );
and ( n58574 , n58522 , n58573 );
or ( n58575 , n58521 , n58574 );
and ( n58576 , n58518 , n58575 );
or ( n58577 , n58517 , n58576 );
and ( n58578 , n58514 , n58577 );
or ( n58579 , n58513 , n58578 );
and ( n58580 , n58510 , n58579 );
or ( n58581 , n58509 , n58580 );
and ( n58582 , n58506 , n58581 );
or ( n58583 , n58505 , n58582 );
and ( n58584 , n58502 , n58583 );
or ( n58585 , n58501 , n58584 );
and ( n58586 , n58498 , n58585 );
or ( n58587 , n58497 , n58586 );
and ( n58588 , n58494 , n58587 );
or ( n58589 , n58493 , n58588 );
and ( n58590 , n58490 , n58589 );
or ( n58591 , n58489 , n58590 );
and ( n58592 , n58486 , n58591 );
or ( n58593 , n58485 , n58592 );
and ( n58594 , n58482 , n58593 );
or ( n58595 , n58481 , n58594 );
and ( n58596 , n58478 , n58595 );
or ( n58597 , n58477 , n58596 );
and ( n58598 , n58474 , n58597 );
or ( n58599 , n58473 , n58598 );
and ( n58600 , n58470 , n58599 );
or ( n58601 , n58469 , n58600 );
and ( n58602 , n58466 , n58601 );
or ( n58603 , n58465 , n58602 );
and ( n58604 , n58462 , n58603 );
or ( n58605 , n58461 , n58604 );
and ( n58606 , n58458 , n58605 );
or ( n58607 , n58457 , n58606 );
and ( n58608 , n58454 , n58607 );
or ( n58609 , n58453 , n58608 );
and ( n58610 , n58450 , n58609 );
or ( n58611 , n58449 , n58610 );
and ( n58612 , n58446 , n58611 );
or ( n58613 , n58445 , n58612 );
and ( n58614 , n58442 , n58613 );
or ( n58615 , n58441 , n58614 );
and ( n58616 , n58438 , n58615 );
or ( n58617 , n58437 , n58616 );
and ( n58618 , n58434 , n58617 );
or ( n58619 , n58433 , n58618 );
and ( n58620 , n58430 , n58619 );
or ( n58621 , n58429 , n58620 );
and ( n58622 , n58426 , n58621 );
or ( n58623 , n58425 , n58622 );
and ( n58624 , n58422 , n58623 );
or ( n58625 , n58421 , n58624 );
and ( n58626 , n58418 , n58625 );
or ( n58627 , n58417 , n58626 );
and ( n58628 , n58414 , n58627 );
or ( n58629 , n58413 , n58628 );
and ( n58630 , n58410 , n58629 );
or ( n58631 , n58409 , n58630 );
and ( n58632 , n58406 , n58631 );
or ( n58633 , n58405 , n58632 );
and ( n58634 , n58402 , n58633 );
or ( n58635 , n58401 , n58634 );
and ( n58636 , n58398 , n58635 );
or ( n58637 , n58397 , n58636 );
and ( n58638 , n58394 , n58637 );
or ( n58639 , n58393 , n58638 );
and ( n58640 , n58390 , n58639 );
or ( n58641 , n58389 , n58640 );
and ( n58642 , n58386 , n58641 );
or ( n58643 , n58385 , n58642 );
and ( n58644 , n58382 , n58643 );
or ( n58645 , n58381 , n58644 );
and ( n58646 , n58378 , n58645 );
or ( n58647 , n58377 , n58646 );
and ( n58648 , n58374 , n58647 );
or ( n58649 , n58373 , n58648 );
and ( n58650 , n58370 , n58649 );
or ( n58651 , n58369 , n58650 );
and ( n58652 , n58366 , n58651 );
or ( n58653 , n58365 , n58652 );
and ( n58654 , n58362 , n58653 );
or ( n58655 , n58361 , n58654 );
and ( n58656 , n58358 , n58655 );
or ( n58657 , n58357 , n58656 );
and ( n58658 , n58354 , n58657 );
or ( n58659 , n58353 , n58658 );
and ( n58660 , n58350 , n58659 );
or ( n58661 , n58349 , n58660 );
and ( n58662 , n58346 , n58661 );
or ( n58663 , n58345 , n58662 );
and ( n58664 , n58342 , n58663 );
or ( n58665 , n58341 , n58664 );
and ( n58666 , n58338 , n58665 );
or ( n58667 , n58337 , n58666 );
and ( n58668 , n58334 , n58667 );
or ( n58669 , n58333 , n58668 );
and ( n58670 , n58330 , n58669 );
or ( n58671 , n58329 , n58670 );
and ( n58672 , n58326 , n58671 );
or ( n58673 , n58325 , n58672 );
and ( n58674 , n58322 , n58673 );
or ( n58675 , n58321 , n58674 );
and ( n58676 , n58318 , n58675 );
or ( n58677 , n58317 , n58676 );
and ( n58678 , n58314 , n58677 );
or ( n58679 , n58313 , n58678 );
and ( n58680 , n58310 , n58679 );
or ( n58681 , n58309 , n58680 );
and ( n58682 , n58306 , n58681 );
or ( n58683 , n58305 , n58682 );
and ( n58684 , n58302 , n58683 );
or ( n58685 , n58301 , n58684 );
and ( n58686 , n58298 , n58685 );
or ( n58687 , n58297 , n58686 );
and ( n58688 , n58294 , n58687 );
or ( n58689 , n58293 , n58688 );
and ( n58690 , n58290 , n58689 );
or ( n58691 , n58289 , n58690 );
and ( n58692 , n58286 , n58691 );
or ( n58693 , n58285 , n58692 );
and ( n58694 , n58282 , n58693 );
or ( n58695 , n58281 , n58694 );
and ( n58696 , n58278 , n58695 );
or ( n58697 , n58277 , n58696 );
and ( n58698 , n58274 , n58697 );
or ( n58699 , n58273 , n58698 );
and ( n58700 , n58270 , n58699 );
or ( n58701 , n58269 , n58700 );
and ( n58702 , n58266 , n58701 );
or ( n58703 , n58265 , n58702 );
and ( n58704 , n58262 , n58703 );
or ( n58705 , n58261 , n58704 );
and ( n58706 , n58258 , n58705 );
or ( n58707 , n58257 , n58706 );
and ( n58708 , n58254 , n58707 );
or ( n58709 , n58253 , n58708 );
and ( n58710 , n58250 , n58709 );
or ( n58711 , n58249 , n58710 );
and ( n58712 , n58246 , n58711 );
or ( n58713 , n58245 , n58712 );
and ( n58714 , n58242 , n58713 );
or ( n58715 , n58241 , n58714 );
and ( n58716 , n58238 , n58715 );
or ( n58717 , n58237 , n58716 );
and ( n58718 , n58234 , n58717 );
or ( n58719 , n58233 , n58718 );
xor ( n58720 , n58230 , n58719 );
and ( n58721 , n33403 , n3299 );
nor ( n58722 , n3300 , n58721 );
nor ( n58723 , n3570 , n32231 );
xor ( n58724 , n58722 , n58723 );
and ( n58725 , n57521 , n57522 );
and ( n58726 , n57523 , n57526 );
or ( n58727 , n58725 , n58726 );
xor ( n58728 , n58724 , n58727 );
nor ( n58729 , n3853 , n31083 );
xor ( n58730 , n58728 , n58729 );
and ( n58731 , n57527 , n57528 );
and ( n58732 , n57529 , n57532 );
or ( n58733 , n58731 , n58732 );
xor ( n58734 , n58730 , n58733 );
nor ( n58735 , n4151 , n29948 );
xor ( n58736 , n58734 , n58735 );
and ( n58737 , n57533 , n57534 );
and ( n58738 , n57535 , n57538 );
or ( n58739 , n58737 , n58738 );
xor ( n58740 , n58736 , n58739 );
nor ( n58741 , n4458 , n28833 );
xor ( n58742 , n58740 , n58741 );
and ( n58743 , n57539 , n57540 );
and ( n58744 , n57541 , n57544 );
or ( n58745 , n58743 , n58744 );
xor ( n58746 , n58742 , n58745 );
nor ( n58747 , n4786 , n27737 );
xor ( n58748 , n58746 , n58747 );
and ( n58749 , n57545 , n57546 );
and ( n58750 , n57547 , n57550 );
or ( n58751 , n58749 , n58750 );
xor ( n58752 , n58748 , n58751 );
nor ( n58753 , n5126 , n26660 );
xor ( n58754 , n58752 , n58753 );
and ( n58755 , n57551 , n57552 );
and ( n58756 , n57553 , n57556 );
or ( n58757 , n58755 , n58756 );
xor ( n58758 , n58754 , n58757 );
nor ( n58759 , n5477 , n25600 );
xor ( n58760 , n58758 , n58759 );
and ( n58761 , n57557 , n57558 );
and ( n58762 , n57559 , n57562 );
or ( n58763 , n58761 , n58762 );
xor ( n58764 , n58760 , n58763 );
nor ( n58765 , n5838 , n24564 );
xor ( n58766 , n58764 , n58765 );
and ( n58767 , n57563 , n57564 );
and ( n58768 , n57565 , n57568 );
or ( n58769 , n58767 , n58768 );
xor ( n58770 , n58766 , n58769 );
nor ( n58771 , n6212 , n23541 );
xor ( n58772 , n58770 , n58771 );
and ( n58773 , n57569 , n57570 );
and ( n58774 , n57571 , n57574 );
or ( n58775 , n58773 , n58774 );
xor ( n58776 , n58772 , n58775 );
nor ( n58777 , n6596 , n22541 );
xor ( n58778 , n58776 , n58777 );
and ( n58779 , n57575 , n57576 );
and ( n58780 , n57577 , n57580 );
or ( n58781 , n58779 , n58780 );
xor ( n58782 , n58778 , n58781 );
nor ( n58783 , n6997 , n21562 );
xor ( n58784 , n58782 , n58783 );
and ( n58785 , n57581 , n57582 );
and ( n58786 , n57583 , n57586 );
or ( n58787 , n58785 , n58786 );
xor ( n58788 , n58784 , n58787 );
nor ( n58789 , n7413 , n20601 );
xor ( n58790 , n58788 , n58789 );
and ( n58791 , n57587 , n57588 );
and ( n58792 , n57589 , n57592 );
or ( n58793 , n58791 , n58792 );
xor ( n58794 , n58790 , n58793 );
nor ( n58795 , n7841 , n19657 );
xor ( n58796 , n58794 , n58795 );
and ( n58797 , n57593 , n57594 );
and ( n58798 , n57595 , n57598 );
or ( n58799 , n58797 , n58798 );
xor ( n58800 , n58796 , n58799 );
nor ( n58801 , n8281 , n18734 );
xor ( n58802 , n58800 , n58801 );
and ( n58803 , n57599 , n57600 );
and ( n58804 , n57601 , n57604 );
or ( n58805 , n58803 , n58804 );
xor ( n58806 , n58802 , n58805 );
nor ( n58807 , n8737 , n17828 );
xor ( n58808 , n58806 , n58807 );
and ( n58809 , n57605 , n57606 );
and ( n58810 , n57607 , n57610 );
or ( n58811 , n58809 , n58810 );
xor ( n58812 , n58808 , n58811 );
nor ( n58813 , n9420 , n16943 );
xor ( n58814 , n58812 , n58813 );
and ( n58815 , n57611 , n57612 );
and ( n58816 , n57613 , n57616 );
or ( n58817 , n58815 , n58816 );
xor ( n58818 , n58814 , n58817 );
nor ( n58819 , n10312 , n16077 );
xor ( n58820 , n58818 , n58819 );
and ( n58821 , n57617 , n57618 );
and ( n58822 , n57619 , n57622 );
or ( n58823 , n58821 , n58822 );
xor ( n58824 , n58820 , n58823 );
nor ( n58825 , n11041 , n15230 );
xor ( n58826 , n58824 , n58825 );
and ( n58827 , n57623 , n57624 );
and ( n58828 , n57625 , n57628 );
or ( n58829 , n58827 , n58828 );
xor ( n58830 , n58826 , n58829 );
nor ( n58831 , n11790 , n14403 );
xor ( n58832 , n58830 , n58831 );
and ( n58833 , n57629 , n57630 );
and ( n58834 , n57631 , n57634 );
or ( n58835 , n58833 , n58834 );
xor ( n58836 , n58832 , n58835 );
nor ( n58837 , n12555 , n13599 );
xor ( n58838 , n58836 , n58837 );
and ( n58839 , n57635 , n57636 );
and ( n58840 , n57637 , n57640 );
or ( n58841 , n58839 , n58840 );
xor ( n58842 , n58838 , n58841 );
nor ( n58843 , n13340 , n12808 );
xor ( n58844 , n58842 , n58843 );
and ( n58845 , n57641 , n57642 );
and ( n58846 , n57643 , n57646 );
or ( n58847 , n58845 , n58846 );
xor ( n58848 , n58844 , n58847 );
nor ( n58849 , n14138 , n12037 );
xor ( n58850 , n58848 , n58849 );
and ( n58851 , n57647 , n57648 );
and ( n58852 , n57649 , n57652 );
or ( n58853 , n58851 , n58852 );
xor ( n58854 , n58850 , n58853 );
nor ( n58855 , n14959 , n11282 );
xor ( n58856 , n58854 , n58855 );
and ( n58857 , n57653 , n57654 );
and ( n58858 , n57655 , n57658 );
or ( n58859 , n58857 , n58858 );
xor ( n58860 , n58856 , n58859 );
nor ( n58861 , n15800 , n10547 );
xor ( n58862 , n58860 , n58861 );
and ( n58863 , n57659 , n57660 );
and ( n58864 , n57661 , n57664 );
or ( n58865 , n58863 , n58864 );
xor ( n58866 , n58862 , n58865 );
nor ( n58867 , n16660 , n9829 );
xor ( n58868 , n58866 , n58867 );
and ( n58869 , n57665 , n57666 );
and ( n58870 , n57667 , n57670 );
or ( n58871 , n58869 , n58870 );
xor ( n58872 , n58868 , n58871 );
nor ( n58873 , n17539 , n8955 );
xor ( n58874 , n58872 , n58873 );
and ( n58875 , n57671 , n57672 );
and ( n58876 , n57673 , n57676 );
or ( n58877 , n58875 , n58876 );
xor ( n58878 , n58874 , n58877 );
nor ( n58879 , n18439 , n603 );
xor ( n58880 , n58878 , n58879 );
and ( n58881 , n57677 , n57678 );
and ( n58882 , n57679 , n57682 );
or ( n58883 , n58881 , n58882 );
xor ( n58884 , n58880 , n58883 );
nor ( n58885 , n19356 , n652 );
xor ( n58886 , n58884 , n58885 );
and ( n58887 , n57683 , n57684 );
and ( n58888 , n57685 , n57688 );
or ( n58889 , n58887 , n58888 );
xor ( n58890 , n58886 , n58889 );
nor ( n58891 , n20294 , n624 );
xor ( n58892 , n58890 , n58891 );
and ( n58893 , n57689 , n57690 );
and ( n58894 , n57691 , n57694 );
or ( n58895 , n58893 , n58894 );
xor ( n58896 , n58892 , n58895 );
nor ( n58897 , n21249 , n648 );
xor ( n58898 , n58896 , n58897 );
and ( n58899 , n57695 , n57696 );
and ( n58900 , n57697 , n57700 );
or ( n58901 , n58899 , n58900 );
xor ( n58902 , n58898 , n58901 );
nor ( n58903 , n22222 , n686 );
xor ( n58904 , n58902 , n58903 );
and ( n58905 , n57701 , n57702 );
and ( n58906 , n57703 , n57706 );
or ( n58907 , n58905 , n58906 );
xor ( n58908 , n58904 , n58907 );
nor ( n58909 , n23216 , n735 );
xor ( n58910 , n58908 , n58909 );
and ( n58911 , n57707 , n57708 );
and ( n58912 , n57709 , n57712 );
or ( n58913 , n58911 , n58912 );
xor ( n58914 , n58910 , n58913 );
nor ( n58915 , n24233 , n798 );
xor ( n58916 , n58914 , n58915 );
and ( n58917 , n57713 , n57714 );
and ( n58918 , n57715 , n57718 );
or ( n58919 , n58917 , n58918 );
xor ( n58920 , n58916 , n58919 );
nor ( n58921 , n25263 , n870 );
xor ( n58922 , n58920 , n58921 );
and ( n58923 , n57719 , n57720 );
and ( n58924 , n57721 , n57724 );
or ( n58925 , n58923 , n58924 );
xor ( n58926 , n58922 , n58925 );
nor ( n58927 , n26317 , n960 );
xor ( n58928 , n58926 , n58927 );
and ( n58929 , n57725 , n57726 );
and ( n58930 , n57727 , n57730 );
or ( n58931 , n58929 , n58930 );
xor ( n58932 , n58928 , n58931 );
nor ( n58933 , n27388 , n1064 );
xor ( n58934 , n58932 , n58933 );
and ( n58935 , n57731 , n57732 );
and ( n58936 , n57733 , n57736 );
or ( n58937 , n58935 , n58936 );
xor ( n58938 , n58934 , n58937 );
nor ( n58939 , n28478 , n1178 );
xor ( n58940 , n58938 , n58939 );
and ( n58941 , n57737 , n57738 );
and ( n58942 , n57739 , n57742 );
or ( n58943 , n58941 , n58942 );
xor ( n58944 , n58940 , n58943 );
nor ( n58945 , n29587 , n1305 );
xor ( n58946 , n58944 , n58945 );
and ( n58947 , n57743 , n57744 );
and ( n58948 , n57745 , n57748 );
or ( n58949 , n58947 , n58948 );
xor ( n58950 , n58946 , n58949 );
nor ( n58951 , n30716 , n1447 );
xor ( n58952 , n58950 , n58951 );
and ( n58953 , n57749 , n57750 );
and ( n58954 , n57751 , n57754 );
or ( n58955 , n58953 , n58954 );
xor ( n58956 , n58952 , n58955 );
nor ( n58957 , n31858 , n1600 );
xor ( n58958 , n58956 , n58957 );
and ( n58959 , n57755 , n57756 );
and ( n58960 , n57757 , n57760 );
or ( n58961 , n58959 , n58960 );
xor ( n58962 , n58958 , n58961 );
nor ( n58963 , n33024 , n1768 );
xor ( n58964 , n58962 , n58963 );
and ( n58965 , n57761 , n57762 );
and ( n58966 , n57763 , n57766 );
or ( n58967 , n58965 , n58966 );
xor ( n58968 , n58964 , n58967 );
nor ( n58969 , n34215 , n1947 );
xor ( n58970 , n58968 , n58969 );
and ( n58971 , n57767 , n57768 );
and ( n58972 , n57769 , n57772 );
or ( n58973 , n58971 , n58972 );
xor ( n58974 , n58970 , n58973 );
nor ( n58975 , n35410 , n2139 );
xor ( n58976 , n58974 , n58975 );
and ( n58977 , n57773 , n57774 );
and ( n58978 , n57775 , n57778 );
or ( n58979 , n58977 , n58978 );
xor ( n58980 , n58976 , n58979 );
nor ( n58981 , n36611 , n2345 );
xor ( n58982 , n58980 , n58981 );
and ( n58983 , n57779 , n57780 );
and ( n58984 , n57781 , n57784 );
or ( n58985 , n58983 , n58984 );
xor ( n58986 , n58982 , n58985 );
nor ( n58987 , n37816 , n2568 );
xor ( n58988 , n58986 , n58987 );
and ( n58989 , n57785 , n57786 );
and ( n58990 , n57787 , n57790 );
or ( n58991 , n58989 , n58990 );
xor ( n58992 , n58988 , n58991 );
nor ( n58993 , n39018 , n2799 );
xor ( n58994 , n58992 , n58993 );
and ( n58995 , n57791 , n57792 );
and ( n58996 , n57793 , n57796 );
or ( n58997 , n58995 , n58996 );
xor ( n58998 , n58994 , n58997 );
nor ( n58999 , n40223 , n3045 );
xor ( n59000 , n58998 , n58999 );
and ( n59001 , n57797 , n57798 );
and ( n59002 , n57799 , n57802 );
or ( n59003 , n59001 , n59002 );
xor ( n59004 , n59000 , n59003 );
nor ( n59005 , n41428 , n3302 );
xor ( n59006 , n59004 , n59005 );
and ( n59007 , n57803 , n57804 );
and ( n59008 , n57805 , n57808 );
or ( n59009 , n59007 , n59008 );
xor ( n59010 , n59006 , n59009 );
nor ( n59011 , n42632 , n3572 );
xor ( n59012 , n59010 , n59011 );
and ( n59013 , n57809 , n57810 );
and ( n59014 , n57811 , n57814 );
or ( n59015 , n59013 , n59014 );
xor ( n59016 , n59012 , n59015 );
nor ( n59017 , n43834 , n3855 );
xor ( n59018 , n59016 , n59017 );
and ( n59019 , n57815 , n57816 );
and ( n59020 , n57817 , n57820 );
or ( n59021 , n59019 , n59020 );
xor ( n59022 , n59018 , n59021 );
nor ( n59023 , n45038 , n4153 );
xor ( n59024 , n59022 , n59023 );
and ( n59025 , n57821 , n57822 );
and ( n59026 , n57823 , n57826 );
or ( n59027 , n59025 , n59026 );
xor ( n59028 , n59024 , n59027 );
nor ( n59029 , n46239 , n4460 );
xor ( n59030 , n59028 , n59029 );
and ( n59031 , n57827 , n57828 );
and ( n59032 , n57829 , n57832 );
or ( n59033 , n59031 , n59032 );
xor ( n59034 , n59030 , n59033 );
nor ( n59035 , n47440 , n4788 );
xor ( n59036 , n59034 , n59035 );
and ( n59037 , n57833 , n57834 );
and ( n59038 , n57835 , n57838 );
or ( n59039 , n59037 , n59038 );
xor ( n59040 , n59036 , n59039 );
nor ( n59041 , n48641 , n5128 );
xor ( n59042 , n59040 , n59041 );
and ( n59043 , n57839 , n57840 );
and ( n59044 , n57841 , n57844 );
or ( n59045 , n59043 , n59044 );
xor ( n59046 , n59042 , n59045 );
nor ( n59047 , n49841 , n5479 );
xor ( n59048 , n59046 , n59047 );
and ( n59049 , n57845 , n57846 );
and ( n59050 , n57847 , n57850 );
or ( n59051 , n59049 , n59050 );
xor ( n59052 , n59048 , n59051 );
nor ( n59053 , n51040 , n5840 );
xor ( n59054 , n59052 , n59053 );
and ( n59055 , n57851 , n57852 );
and ( n59056 , n57853 , n57856 );
or ( n59057 , n59055 , n59056 );
xor ( n59058 , n59054 , n59057 );
nor ( n59059 , n52238 , n6214 );
xor ( n59060 , n59058 , n59059 );
and ( n59061 , n57857 , n57858 );
and ( n59062 , n57859 , n57862 );
or ( n59063 , n59061 , n59062 );
xor ( n59064 , n59060 , n59063 );
nor ( n59065 , n53432 , n6598 );
xor ( n59066 , n59064 , n59065 );
and ( n59067 , n57863 , n57864 );
and ( n59068 , n57865 , n57868 );
or ( n59069 , n59067 , n59068 );
xor ( n59070 , n59066 , n59069 );
nor ( n59071 , n54629 , n6999 );
xor ( n59072 , n59070 , n59071 );
and ( n59073 , n57869 , n57870 );
and ( n59074 , n57871 , n57874 );
or ( n59075 , n59073 , n59074 );
xor ( n59076 , n59072 , n59075 );
nor ( n59077 , n55826 , n7415 );
xor ( n59078 , n59076 , n59077 );
and ( n59079 , n57875 , n57876 );
and ( n59080 , n57877 , n57880 );
or ( n59081 , n59079 , n59080 );
xor ( n59082 , n59078 , n59081 );
nor ( n59083 , n57022 , n7843 );
xor ( n59084 , n59082 , n59083 );
and ( n59085 , n57881 , n57882 );
and ( n59086 , n57883 , n57886 );
or ( n59087 , n59085 , n59086 );
xor ( n59088 , n59084 , n59087 );
nor ( n59089 , n58217 , n8283 );
xor ( n59090 , n59088 , n59089 );
and ( n59091 , n57887 , n57888 );
and ( n59092 , n57889 , n57892 );
or ( n59093 , n59091 , n59092 );
xor ( n59094 , n59090 , n59093 );
and ( n59095 , n57905 , n57909 );
and ( n59096 , n57909 , n58203 );
and ( n59097 , n57905 , n58203 );
or ( n59098 , n59095 , n59096 , n59097 );
and ( n59099 , n33774 , n3271 );
not ( n59100 , n3271 );
nor ( n59101 , n59099 , n59100 );
xor ( n59102 , n59098 , n59101 );
and ( n59103 , n57918 , n57922 );
and ( n59104 , n57922 , n57990 );
and ( n59105 , n57918 , n57990 );
or ( n59106 , n59103 , n59104 , n59105 );
and ( n59107 , n57914 , n57991 );
and ( n59108 , n57991 , n58202 );
and ( n59109 , n57914 , n58202 );
or ( n59110 , n59107 , n59108 , n59109 );
xor ( n59111 , n59106 , n59110 );
and ( n59112 , n57993 , n58113 );
and ( n59113 , n58113 , n58201 );
and ( n59114 , n57993 , n58201 );
or ( n59115 , n59112 , n59113 , n59114 );
and ( n59116 , n57927 , n57931 );
and ( n59117 , n57931 , n57989 );
and ( n59118 , n57927 , n57989 );
or ( n59119 , n59116 , n59117 , n59118 );
and ( n59120 , n57997 , n58001 );
and ( n59121 , n58001 , n58112 );
and ( n59122 , n57997 , n58112 );
or ( n59123 , n59120 , n59121 , n59122 );
xor ( n59124 , n59119 , n59123 );
and ( n59125 , n57958 , n57962 );
and ( n59126 , n57962 , n57968 );
and ( n59127 , n57958 , n57968 );
or ( n59128 , n59125 , n59126 , n59127 );
and ( n59129 , n57936 , n57940 );
and ( n59130 , n57940 , n57988 );
and ( n59131 , n57936 , n57988 );
or ( n59132 , n59129 , n59130 , n59131 );
xor ( n59133 , n59128 , n59132 );
and ( n59134 , n57945 , n57949 );
and ( n59135 , n57949 , n57987 );
and ( n59136 , n57945 , n57987 );
or ( n59137 , n59134 , n59135 , n59136 );
and ( n59138 , n58010 , n58035 );
and ( n59139 , n58035 , n58073 );
and ( n59140 , n58010 , n58073 );
or ( n59141 , n59138 , n59139 , n59140 );
xor ( n59142 , n59137 , n59141 );
and ( n59143 , n57954 , n57969 );
and ( n59144 , n57969 , n57986 );
and ( n59145 , n57954 , n57986 );
or ( n59146 , n59143 , n59144 , n59145 );
and ( n59147 , n58014 , n58018 );
and ( n59148 , n58018 , n58034 );
and ( n59149 , n58014 , n58034 );
or ( n59150 , n59147 , n59148 , n59149 );
xor ( n59151 , n59146 , n59150 );
and ( n59152 , n57974 , n57979 );
and ( n59153 , n57979 , n57985 );
and ( n59154 , n57974 , n57985 );
or ( n59155 , n59152 , n59153 , n59154 );
and ( n59156 , n57964 , n57965 );
and ( n59157 , n57965 , n57967 );
and ( n59158 , n57964 , n57967 );
or ( n59159 , n59156 , n59157 , n59158 );
and ( n59160 , n57975 , n57976 );
and ( n59161 , n57976 , n57978 );
and ( n59162 , n57975 , n57978 );
or ( n59163 , n59160 , n59161 , n59162 );
xor ( n59164 , n59159 , n59163 );
and ( n59165 , n30695 , n4102 );
and ( n59166 , n31836 , n3749 );
xor ( n59167 , n59165 , n59166 );
and ( n59168 , n32649 , n3495 );
xor ( n59169 , n59167 , n59168 );
xor ( n59170 , n59164 , n59169 );
xor ( n59171 , n59155 , n59170 );
and ( n59172 , n57981 , n57982 );
and ( n59173 , n57982 , n57984 );
and ( n59174 , n57981 , n57984 );
or ( n59175 , n59172 , n59173 , n59174 );
and ( n59176 , n27361 , n5103 );
and ( n59177 , n28456 , n4730 );
xor ( n59178 , n59176 , n59177 );
and ( n59179 , n29559 , n4403 );
xor ( n59180 , n59178 , n59179 );
xor ( n59181 , n59175 , n59180 );
and ( n59182 , n24214 , n6132 );
and ( n59183 , n25243 , n5765 );
xor ( n59184 , n59182 , n59183 );
and ( n59185 , n26296 , n5408 );
xor ( n59186 , n59184 , n59185 );
xor ( n59187 , n59181 , n59186 );
xor ( n59188 , n59171 , n59187 );
xor ( n59189 , n59151 , n59188 );
xor ( n59190 , n59142 , n59189 );
xor ( n59191 , n59133 , n59190 );
xor ( n59192 , n59124 , n59191 );
xor ( n59193 , n59115 , n59192 );
and ( n59194 , n58125 , n58200 );
and ( n59195 , n58129 , n58130 );
and ( n59196 , n58130 , n58199 );
and ( n59197 , n58129 , n58199 );
or ( n59198 , n59195 , n59196 , n59197 );
and ( n59199 , n58006 , n58074 );
and ( n59200 , n58074 , n58111 );
and ( n59201 , n58006 , n58111 );
or ( n59202 , n59199 , n59200 , n59201 );
xor ( n59203 , n59198 , n59202 );
and ( n59204 , n58079 , n58083 );
and ( n59205 , n58083 , n58110 );
and ( n59206 , n58079 , n58110 );
or ( n59207 , n59204 , n59205 , n59206 );
and ( n59208 , n58040 , n58056 );
and ( n59209 , n58056 , n58072 );
and ( n59210 , n58040 , n58072 );
or ( n59211 , n59208 , n59209 , n59210 );
and ( n59212 , n58023 , n58027 );
and ( n59213 , n58027 , n58033 );
and ( n59214 , n58023 , n58033 );
or ( n59215 , n59212 , n59213 , n59214 );
and ( n59216 , n58044 , n58049 );
and ( n59217 , n58049 , n58055 );
and ( n59218 , n58044 , n58055 );
or ( n59219 , n59216 , n59217 , n59218 );
xor ( n59220 , n59215 , n59219 );
and ( n59221 , n58029 , n58030 );
and ( n59222 , n58030 , n58032 );
and ( n59223 , n58029 , n58032 );
or ( n59224 , n59221 , n59222 , n59223 );
and ( n59225 , n58045 , n58046 );
and ( n59226 , n58046 , n58048 );
and ( n59227 , n58045 , n58048 );
or ( n59228 , n59225 , n59226 , n59227 );
xor ( n59229 , n59224 , n59228 );
and ( n59230 , n21216 , n7310 );
and ( n59231 , n22186 , n6971 );
xor ( n59232 , n59230 , n59231 );
and ( n59233 , n22892 , n6504 );
xor ( n59234 , n59232 , n59233 );
xor ( n59235 , n59229 , n59234 );
xor ( n59236 , n59220 , n59235 );
xor ( n59237 , n59211 , n59236 );
and ( n59238 , n58061 , n58065 );
and ( n59239 , n58065 , n58071 );
and ( n59240 , n58061 , n58071 );
or ( n59241 , n59238 , n59239 , n59240 );
and ( n59242 , n58051 , n58052 );
and ( n59243 , n58052 , n58054 );
and ( n59244 , n58051 , n58054 );
or ( n59245 , n59242 , n59243 , n59244 );
and ( n59246 , n18144 , n8669 );
and ( n59247 , n19324 , n8243 );
xor ( n59248 , n59246 , n59247 );
and ( n59249 , n20233 , n7662 );
xor ( n59250 , n59248 , n59249 );
xor ( n59251 , n59245 , n59250 );
and ( n59252 , n15758 , n10977 );
and ( n59253 , n16637 , n10239 );
xor ( n59254 , n59252 , n59253 );
and ( n59255 , n17512 , n9348 );
xor ( n59256 , n59254 , n59255 );
xor ( n59257 , n59251 , n59256 );
xor ( n59258 , n59241 , n59257 );
and ( n59259 , n58067 , n58068 );
and ( n59260 , n58068 , n58070 );
and ( n59261 , n58067 , n58070 );
or ( n59262 , n59259 , n59260 , n59261 );
and ( n59263 , n58098 , n58099 );
and ( n59264 , n58099 , n58101 );
and ( n59265 , n58098 , n58101 );
or ( n59266 , n59263 , n59264 , n59265 );
xor ( n59267 , n59262 , n59266 );
buf ( n59268 , n13322 );
and ( n59269 , n14118 , n12531 );
xor ( n59270 , n59268 , n59269 );
and ( n59271 , n14938 , n11718 );
xor ( n59272 , n59270 , n59271 );
xor ( n59273 , n59267 , n59272 );
xor ( n59274 , n59258 , n59273 );
xor ( n59275 , n59237 , n59274 );
xor ( n59276 , n59207 , n59275 );
and ( n59277 , n58088 , n58092 );
and ( n59278 , n58092 , n58109 );
and ( n59279 , n58088 , n58109 );
or ( n59280 , n59277 , n59278 , n59279 );
and ( n59281 , n58139 , n58154 );
and ( n59282 , n58154 , n58171 );
and ( n59283 , n58139 , n58171 );
or ( n59284 , n59281 , n59282 , n59283 );
xor ( n59285 , n59280 , n59284 );
and ( n59286 , n58097 , n58102 );
and ( n59287 , n58102 , n58108 );
and ( n59288 , n58097 , n58108 );
or ( n59289 , n59286 , n59287 , n59288 );
and ( n59290 , n58143 , n58147 );
and ( n59291 , n58147 , n58153 );
and ( n59292 , n58143 , n58153 );
or ( n59293 , n59290 , n59291 , n59292 );
xor ( n59294 , n59289 , n59293 );
and ( n59295 , n58104 , n58105 );
and ( n59296 , n58105 , n58107 );
and ( n59297 , n58104 , n58107 );
or ( n59298 , n59295 , n59296 , n59297 );
and ( n59299 , n11015 , n15691 );
and ( n59300 , n11769 , n14838 );
xor ( n59301 , n59299 , n59300 );
and ( n59302 , n12320 , n14044 );
xor ( n59303 , n59301 , n59302 );
xor ( n59304 , n59298 , n59303 );
and ( n59305 , n8718 , n18407 );
and ( n59306 , n9400 , n17422 );
xor ( n59307 , n59305 , n59306 );
and ( n59308 , n10291 , n16550 );
xor ( n59309 , n59307 , n59308 );
xor ( n59310 , n59304 , n59309 );
xor ( n59311 , n59294 , n59310 );
xor ( n59312 , n59285 , n59311 );
xor ( n59313 , n59276 , n59312 );
xor ( n59314 , n59203 , n59313 );
xor ( n59315 , n59194 , n59314 );
not ( n59316 , n3182 );
and ( n59317 , n34193 , n3182 );
nor ( n59318 , n59316 , n59317 );
and ( n59319 , n3545 , n32999 );
xor ( n59320 , n59318 , n59319 );
and ( n59321 , n3801 , n31761 );
xor ( n59322 , n59320 , n59321 );
and ( n59323 , n58135 , n58172 );
and ( n59324 , n58172 , n58198 );
and ( n59325 , n58135 , n58198 );
or ( n59326 , n59323 , n59324 , n59325 );
and ( n59327 , n58177 , n58181 );
and ( n59328 , n58181 , n58197 );
and ( n59329 , n58177 , n58197 );
or ( n59330 , n59327 , n59328 , n59329 );
and ( n59331 , n58159 , n58164 );
and ( n59332 , n58164 , n58170 );
and ( n59333 , n58159 , n58170 );
or ( n59334 , n59331 , n59332 , n59333 );
and ( n59335 , n58149 , n58150 );
and ( n59336 , n58150 , n58152 );
and ( n59337 , n58149 , n58152 );
or ( n59338 , n59335 , n59336 , n59337 );
and ( n59339 , n58160 , n58161 );
and ( n59340 , n58161 , n58163 );
and ( n59341 , n58160 , n58163 );
or ( n59342 , n59339 , n59340 , n59341 );
xor ( n59343 , n59338 , n59342 );
and ( n59344 , n7385 , n20976 );
and ( n59345 , n7808 , n20156 );
xor ( n59346 , n59344 , n59345 );
and ( n59347 , n8079 , n19222 );
xor ( n59348 , n59346 , n59347 );
xor ( n59349 , n59343 , n59348 );
xor ( n59350 , n59334 , n59349 );
and ( n59351 , n58166 , n58167 );
and ( n59352 , n58167 , n58169 );
and ( n59353 , n58166 , n58169 );
or ( n59354 , n59351 , n59352 , n59353 );
and ( n59355 , n6187 , n24137 );
and ( n59356 , n6569 , n23075 );
xor ( n59357 , n59355 , n59356 );
and ( n59358 , n6816 , n22065 );
xor ( n59359 , n59357 , n59358 );
xor ( n59360 , n59354 , n59359 );
and ( n59361 , n4959 , n27296 );
and ( n59362 , n5459 , n26216 );
xor ( n59363 , n59361 , n59362 );
and ( n59364 , n5819 , n25163 );
xor ( n59365 , n59363 , n59364 );
xor ( n59366 , n59360 , n59365 );
xor ( n59367 , n59350 , n59366 );
xor ( n59368 , n59330 , n59367 );
and ( n59369 , n58115 , n58118 );
and ( n59370 , n58118 , n58124 );
and ( n59371 , n58115 , n58124 );
or ( n59372 , n59369 , n59370 , n59371 );
and ( n59373 , n58186 , n58190 );
and ( n59374 , n58190 , n58196 );
and ( n59375 , n58186 , n58196 );
or ( n59376 , n59373 , n59374 , n59375 );
xor ( n59377 , n59372 , n59376 );
and ( n59378 , n58192 , n58193 );
and ( n59379 , n58193 , n58195 );
and ( n59380 , n58192 , n58195 );
or ( n59381 , n59378 , n59379 , n59380 );
and ( n59382 , n58120 , n58121 );
and ( n59383 , n58121 , n58123 );
and ( n59384 , n58120 , n58123 );
or ( n59385 , n59382 , n59383 , n59384 );
xor ( n59386 , n59381 , n59385 );
and ( n59387 , n4132 , n30629 );
and ( n59388 , n4438 , n29508 );
xor ( n59389 , n59387 , n59388 );
and ( n59390 , n4766 , n28406 );
xor ( n59391 , n59389 , n59390 );
xor ( n59392 , n59386 , n59391 );
xor ( n59393 , n59377 , n59392 );
xor ( n59394 , n59368 , n59393 );
xor ( n59395 , n59326 , n59394 );
xor ( n59396 , n59322 , n59395 );
xor ( n59397 , n59315 , n59396 );
xor ( n59398 , n59193 , n59397 );
xor ( n59399 , n59111 , n59398 );
xor ( n59400 , n59102 , n59399 );
and ( n59401 , n57897 , n57900 );
and ( n59402 , n57900 , n58204 );
and ( n59403 , n57897 , n58204 );
or ( n59404 , n59401 , n59402 , n59403 );
xor ( n59405 , n59400 , n59404 );
and ( n59406 , n58205 , n58209 );
and ( n59407 , n58210 , n58213 );
or ( n59408 , n59406 , n59407 );
xor ( n59409 , n59405 , n59408 );
buf ( n59410 , n59409 );
buf ( n59411 , n59410 );
not ( n59412 , n59411 );
nor ( n59413 , n59412 , n8739 );
xor ( n59414 , n59094 , n59413 );
and ( n59415 , n57893 , n58218 );
and ( n59416 , n58219 , n58222 );
or ( n59417 , n59415 , n59416 );
xor ( n59418 , n59414 , n59417 );
buf ( n59419 , n59418 );
buf ( n59420 , n59419 );
not ( n59421 , n59420 );
buf ( n59422 , n583 );
not ( n59423 , n59422 );
nor ( n59424 , n59421 , n59423 );
xor ( n59425 , n58720 , n59424 );
xor ( n59426 , n58234 , n58717 );
nor ( n59427 , n58226 , n59423 );
and ( n59428 , n59426 , n59427 );
xor ( n59429 , n59426 , n59427 );
xor ( n59430 , n58238 , n58715 );
nor ( n59431 , n57031 , n59423 );
and ( n59432 , n59430 , n59431 );
xor ( n59433 , n59430 , n59431 );
xor ( n59434 , n58242 , n58713 );
nor ( n59435 , n55835 , n59423 );
and ( n59436 , n59434 , n59435 );
xor ( n59437 , n59434 , n59435 );
xor ( n59438 , n58246 , n58711 );
nor ( n59439 , n54638 , n59423 );
and ( n59440 , n59438 , n59439 );
xor ( n59441 , n59438 , n59439 );
xor ( n59442 , n58250 , n58709 );
nor ( n59443 , n53441 , n59423 );
and ( n59444 , n59442 , n59443 );
xor ( n59445 , n59442 , n59443 );
xor ( n59446 , n58254 , n58707 );
nor ( n59447 , n52247 , n59423 );
and ( n59448 , n59446 , n59447 );
xor ( n59449 , n59446 , n59447 );
xor ( n59450 , n58258 , n58705 );
nor ( n59451 , n51049 , n59423 );
and ( n59452 , n59450 , n59451 );
xor ( n59453 , n59450 , n59451 );
xor ( n59454 , n58262 , n58703 );
nor ( n59455 , n49850 , n59423 );
and ( n59456 , n59454 , n59455 );
xor ( n59457 , n59454 , n59455 );
xor ( n59458 , n58266 , n58701 );
nor ( n59459 , n48650 , n59423 );
and ( n59460 , n59458 , n59459 );
xor ( n59461 , n59458 , n59459 );
xor ( n59462 , n58270 , n58699 );
nor ( n59463 , n47449 , n59423 );
and ( n59464 , n59462 , n59463 );
xor ( n59465 , n59462 , n59463 );
xor ( n59466 , n58274 , n58697 );
nor ( n59467 , n46248 , n59423 );
and ( n59468 , n59466 , n59467 );
xor ( n59469 , n59466 , n59467 );
xor ( n59470 , n58278 , n58695 );
nor ( n59471 , n45047 , n59423 );
and ( n59472 , n59470 , n59471 );
xor ( n59473 , n59470 , n59471 );
xor ( n59474 , n58282 , n58693 );
nor ( n59475 , n43843 , n59423 );
and ( n59476 , n59474 , n59475 );
xor ( n59477 , n59474 , n59475 );
xor ( n59478 , n58286 , n58691 );
nor ( n59479 , n42641 , n59423 );
and ( n59480 , n59478 , n59479 );
xor ( n59481 , n59478 , n59479 );
xor ( n59482 , n58290 , n58689 );
nor ( n59483 , n41437 , n59423 );
and ( n59484 , n59482 , n59483 );
xor ( n59485 , n59482 , n59483 );
xor ( n59486 , n58294 , n58687 );
nor ( n59487 , n40232 , n59423 );
and ( n59488 , n59486 , n59487 );
xor ( n59489 , n59486 , n59487 );
xor ( n59490 , n58298 , n58685 );
nor ( n59491 , n39027 , n59423 );
and ( n59492 , n59490 , n59491 );
xor ( n59493 , n59490 , n59491 );
xor ( n59494 , n58302 , n58683 );
nor ( n59495 , n37825 , n59423 );
and ( n59496 , n59494 , n59495 );
xor ( n59497 , n59494 , n59495 );
xor ( n59498 , n58306 , n58681 );
nor ( n59499 , n36620 , n59423 );
and ( n59500 , n59498 , n59499 );
xor ( n59501 , n59498 , n59499 );
xor ( n59502 , n58310 , n58679 );
nor ( n59503 , n35419 , n59423 );
and ( n59504 , n59502 , n59503 );
xor ( n59505 , n59502 , n59503 );
xor ( n59506 , n58314 , n58677 );
nor ( n59507 , n34224 , n59423 );
and ( n59508 , n59506 , n59507 );
xor ( n59509 , n59506 , n59507 );
xor ( n59510 , n58318 , n58675 );
nor ( n59511 , n33033 , n59423 );
and ( n59512 , n59510 , n59511 );
xor ( n59513 , n59510 , n59511 );
xor ( n59514 , n58322 , n58673 );
nor ( n59515 , n31867 , n59423 );
and ( n59516 , n59514 , n59515 );
xor ( n59517 , n59514 , n59515 );
xor ( n59518 , n58326 , n58671 );
nor ( n59519 , n30725 , n59423 );
and ( n59520 , n59518 , n59519 );
xor ( n59521 , n59518 , n59519 );
xor ( n59522 , n58330 , n58669 );
nor ( n59523 , n29596 , n59423 );
and ( n59524 , n59522 , n59523 );
xor ( n59525 , n59522 , n59523 );
xor ( n59526 , n58334 , n58667 );
nor ( n59527 , n28487 , n59423 );
and ( n59528 , n59526 , n59527 );
xor ( n59529 , n59526 , n59527 );
xor ( n59530 , n58338 , n58665 );
nor ( n59531 , n27397 , n59423 );
and ( n59532 , n59530 , n59531 );
xor ( n59533 , n59530 , n59531 );
xor ( n59534 , n58342 , n58663 );
nor ( n59535 , n26326 , n59423 );
and ( n59536 , n59534 , n59535 );
xor ( n59537 , n59534 , n59535 );
xor ( n59538 , n58346 , n58661 );
nor ( n59539 , n25272 , n59423 );
and ( n59540 , n59538 , n59539 );
xor ( n59541 , n59538 , n59539 );
xor ( n59542 , n58350 , n58659 );
nor ( n59543 , n24242 , n59423 );
and ( n59544 , n59542 , n59543 );
xor ( n59545 , n59542 , n59543 );
xor ( n59546 , n58354 , n58657 );
nor ( n59547 , n23225 , n59423 );
and ( n59548 , n59546 , n59547 );
xor ( n59549 , n59546 , n59547 );
xor ( n59550 , n58358 , n58655 );
nor ( n59551 , n22231 , n59423 );
and ( n59552 , n59550 , n59551 );
xor ( n59553 , n59550 , n59551 );
xor ( n59554 , n58362 , n58653 );
nor ( n59555 , n21258 , n59423 );
and ( n59556 , n59554 , n59555 );
xor ( n59557 , n59554 , n59555 );
xor ( n59558 , n58366 , n58651 );
nor ( n59559 , n20303 , n59423 );
and ( n59560 , n59558 , n59559 );
xor ( n59561 , n59558 , n59559 );
xor ( n59562 , n58370 , n58649 );
nor ( n59563 , n19365 , n59423 );
and ( n59564 , n59562 , n59563 );
xor ( n59565 , n59562 , n59563 );
xor ( n59566 , n58374 , n58647 );
nor ( n59567 , n18448 , n59423 );
and ( n59568 , n59566 , n59567 );
xor ( n59569 , n59566 , n59567 );
xor ( n59570 , n58378 , n58645 );
nor ( n59571 , n17548 , n59423 );
and ( n59572 , n59570 , n59571 );
xor ( n59573 , n59570 , n59571 );
xor ( n59574 , n58382 , n58643 );
nor ( n59575 , n16669 , n59423 );
and ( n59576 , n59574 , n59575 );
xor ( n59577 , n59574 , n59575 );
xor ( n59578 , n58386 , n58641 );
nor ( n59579 , n15809 , n59423 );
and ( n59580 , n59578 , n59579 );
xor ( n59581 , n59578 , n59579 );
xor ( n59582 , n58390 , n58639 );
nor ( n59583 , n14968 , n59423 );
and ( n59584 , n59582 , n59583 );
xor ( n59585 , n59582 , n59583 );
xor ( n59586 , n58394 , n58637 );
nor ( n59587 , n14147 , n59423 );
and ( n59588 , n59586 , n59587 );
xor ( n59589 , n59586 , n59587 );
xor ( n59590 , n58398 , n58635 );
nor ( n59591 , n13349 , n59423 );
and ( n59592 , n59590 , n59591 );
xor ( n59593 , n59590 , n59591 );
xor ( n59594 , n58402 , n58633 );
nor ( n59595 , n12564 , n59423 );
and ( n59596 , n59594 , n59595 );
xor ( n59597 , n59594 , n59595 );
xor ( n59598 , n58406 , n58631 );
nor ( n59599 , n11799 , n59423 );
and ( n59600 , n59598 , n59599 );
xor ( n59601 , n59598 , n59599 );
xor ( n59602 , n58410 , n58629 );
nor ( n59603 , n11050 , n59423 );
and ( n59604 , n59602 , n59603 );
xor ( n59605 , n59602 , n59603 );
xor ( n59606 , n58414 , n58627 );
nor ( n59607 , n10321 , n59423 );
and ( n59608 , n59606 , n59607 );
xor ( n59609 , n59606 , n59607 );
xor ( n59610 , n58418 , n58625 );
nor ( n59611 , n9429 , n59423 );
and ( n59612 , n59610 , n59611 );
xor ( n59613 , n59610 , n59611 );
xor ( n59614 , n58422 , n58623 );
nor ( n59615 , n8949 , n59423 );
and ( n59616 , n59614 , n59615 );
xor ( n59617 , n59614 , n59615 );
xor ( n59618 , n58426 , n58621 );
nor ( n59619 , n9437 , n59423 );
and ( n59620 , n59618 , n59619 );
xor ( n59621 , n59618 , n59619 );
xor ( n59622 , n58430 , n58619 );
nor ( n59623 , n9446 , n59423 );
and ( n59624 , n59622 , n59623 );
xor ( n59625 , n59622 , n59623 );
xor ( n59626 , n58434 , n58617 );
nor ( n59627 , n9455 , n59423 );
and ( n59628 , n59626 , n59627 );
xor ( n59629 , n59626 , n59627 );
xor ( n59630 , n58438 , n58615 );
nor ( n59631 , n9464 , n59423 );
and ( n59632 , n59630 , n59631 );
xor ( n59633 , n59630 , n59631 );
xor ( n59634 , n58442 , n58613 );
nor ( n59635 , n9473 , n59423 );
and ( n59636 , n59634 , n59635 );
xor ( n59637 , n59634 , n59635 );
xor ( n59638 , n58446 , n58611 );
nor ( n59639 , n9482 , n59423 );
and ( n59640 , n59638 , n59639 );
xor ( n59641 , n59638 , n59639 );
xor ( n59642 , n58450 , n58609 );
nor ( n59643 , n9491 , n59423 );
and ( n59644 , n59642 , n59643 );
xor ( n59645 , n59642 , n59643 );
xor ( n59646 , n58454 , n58607 );
nor ( n59647 , n9500 , n59423 );
and ( n59648 , n59646 , n59647 );
xor ( n59649 , n59646 , n59647 );
xor ( n59650 , n58458 , n58605 );
nor ( n59651 , n9509 , n59423 );
and ( n59652 , n59650 , n59651 );
xor ( n59653 , n59650 , n59651 );
xor ( n59654 , n58462 , n58603 );
nor ( n59655 , n9518 , n59423 );
and ( n59656 , n59654 , n59655 );
xor ( n59657 , n59654 , n59655 );
xor ( n59658 , n58466 , n58601 );
nor ( n59659 , n9527 , n59423 );
and ( n59660 , n59658 , n59659 );
xor ( n59661 , n59658 , n59659 );
xor ( n59662 , n58470 , n58599 );
nor ( n59663 , n9536 , n59423 );
and ( n59664 , n59662 , n59663 );
xor ( n59665 , n59662 , n59663 );
xor ( n59666 , n58474 , n58597 );
nor ( n59667 , n9545 , n59423 );
and ( n59668 , n59666 , n59667 );
xor ( n59669 , n59666 , n59667 );
xor ( n59670 , n58478 , n58595 );
nor ( n59671 , n9554 , n59423 );
and ( n59672 , n59670 , n59671 );
xor ( n59673 , n59670 , n59671 );
xor ( n59674 , n58482 , n58593 );
nor ( n59675 , n9563 , n59423 );
and ( n59676 , n59674 , n59675 );
xor ( n59677 , n59674 , n59675 );
xor ( n59678 , n58486 , n58591 );
nor ( n59679 , n9572 , n59423 );
and ( n59680 , n59678 , n59679 );
xor ( n59681 , n59678 , n59679 );
xor ( n59682 , n58490 , n58589 );
nor ( n59683 , n9581 , n59423 );
and ( n59684 , n59682 , n59683 );
xor ( n59685 , n59682 , n59683 );
xor ( n59686 , n58494 , n58587 );
nor ( n59687 , n9590 , n59423 );
and ( n59688 , n59686 , n59687 );
xor ( n59689 , n59686 , n59687 );
xor ( n59690 , n58498 , n58585 );
nor ( n59691 , n9599 , n59423 );
and ( n59692 , n59690 , n59691 );
xor ( n59693 , n59690 , n59691 );
xor ( n59694 , n58502 , n58583 );
nor ( n59695 , n9608 , n59423 );
and ( n59696 , n59694 , n59695 );
xor ( n59697 , n59694 , n59695 );
xor ( n59698 , n58506 , n58581 );
nor ( n59699 , n9617 , n59423 );
and ( n59700 , n59698 , n59699 );
xor ( n59701 , n59698 , n59699 );
xor ( n59702 , n58510 , n58579 );
nor ( n59703 , n9626 , n59423 );
and ( n59704 , n59702 , n59703 );
xor ( n59705 , n59702 , n59703 );
xor ( n59706 , n58514 , n58577 );
nor ( n59707 , n9635 , n59423 );
and ( n59708 , n59706 , n59707 );
xor ( n59709 , n59706 , n59707 );
xor ( n59710 , n58518 , n58575 );
nor ( n59711 , n9644 , n59423 );
and ( n59712 , n59710 , n59711 );
xor ( n59713 , n59710 , n59711 );
xor ( n59714 , n58522 , n58573 );
nor ( n59715 , n9653 , n59423 );
and ( n59716 , n59714 , n59715 );
xor ( n59717 , n59714 , n59715 );
xor ( n59718 , n58526 , n58571 );
nor ( n59719 , n9662 , n59423 );
and ( n59720 , n59718 , n59719 );
xor ( n59721 , n59718 , n59719 );
xor ( n59722 , n58530 , n58569 );
nor ( n59723 , n9671 , n59423 );
and ( n59724 , n59722 , n59723 );
xor ( n59725 , n59722 , n59723 );
xor ( n59726 , n58534 , n58567 );
nor ( n59727 , n9680 , n59423 );
and ( n59728 , n59726 , n59727 );
xor ( n59729 , n59726 , n59727 );
xor ( n59730 , n58538 , n58565 );
nor ( n59731 , n9689 , n59423 );
and ( n59732 , n59730 , n59731 );
xor ( n59733 , n59730 , n59731 );
xor ( n59734 , n58542 , n58563 );
nor ( n59735 , n9698 , n59423 );
and ( n59736 , n59734 , n59735 );
xor ( n59737 , n59734 , n59735 );
xor ( n59738 , n58546 , n58561 );
nor ( n59739 , n9707 , n59423 );
and ( n59740 , n59738 , n59739 );
xor ( n59741 , n59738 , n59739 );
xor ( n59742 , n58550 , n58559 );
nor ( n59743 , n9716 , n59423 );
and ( n59744 , n59742 , n59743 );
xor ( n59745 , n59742 , n59743 );
xor ( n59746 , n58554 , n58557 );
nor ( n59747 , n9725 , n59423 );
and ( n59748 , n59746 , n59747 );
xor ( n59749 , n59746 , n59747 );
xor ( n59750 , n58555 , n58556 );
nor ( n59751 , n9734 , n59423 );
and ( n59752 , n59750 , n59751 );
xor ( n59753 , n59750 , n59751 );
nor ( n59754 , n9752 , n58228 );
nor ( n59755 , n9743 , n59423 );
and ( n59756 , n59754 , n59755 );
and ( n59757 , n59753 , n59756 );
or ( n59758 , n59752 , n59757 );
and ( n59759 , n59749 , n59758 );
or ( n59760 , n59748 , n59759 );
and ( n59761 , n59745 , n59760 );
or ( n59762 , n59744 , n59761 );
and ( n59763 , n59741 , n59762 );
or ( n59764 , n59740 , n59763 );
and ( n59765 , n59737 , n59764 );
or ( n59766 , n59736 , n59765 );
and ( n59767 , n59733 , n59766 );
or ( n59768 , n59732 , n59767 );
and ( n59769 , n59729 , n59768 );
or ( n59770 , n59728 , n59769 );
and ( n59771 , n59725 , n59770 );
or ( n59772 , n59724 , n59771 );
and ( n59773 , n59721 , n59772 );
or ( n59774 , n59720 , n59773 );
and ( n59775 , n59717 , n59774 );
or ( n59776 , n59716 , n59775 );
and ( n59777 , n59713 , n59776 );
or ( n59778 , n59712 , n59777 );
and ( n59779 , n59709 , n59778 );
or ( n59780 , n59708 , n59779 );
and ( n59781 , n59705 , n59780 );
or ( n59782 , n59704 , n59781 );
and ( n59783 , n59701 , n59782 );
or ( n59784 , n59700 , n59783 );
and ( n59785 , n59697 , n59784 );
or ( n59786 , n59696 , n59785 );
and ( n59787 , n59693 , n59786 );
or ( n59788 , n59692 , n59787 );
and ( n59789 , n59689 , n59788 );
or ( n59790 , n59688 , n59789 );
and ( n59791 , n59685 , n59790 );
or ( n59792 , n59684 , n59791 );
and ( n59793 , n59681 , n59792 );
or ( n59794 , n59680 , n59793 );
and ( n59795 , n59677 , n59794 );
or ( n59796 , n59676 , n59795 );
and ( n59797 , n59673 , n59796 );
or ( n59798 , n59672 , n59797 );
and ( n59799 , n59669 , n59798 );
or ( n59800 , n59668 , n59799 );
and ( n59801 , n59665 , n59800 );
or ( n59802 , n59664 , n59801 );
and ( n59803 , n59661 , n59802 );
or ( n59804 , n59660 , n59803 );
and ( n59805 , n59657 , n59804 );
or ( n59806 , n59656 , n59805 );
and ( n59807 , n59653 , n59806 );
or ( n59808 , n59652 , n59807 );
and ( n59809 , n59649 , n59808 );
or ( n59810 , n59648 , n59809 );
and ( n59811 , n59645 , n59810 );
or ( n59812 , n59644 , n59811 );
and ( n59813 , n59641 , n59812 );
or ( n59814 , n59640 , n59813 );
and ( n59815 , n59637 , n59814 );
or ( n59816 , n59636 , n59815 );
and ( n59817 , n59633 , n59816 );
or ( n59818 , n59632 , n59817 );
and ( n59819 , n59629 , n59818 );
or ( n59820 , n59628 , n59819 );
and ( n59821 , n59625 , n59820 );
or ( n59822 , n59624 , n59821 );
and ( n59823 , n59621 , n59822 );
or ( n59824 , n59620 , n59823 );
and ( n59825 , n59617 , n59824 );
or ( n59826 , n59616 , n59825 );
and ( n59827 , n59613 , n59826 );
or ( n59828 , n59612 , n59827 );
and ( n59829 , n59609 , n59828 );
or ( n59830 , n59608 , n59829 );
and ( n59831 , n59605 , n59830 );
or ( n59832 , n59604 , n59831 );
and ( n59833 , n59601 , n59832 );
or ( n59834 , n59600 , n59833 );
and ( n59835 , n59597 , n59834 );
or ( n59836 , n59596 , n59835 );
and ( n59837 , n59593 , n59836 );
or ( n59838 , n59592 , n59837 );
and ( n59839 , n59589 , n59838 );
or ( n59840 , n59588 , n59839 );
and ( n59841 , n59585 , n59840 );
or ( n59842 , n59584 , n59841 );
and ( n59843 , n59581 , n59842 );
or ( n59844 , n59580 , n59843 );
and ( n59845 , n59577 , n59844 );
or ( n59846 , n59576 , n59845 );
and ( n59847 , n59573 , n59846 );
or ( n59848 , n59572 , n59847 );
and ( n59849 , n59569 , n59848 );
or ( n59850 , n59568 , n59849 );
and ( n59851 , n59565 , n59850 );
or ( n59852 , n59564 , n59851 );
and ( n59853 , n59561 , n59852 );
or ( n59854 , n59560 , n59853 );
and ( n59855 , n59557 , n59854 );
or ( n59856 , n59556 , n59855 );
and ( n59857 , n59553 , n59856 );
or ( n59858 , n59552 , n59857 );
and ( n59859 , n59549 , n59858 );
or ( n59860 , n59548 , n59859 );
and ( n59861 , n59545 , n59860 );
or ( n59862 , n59544 , n59861 );
and ( n59863 , n59541 , n59862 );
or ( n59864 , n59540 , n59863 );
and ( n59865 , n59537 , n59864 );
or ( n59866 , n59536 , n59865 );
and ( n59867 , n59533 , n59866 );
or ( n59868 , n59532 , n59867 );
and ( n59869 , n59529 , n59868 );
or ( n59870 , n59528 , n59869 );
and ( n59871 , n59525 , n59870 );
or ( n59872 , n59524 , n59871 );
and ( n59873 , n59521 , n59872 );
or ( n59874 , n59520 , n59873 );
and ( n59875 , n59517 , n59874 );
or ( n59876 , n59516 , n59875 );
and ( n59877 , n59513 , n59876 );
or ( n59878 , n59512 , n59877 );
and ( n59879 , n59509 , n59878 );
or ( n59880 , n59508 , n59879 );
and ( n59881 , n59505 , n59880 );
or ( n59882 , n59504 , n59881 );
and ( n59883 , n59501 , n59882 );
or ( n59884 , n59500 , n59883 );
and ( n59885 , n59497 , n59884 );
or ( n59886 , n59496 , n59885 );
and ( n59887 , n59493 , n59886 );
or ( n59888 , n59492 , n59887 );
and ( n59889 , n59489 , n59888 );
or ( n59890 , n59488 , n59889 );
and ( n59891 , n59485 , n59890 );
or ( n59892 , n59484 , n59891 );
and ( n59893 , n59481 , n59892 );
or ( n59894 , n59480 , n59893 );
and ( n59895 , n59477 , n59894 );
or ( n59896 , n59476 , n59895 );
and ( n59897 , n59473 , n59896 );
or ( n59898 , n59472 , n59897 );
and ( n59899 , n59469 , n59898 );
or ( n59900 , n59468 , n59899 );
and ( n59901 , n59465 , n59900 );
or ( n59902 , n59464 , n59901 );
and ( n59903 , n59461 , n59902 );
or ( n59904 , n59460 , n59903 );
and ( n59905 , n59457 , n59904 );
or ( n59906 , n59456 , n59905 );
and ( n59907 , n59453 , n59906 );
or ( n59908 , n59452 , n59907 );
and ( n59909 , n59449 , n59908 );
or ( n59910 , n59448 , n59909 );
and ( n59911 , n59445 , n59910 );
or ( n59912 , n59444 , n59911 );
and ( n59913 , n59441 , n59912 );
or ( n59914 , n59440 , n59913 );
and ( n59915 , n59437 , n59914 );
or ( n59916 , n59436 , n59915 );
and ( n59917 , n59433 , n59916 );
or ( n59918 , n59432 , n59917 );
and ( n59919 , n59429 , n59918 );
or ( n59920 , n59428 , n59919 );
xor ( n59921 , n59425 , n59920 );
and ( n59922 , n33403 , n3569 );
nor ( n59923 , n3570 , n59922 );
nor ( n59924 , n3853 , n32231 );
xor ( n59925 , n59923 , n59924 );
and ( n59926 , n58722 , n58723 );
and ( n59927 , n58724 , n58727 );
or ( n59928 , n59926 , n59927 );
xor ( n59929 , n59925 , n59928 );
nor ( n59930 , n4151 , n31083 );
xor ( n59931 , n59929 , n59930 );
and ( n59932 , n58728 , n58729 );
and ( n59933 , n58730 , n58733 );
or ( n59934 , n59932 , n59933 );
xor ( n59935 , n59931 , n59934 );
nor ( n59936 , n4458 , n29948 );
xor ( n59937 , n59935 , n59936 );
and ( n59938 , n58734 , n58735 );
and ( n59939 , n58736 , n58739 );
or ( n59940 , n59938 , n59939 );
xor ( n59941 , n59937 , n59940 );
nor ( n59942 , n4786 , n28833 );
xor ( n59943 , n59941 , n59942 );
and ( n59944 , n58740 , n58741 );
and ( n59945 , n58742 , n58745 );
or ( n59946 , n59944 , n59945 );
xor ( n59947 , n59943 , n59946 );
nor ( n59948 , n5126 , n27737 );
xor ( n59949 , n59947 , n59948 );
and ( n59950 , n58746 , n58747 );
and ( n59951 , n58748 , n58751 );
or ( n59952 , n59950 , n59951 );
xor ( n59953 , n59949 , n59952 );
nor ( n59954 , n5477 , n26660 );
xor ( n59955 , n59953 , n59954 );
and ( n59956 , n58752 , n58753 );
and ( n59957 , n58754 , n58757 );
or ( n59958 , n59956 , n59957 );
xor ( n59959 , n59955 , n59958 );
nor ( n59960 , n5838 , n25600 );
xor ( n59961 , n59959 , n59960 );
and ( n59962 , n58758 , n58759 );
and ( n59963 , n58760 , n58763 );
or ( n59964 , n59962 , n59963 );
xor ( n59965 , n59961 , n59964 );
nor ( n59966 , n6212 , n24564 );
xor ( n59967 , n59965 , n59966 );
and ( n59968 , n58764 , n58765 );
and ( n59969 , n58766 , n58769 );
or ( n59970 , n59968 , n59969 );
xor ( n59971 , n59967 , n59970 );
nor ( n59972 , n6596 , n23541 );
xor ( n59973 , n59971 , n59972 );
and ( n59974 , n58770 , n58771 );
and ( n59975 , n58772 , n58775 );
or ( n59976 , n59974 , n59975 );
xor ( n59977 , n59973 , n59976 );
nor ( n59978 , n6997 , n22541 );
xor ( n59979 , n59977 , n59978 );
and ( n59980 , n58776 , n58777 );
and ( n59981 , n58778 , n58781 );
or ( n59982 , n59980 , n59981 );
xor ( n59983 , n59979 , n59982 );
nor ( n59984 , n7413 , n21562 );
xor ( n59985 , n59983 , n59984 );
and ( n59986 , n58782 , n58783 );
and ( n59987 , n58784 , n58787 );
or ( n59988 , n59986 , n59987 );
xor ( n59989 , n59985 , n59988 );
nor ( n59990 , n7841 , n20601 );
xor ( n59991 , n59989 , n59990 );
and ( n59992 , n58788 , n58789 );
and ( n59993 , n58790 , n58793 );
or ( n59994 , n59992 , n59993 );
xor ( n59995 , n59991 , n59994 );
nor ( n59996 , n8281 , n19657 );
xor ( n59997 , n59995 , n59996 );
and ( n59998 , n58794 , n58795 );
and ( n59999 , n58796 , n58799 );
or ( n60000 , n59998 , n59999 );
xor ( n60001 , n59997 , n60000 );
nor ( n60002 , n8737 , n18734 );
xor ( n60003 , n60001 , n60002 );
and ( n60004 , n58800 , n58801 );
and ( n60005 , n58802 , n58805 );
or ( n60006 , n60004 , n60005 );
xor ( n60007 , n60003 , n60006 );
nor ( n60008 , n9420 , n17828 );
xor ( n60009 , n60007 , n60008 );
and ( n60010 , n58806 , n58807 );
and ( n60011 , n58808 , n58811 );
or ( n60012 , n60010 , n60011 );
xor ( n60013 , n60009 , n60012 );
nor ( n60014 , n10312 , n16943 );
xor ( n60015 , n60013 , n60014 );
and ( n60016 , n58812 , n58813 );
and ( n60017 , n58814 , n58817 );
or ( n60018 , n60016 , n60017 );
xor ( n60019 , n60015 , n60018 );
nor ( n60020 , n11041 , n16077 );
xor ( n60021 , n60019 , n60020 );
and ( n60022 , n58818 , n58819 );
and ( n60023 , n58820 , n58823 );
or ( n60024 , n60022 , n60023 );
xor ( n60025 , n60021 , n60024 );
nor ( n60026 , n11790 , n15230 );
xor ( n60027 , n60025 , n60026 );
and ( n60028 , n58824 , n58825 );
and ( n60029 , n58826 , n58829 );
or ( n60030 , n60028 , n60029 );
xor ( n60031 , n60027 , n60030 );
nor ( n60032 , n12555 , n14403 );
xor ( n60033 , n60031 , n60032 );
and ( n60034 , n58830 , n58831 );
and ( n60035 , n58832 , n58835 );
or ( n60036 , n60034 , n60035 );
xor ( n60037 , n60033 , n60036 );
nor ( n60038 , n13340 , n13599 );
xor ( n60039 , n60037 , n60038 );
and ( n60040 , n58836 , n58837 );
and ( n60041 , n58838 , n58841 );
or ( n60042 , n60040 , n60041 );
xor ( n60043 , n60039 , n60042 );
nor ( n60044 , n14138 , n12808 );
xor ( n60045 , n60043 , n60044 );
and ( n60046 , n58842 , n58843 );
and ( n60047 , n58844 , n58847 );
or ( n60048 , n60046 , n60047 );
xor ( n60049 , n60045 , n60048 );
nor ( n60050 , n14959 , n12037 );
xor ( n60051 , n60049 , n60050 );
and ( n60052 , n58848 , n58849 );
and ( n60053 , n58850 , n58853 );
or ( n60054 , n60052 , n60053 );
xor ( n60055 , n60051 , n60054 );
nor ( n60056 , n15800 , n11282 );
xor ( n60057 , n60055 , n60056 );
and ( n60058 , n58854 , n58855 );
and ( n60059 , n58856 , n58859 );
or ( n60060 , n60058 , n60059 );
xor ( n60061 , n60057 , n60060 );
nor ( n60062 , n16660 , n10547 );
xor ( n60063 , n60061 , n60062 );
and ( n60064 , n58860 , n58861 );
and ( n60065 , n58862 , n58865 );
or ( n60066 , n60064 , n60065 );
xor ( n60067 , n60063 , n60066 );
nor ( n60068 , n17539 , n9829 );
xor ( n60069 , n60067 , n60068 );
and ( n60070 , n58866 , n58867 );
and ( n60071 , n58868 , n58871 );
or ( n60072 , n60070 , n60071 );
xor ( n60073 , n60069 , n60072 );
nor ( n60074 , n18439 , n8955 );
xor ( n60075 , n60073 , n60074 );
and ( n60076 , n58872 , n58873 );
and ( n60077 , n58874 , n58877 );
or ( n60078 , n60076 , n60077 );
xor ( n60079 , n60075 , n60078 );
nor ( n60080 , n19356 , n603 );
xor ( n60081 , n60079 , n60080 );
and ( n60082 , n58878 , n58879 );
and ( n60083 , n58880 , n58883 );
or ( n60084 , n60082 , n60083 );
xor ( n60085 , n60081 , n60084 );
nor ( n60086 , n20294 , n652 );
xor ( n60087 , n60085 , n60086 );
and ( n60088 , n58884 , n58885 );
and ( n60089 , n58886 , n58889 );
or ( n60090 , n60088 , n60089 );
xor ( n60091 , n60087 , n60090 );
nor ( n60092 , n21249 , n624 );
xor ( n60093 , n60091 , n60092 );
and ( n60094 , n58890 , n58891 );
and ( n60095 , n58892 , n58895 );
or ( n60096 , n60094 , n60095 );
xor ( n60097 , n60093 , n60096 );
nor ( n60098 , n22222 , n648 );
xor ( n60099 , n60097 , n60098 );
and ( n60100 , n58896 , n58897 );
and ( n60101 , n58898 , n58901 );
or ( n60102 , n60100 , n60101 );
xor ( n60103 , n60099 , n60102 );
nor ( n60104 , n23216 , n686 );
xor ( n60105 , n60103 , n60104 );
and ( n60106 , n58902 , n58903 );
and ( n60107 , n58904 , n58907 );
or ( n60108 , n60106 , n60107 );
xor ( n60109 , n60105 , n60108 );
nor ( n60110 , n24233 , n735 );
xor ( n60111 , n60109 , n60110 );
and ( n60112 , n58908 , n58909 );
and ( n60113 , n58910 , n58913 );
or ( n60114 , n60112 , n60113 );
xor ( n60115 , n60111 , n60114 );
nor ( n60116 , n25263 , n798 );
xor ( n60117 , n60115 , n60116 );
and ( n60118 , n58914 , n58915 );
and ( n60119 , n58916 , n58919 );
or ( n60120 , n60118 , n60119 );
xor ( n60121 , n60117 , n60120 );
nor ( n60122 , n26317 , n870 );
xor ( n60123 , n60121 , n60122 );
and ( n60124 , n58920 , n58921 );
and ( n60125 , n58922 , n58925 );
or ( n60126 , n60124 , n60125 );
xor ( n60127 , n60123 , n60126 );
nor ( n60128 , n27388 , n960 );
xor ( n60129 , n60127 , n60128 );
and ( n60130 , n58926 , n58927 );
and ( n60131 , n58928 , n58931 );
or ( n60132 , n60130 , n60131 );
xor ( n60133 , n60129 , n60132 );
nor ( n60134 , n28478 , n1064 );
xor ( n60135 , n60133 , n60134 );
and ( n60136 , n58932 , n58933 );
and ( n60137 , n58934 , n58937 );
or ( n60138 , n60136 , n60137 );
xor ( n60139 , n60135 , n60138 );
nor ( n60140 , n29587 , n1178 );
xor ( n60141 , n60139 , n60140 );
and ( n60142 , n58938 , n58939 );
and ( n60143 , n58940 , n58943 );
or ( n60144 , n60142 , n60143 );
xor ( n60145 , n60141 , n60144 );
nor ( n60146 , n30716 , n1305 );
xor ( n60147 , n60145 , n60146 );
and ( n60148 , n58944 , n58945 );
and ( n60149 , n58946 , n58949 );
or ( n60150 , n60148 , n60149 );
xor ( n60151 , n60147 , n60150 );
nor ( n60152 , n31858 , n1447 );
xor ( n60153 , n60151 , n60152 );
and ( n60154 , n58950 , n58951 );
and ( n60155 , n58952 , n58955 );
or ( n60156 , n60154 , n60155 );
xor ( n60157 , n60153 , n60156 );
nor ( n60158 , n33024 , n1600 );
xor ( n60159 , n60157 , n60158 );
and ( n60160 , n58956 , n58957 );
and ( n60161 , n58958 , n58961 );
or ( n60162 , n60160 , n60161 );
xor ( n60163 , n60159 , n60162 );
nor ( n60164 , n34215 , n1768 );
xor ( n60165 , n60163 , n60164 );
and ( n60166 , n58962 , n58963 );
and ( n60167 , n58964 , n58967 );
or ( n60168 , n60166 , n60167 );
xor ( n60169 , n60165 , n60168 );
nor ( n60170 , n35410 , n1947 );
xor ( n60171 , n60169 , n60170 );
and ( n60172 , n58968 , n58969 );
and ( n60173 , n58970 , n58973 );
or ( n60174 , n60172 , n60173 );
xor ( n60175 , n60171 , n60174 );
nor ( n60176 , n36611 , n2139 );
xor ( n60177 , n60175 , n60176 );
and ( n60178 , n58974 , n58975 );
and ( n60179 , n58976 , n58979 );
or ( n60180 , n60178 , n60179 );
xor ( n60181 , n60177 , n60180 );
nor ( n60182 , n37816 , n2345 );
xor ( n60183 , n60181 , n60182 );
and ( n60184 , n58980 , n58981 );
and ( n60185 , n58982 , n58985 );
or ( n60186 , n60184 , n60185 );
xor ( n60187 , n60183 , n60186 );
nor ( n60188 , n39018 , n2568 );
xor ( n60189 , n60187 , n60188 );
and ( n60190 , n58986 , n58987 );
and ( n60191 , n58988 , n58991 );
or ( n60192 , n60190 , n60191 );
xor ( n60193 , n60189 , n60192 );
nor ( n60194 , n40223 , n2799 );
xor ( n60195 , n60193 , n60194 );
and ( n60196 , n58992 , n58993 );
and ( n60197 , n58994 , n58997 );
or ( n60198 , n60196 , n60197 );
xor ( n60199 , n60195 , n60198 );
nor ( n60200 , n41428 , n3045 );
xor ( n60201 , n60199 , n60200 );
and ( n60202 , n58998 , n58999 );
and ( n60203 , n59000 , n59003 );
or ( n60204 , n60202 , n60203 );
xor ( n60205 , n60201 , n60204 );
nor ( n60206 , n42632 , n3302 );
xor ( n60207 , n60205 , n60206 );
and ( n60208 , n59004 , n59005 );
and ( n60209 , n59006 , n59009 );
or ( n60210 , n60208 , n60209 );
xor ( n60211 , n60207 , n60210 );
nor ( n60212 , n43834 , n3572 );
xor ( n60213 , n60211 , n60212 );
and ( n60214 , n59010 , n59011 );
and ( n60215 , n59012 , n59015 );
or ( n60216 , n60214 , n60215 );
xor ( n60217 , n60213 , n60216 );
nor ( n60218 , n45038 , n3855 );
xor ( n60219 , n60217 , n60218 );
and ( n60220 , n59016 , n59017 );
and ( n60221 , n59018 , n59021 );
or ( n60222 , n60220 , n60221 );
xor ( n60223 , n60219 , n60222 );
nor ( n60224 , n46239 , n4153 );
xor ( n60225 , n60223 , n60224 );
and ( n60226 , n59022 , n59023 );
and ( n60227 , n59024 , n59027 );
or ( n60228 , n60226 , n60227 );
xor ( n60229 , n60225 , n60228 );
nor ( n60230 , n47440 , n4460 );
xor ( n60231 , n60229 , n60230 );
and ( n60232 , n59028 , n59029 );
and ( n60233 , n59030 , n59033 );
or ( n60234 , n60232 , n60233 );
xor ( n60235 , n60231 , n60234 );
nor ( n60236 , n48641 , n4788 );
xor ( n60237 , n60235 , n60236 );
and ( n60238 , n59034 , n59035 );
and ( n60239 , n59036 , n59039 );
or ( n60240 , n60238 , n60239 );
xor ( n60241 , n60237 , n60240 );
nor ( n60242 , n49841 , n5128 );
xor ( n60243 , n60241 , n60242 );
and ( n60244 , n59040 , n59041 );
and ( n60245 , n59042 , n59045 );
or ( n60246 , n60244 , n60245 );
xor ( n60247 , n60243 , n60246 );
nor ( n60248 , n51040 , n5479 );
xor ( n60249 , n60247 , n60248 );
and ( n60250 , n59046 , n59047 );
and ( n60251 , n59048 , n59051 );
or ( n60252 , n60250 , n60251 );
xor ( n60253 , n60249 , n60252 );
nor ( n60254 , n52238 , n5840 );
xor ( n60255 , n60253 , n60254 );
and ( n60256 , n59052 , n59053 );
and ( n60257 , n59054 , n59057 );
or ( n60258 , n60256 , n60257 );
xor ( n60259 , n60255 , n60258 );
nor ( n60260 , n53432 , n6214 );
xor ( n60261 , n60259 , n60260 );
and ( n60262 , n59058 , n59059 );
and ( n60263 , n59060 , n59063 );
or ( n60264 , n60262 , n60263 );
xor ( n60265 , n60261 , n60264 );
nor ( n60266 , n54629 , n6598 );
xor ( n60267 , n60265 , n60266 );
and ( n60268 , n59064 , n59065 );
and ( n60269 , n59066 , n59069 );
or ( n60270 , n60268 , n60269 );
xor ( n60271 , n60267 , n60270 );
nor ( n60272 , n55826 , n6999 );
xor ( n60273 , n60271 , n60272 );
and ( n60274 , n59070 , n59071 );
and ( n60275 , n59072 , n59075 );
or ( n60276 , n60274 , n60275 );
xor ( n60277 , n60273 , n60276 );
nor ( n60278 , n57022 , n7415 );
xor ( n60279 , n60277 , n60278 );
and ( n60280 , n59076 , n59077 );
and ( n60281 , n59078 , n59081 );
or ( n60282 , n60280 , n60281 );
xor ( n60283 , n60279 , n60282 );
nor ( n60284 , n58217 , n7843 );
xor ( n60285 , n60283 , n60284 );
and ( n60286 , n59082 , n59083 );
and ( n60287 , n59084 , n59087 );
or ( n60288 , n60286 , n60287 );
xor ( n60289 , n60285 , n60288 );
nor ( n60290 , n59412 , n8283 );
xor ( n60291 , n60289 , n60290 );
and ( n60292 , n59088 , n59089 );
and ( n60293 , n59090 , n59093 );
or ( n60294 , n60292 , n60293 );
xor ( n60295 , n60291 , n60294 );
and ( n60296 , n59106 , n59110 );
and ( n60297 , n59110 , n59398 );
and ( n60298 , n59106 , n59398 );
or ( n60299 , n60296 , n60297 , n60298 );
and ( n60300 , n33774 , n3495 );
not ( n60301 , n3495 );
nor ( n60302 , n60300 , n60301 );
xor ( n60303 , n60299 , n60302 );
and ( n60304 , n59119 , n59123 );
and ( n60305 , n59123 , n59191 );
and ( n60306 , n59119 , n59191 );
or ( n60307 , n60304 , n60305 , n60306 );
and ( n60308 , n59115 , n59192 );
and ( n60309 , n59192 , n59397 );
and ( n60310 , n59115 , n59397 );
or ( n60311 , n60308 , n60309 , n60310 );
xor ( n60312 , n60307 , n60311 );
and ( n60313 , n59194 , n59314 );
and ( n60314 , n59314 , n59396 );
and ( n60315 , n59194 , n59396 );
or ( n60316 , n60313 , n60314 , n60315 );
and ( n60317 , n59128 , n59132 );
and ( n60318 , n59132 , n59190 );
and ( n60319 , n59128 , n59190 );
or ( n60320 , n60317 , n60318 , n60319 );
and ( n60321 , n59198 , n59202 );
and ( n60322 , n59202 , n59313 );
and ( n60323 , n59198 , n59313 );
or ( n60324 , n60321 , n60322 , n60323 );
xor ( n60325 , n60320 , n60324 );
and ( n60326 , n59159 , n59163 );
and ( n60327 , n59163 , n59169 );
and ( n60328 , n59159 , n59169 );
or ( n60329 , n60326 , n60327 , n60328 );
and ( n60330 , n59137 , n59141 );
and ( n60331 , n59141 , n59189 );
and ( n60332 , n59137 , n59189 );
or ( n60333 , n60330 , n60331 , n60332 );
xor ( n60334 , n60329 , n60333 );
and ( n60335 , n59146 , n59150 );
and ( n60336 , n59150 , n59188 );
and ( n60337 , n59146 , n59188 );
or ( n60338 , n60335 , n60336 , n60337 );
and ( n60339 , n59211 , n59236 );
and ( n60340 , n59236 , n59274 );
and ( n60341 , n59211 , n59274 );
or ( n60342 , n60339 , n60340 , n60341 );
xor ( n60343 , n60338 , n60342 );
and ( n60344 , n59155 , n59170 );
and ( n60345 , n59170 , n59187 );
and ( n60346 , n59155 , n59187 );
or ( n60347 , n60344 , n60345 , n60346 );
and ( n60348 , n59215 , n59219 );
and ( n60349 , n59219 , n59235 );
and ( n60350 , n59215 , n59235 );
or ( n60351 , n60348 , n60349 , n60350 );
xor ( n60352 , n60347 , n60351 );
and ( n60353 , n59175 , n59180 );
and ( n60354 , n59180 , n59186 );
and ( n60355 , n59175 , n59186 );
or ( n60356 , n60353 , n60354 , n60355 );
and ( n60357 , n59165 , n59166 );
and ( n60358 , n59166 , n59168 );
and ( n60359 , n59165 , n59168 );
or ( n60360 , n60357 , n60358 , n60359 );
and ( n60361 , n59176 , n59177 );
and ( n60362 , n59177 , n59179 );
and ( n60363 , n59176 , n59179 );
or ( n60364 , n60361 , n60362 , n60363 );
xor ( n60365 , n60360 , n60364 );
and ( n60366 , n30695 , n4403 );
and ( n60367 , n31836 , n4102 );
xor ( n60368 , n60366 , n60367 );
and ( n60369 , n32649 , n3749 );
xor ( n60370 , n60368 , n60369 );
xor ( n60371 , n60365 , n60370 );
xor ( n60372 , n60356 , n60371 );
and ( n60373 , n59182 , n59183 );
and ( n60374 , n59183 , n59185 );
and ( n60375 , n59182 , n59185 );
or ( n60376 , n60373 , n60374 , n60375 );
and ( n60377 , n27361 , n5408 );
and ( n60378 , n28456 , n5103 );
xor ( n60379 , n60377 , n60378 );
and ( n60380 , n29559 , n4730 );
xor ( n60381 , n60379 , n60380 );
xor ( n60382 , n60376 , n60381 );
and ( n60383 , n24214 , n6504 );
and ( n60384 , n25243 , n6132 );
xor ( n60385 , n60383 , n60384 );
and ( n60386 , n26296 , n5765 );
xor ( n60387 , n60385 , n60386 );
xor ( n60388 , n60382 , n60387 );
xor ( n60389 , n60372 , n60388 );
xor ( n60390 , n60352 , n60389 );
xor ( n60391 , n60343 , n60390 );
xor ( n60392 , n60334 , n60391 );
xor ( n60393 , n60325 , n60392 );
xor ( n60394 , n60316 , n60393 );
and ( n60395 , n59322 , n59395 );
and ( n60396 , n59207 , n59275 );
and ( n60397 , n59275 , n59312 );
and ( n60398 , n59207 , n59312 );
or ( n60399 , n60396 , n60397 , n60398 );
and ( n60400 , n59326 , n59394 );
xor ( n60401 , n60399 , n60400 );
and ( n60402 , n59280 , n59284 );
and ( n60403 , n59284 , n59311 );
and ( n60404 , n59280 , n59311 );
or ( n60405 , n60402 , n60403 , n60404 );
and ( n60406 , n59241 , n59257 );
and ( n60407 , n59257 , n59273 );
and ( n60408 , n59241 , n59273 );
or ( n60409 , n60406 , n60407 , n60408 );
and ( n60410 , n59224 , n59228 );
and ( n60411 , n59228 , n59234 );
and ( n60412 , n59224 , n59234 );
or ( n60413 , n60410 , n60411 , n60412 );
and ( n60414 , n59245 , n59250 );
and ( n60415 , n59250 , n59256 );
and ( n60416 , n59245 , n59256 );
or ( n60417 , n60414 , n60415 , n60416 );
xor ( n60418 , n60413 , n60417 );
and ( n60419 , n59230 , n59231 );
and ( n60420 , n59231 , n59233 );
and ( n60421 , n59230 , n59233 );
or ( n60422 , n60419 , n60420 , n60421 );
and ( n60423 , n59246 , n59247 );
and ( n60424 , n59247 , n59249 );
and ( n60425 , n59246 , n59249 );
or ( n60426 , n60423 , n60424 , n60425 );
xor ( n60427 , n60422 , n60426 );
and ( n60428 , n21216 , n7662 );
and ( n60429 , n22186 , n7310 );
xor ( n60430 , n60428 , n60429 );
and ( n60431 , n22892 , n6971 );
xor ( n60432 , n60430 , n60431 );
xor ( n60433 , n60427 , n60432 );
xor ( n60434 , n60418 , n60433 );
xor ( n60435 , n60409 , n60434 );
and ( n60436 , n59262 , n59266 );
and ( n60437 , n59266 , n59272 );
and ( n60438 , n59262 , n59272 );
or ( n60439 , n60436 , n60437 , n60438 );
and ( n60440 , n59252 , n59253 );
and ( n60441 , n59253 , n59255 );
and ( n60442 , n59252 , n59255 );
or ( n60443 , n60440 , n60441 , n60442 );
and ( n60444 , n18144 , n9348 );
and ( n60445 , n19324 , n8669 );
xor ( n60446 , n60444 , n60445 );
and ( n60447 , n20233 , n8243 );
xor ( n60448 , n60446 , n60447 );
xor ( n60449 , n60443 , n60448 );
and ( n60450 , n15758 , n11718 );
and ( n60451 , n16637 , n10977 );
xor ( n60452 , n60450 , n60451 );
and ( n60453 , n17512 , n10239 );
xor ( n60454 , n60452 , n60453 );
xor ( n60455 , n60449 , n60454 );
xor ( n60456 , n60439 , n60455 );
and ( n60457 , n59268 , n59269 );
and ( n60458 , n59269 , n59271 );
and ( n60459 , n59268 , n59271 );
or ( n60460 , n60457 , n60458 , n60459 );
and ( n60461 , n59299 , n59300 );
and ( n60462 , n59300 , n59302 );
and ( n60463 , n59299 , n59302 );
or ( n60464 , n60461 , n60462 , n60463 );
xor ( n60465 , n60460 , n60464 );
and ( n60466 , n14938 , n12531 );
buf ( n60467 , n60466 );
xor ( n60468 , n60465 , n60467 );
xor ( n60469 , n60456 , n60468 );
xor ( n60470 , n60435 , n60469 );
xor ( n60471 , n60405 , n60470 );
and ( n60472 , n59289 , n59293 );
and ( n60473 , n59293 , n59310 );
and ( n60474 , n59289 , n59310 );
or ( n60475 , n60472 , n60473 , n60474 );
and ( n60476 , n59334 , n59349 );
and ( n60477 , n59349 , n59366 );
and ( n60478 , n59334 , n59366 );
or ( n60479 , n60476 , n60477 , n60478 );
xor ( n60480 , n60475 , n60479 );
and ( n60481 , n59298 , n59303 );
and ( n60482 , n59303 , n59309 );
and ( n60483 , n59298 , n59309 );
or ( n60484 , n60481 , n60482 , n60483 );
and ( n60485 , n59338 , n59342 );
and ( n60486 , n59342 , n59348 );
and ( n60487 , n59338 , n59348 );
or ( n60488 , n60485 , n60486 , n60487 );
xor ( n60489 , n60484 , n60488 );
and ( n60490 , n59305 , n59306 );
and ( n60491 , n59306 , n59308 );
and ( n60492 , n59305 , n59308 );
or ( n60493 , n60490 , n60491 , n60492 );
and ( n60494 , n11015 , n16550 );
and ( n60495 , n11769 , n15691 );
xor ( n60496 , n60494 , n60495 );
and ( n60497 , n12320 , n14838 );
xor ( n60498 , n60496 , n60497 );
xor ( n60499 , n60493 , n60498 );
and ( n60500 , n8718 , n19222 );
and ( n60501 , n9400 , n18407 );
xor ( n60502 , n60500 , n60501 );
and ( n60503 , n10291 , n17422 );
xor ( n60504 , n60502 , n60503 );
xor ( n60505 , n60499 , n60504 );
xor ( n60506 , n60489 , n60505 );
xor ( n60507 , n60480 , n60506 );
xor ( n60508 , n60471 , n60507 );
xor ( n60509 , n60401 , n60508 );
xor ( n60510 , n60395 , n60509 );
not ( n60511 , n3545 );
and ( n60512 , n34193 , n3545 );
nor ( n60513 , n60511 , n60512 );
and ( n60514 , n3801 , n32999 );
xor ( n60515 , n60513 , n60514 );
and ( n60516 , n59330 , n59367 );
and ( n60517 , n59367 , n59393 );
and ( n60518 , n59330 , n59393 );
or ( n60519 , n60516 , n60517 , n60518 );
and ( n60520 , n59372 , n59376 );
and ( n60521 , n59376 , n59392 );
and ( n60522 , n59372 , n59392 );
or ( n60523 , n60520 , n60521 , n60522 );
and ( n60524 , n59354 , n59359 );
and ( n60525 , n59359 , n59365 );
and ( n60526 , n59354 , n59365 );
or ( n60527 , n60524 , n60525 , n60526 );
and ( n60528 , n59344 , n59345 );
and ( n60529 , n59345 , n59347 );
and ( n60530 , n59344 , n59347 );
or ( n60531 , n60528 , n60529 , n60530 );
and ( n60532 , n59355 , n59356 );
and ( n60533 , n59356 , n59358 );
and ( n60534 , n59355 , n59358 );
or ( n60535 , n60532 , n60533 , n60534 );
xor ( n60536 , n60531 , n60535 );
and ( n60537 , n7385 , n22065 );
and ( n60538 , n7808 , n20976 );
xor ( n60539 , n60537 , n60538 );
and ( n60540 , n8079 , n20156 );
xor ( n60541 , n60539 , n60540 );
xor ( n60542 , n60536 , n60541 );
xor ( n60543 , n60527 , n60542 );
and ( n60544 , n59361 , n59362 );
and ( n60545 , n59362 , n59364 );
and ( n60546 , n59361 , n59364 );
or ( n60547 , n60544 , n60545 , n60546 );
and ( n60548 , n6187 , n25163 );
and ( n60549 , n6569 , n24137 );
xor ( n60550 , n60548 , n60549 );
and ( n60551 , n6816 , n23075 );
xor ( n60552 , n60550 , n60551 );
xor ( n60553 , n60547 , n60552 );
and ( n60554 , n4959 , n28406 );
and ( n60555 , n5459 , n27296 );
xor ( n60556 , n60554 , n60555 );
and ( n60557 , n5819 , n26216 );
xor ( n60558 , n60556 , n60557 );
xor ( n60559 , n60553 , n60558 );
xor ( n60560 , n60543 , n60559 );
xor ( n60561 , n60523 , n60560 );
and ( n60562 , n59381 , n59385 );
and ( n60563 , n59385 , n59391 );
and ( n60564 , n59381 , n59391 );
or ( n60565 , n60562 , n60563 , n60564 );
and ( n60566 , n59318 , n59319 );
and ( n60567 , n59319 , n59321 );
and ( n60568 , n59318 , n59321 );
or ( n60569 , n60566 , n60567 , n60568 );
and ( n60570 , n59387 , n59388 );
and ( n60571 , n59388 , n59390 );
and ( n60572 , n59387 , n59390 );
or ( n60573 , n60570 , n60571 , n60572 );
xor ( n60574 , n60569 , n60573 );
and ( n60575 , n4132 , n31761 );
and ( n60576 , n4438 , n30629 );
xor ( n60577 , n60575 , n60576 );
and ( n60578 , n4766 , n29508 );
xor ( n60579 , n60577 , n60578 );
xor ( n60580 , n60574 , n60579 );
xor ( n60581 , n60565 , n60580 );
xor ( n60582 , n60561 , n60581 );
xor ( n60583 , n60519 , n60582 );
xor ( n60584 , n60515 , n60583 );
xor ( n60585 , n60510 , n60584 );
xor ( n60586 , n60394 , n60585 );
xor ( n60587 , n60312 , n60586 );
xor ( n60588 , n60303 , n60587 );
and ( n60589 , n59098 , n59101 );
and ( n60590 , n59101 , n59399 );
and ( n60591 , n59098 , n59399 );
or ( n60592 , n60589 , n60590 , n60591 );
xor ( n60593 , n60588 , n60592 );
and ( n60594 , n59400 , n59404 );
and ( n60595 , n59405 , n59408 );
or ( n60596 , n60594 , n60595 );
xor ( n60597 , n60593 , n60596 );
buf ( n60598 , n60597 );
buf ( n60599 , n60598 );
not ( n60600 , n60599 );
nor ( n60601 , n60600 , n8739 );
xor ( n60602 , n60295 , n60601 );
and ( n60603 , n59094 , n59413 );
and ( n60604 , n59414 , n59417 );
or ( n60605 , n60603 , n60604 );
xor ( n60606 , n60602 , n60605 );
buf ( n60607 , n60606 );
buf ( n60608 , n60607 );
not ( n60609 , n60608 );
buf ( n60610 , n584 );
not ( n60611 , n60610 );
nor ( n60612 , n60609 , n60611 );
xor ( n60613 , n59921 , n60612 );
xor ( n60614 , n59429 , n59918 );
nor ( n60615 , n59421 , n60611 );
and ( n60616 , n60614 , n60615 );
xor ( n60617 , n60614 , n60615 );
xor ( n60618 , n59433 , n59916 );
nor ( n60619 , n58226 , n60611 );
and ( n60620 , n60618 , n60619 );
xor ( n60621 , n60618 , n60619 );
xor ( n60622 , n59437 , n59914 );
nor ( n60623 , n57031 , n60611 );
and ( n60624 , n60622 , n60623 );
xor ( n60625 , n60622 , n60623 );
xor ( n60626 , n59441 , n59912 );
nor ( n60627 , n55835 , n60611 );
and ( n60628 , n60626 , n60627 );
xor ( n60629 , n60626 , n60627 );
xor ( n60630 , n59445 , n59910 );
nor ( n60631 , n54638 , n60611 );
and ( n60632 , n60630 , n60631 );
xor ( n60633 , n60630 , n60631 );
xor ( n60634 , n59449 , n59908 );
nor ( n60635 , n53441 , n60611 );
and ( n60636 , n60634 , n60635 );
xor ( n60637 , n60634 , n60635 );
xor ( n60638 , n59453 , n59906 );
nor ( n60639 , n52247 , n60611 );
and ( n60640 , n60638 , n60639 );
xor ( n60641 , n60638 , n60639 );
xor ( n60642 , n59457 , n59904 );
nor ( n60643 , n51049 , n60611 );
and ( n60644 , n60642 , n60643 );
xor ( n60645 , n60642 , n60643 );
xor ( n60646 , n59461 , n59902 );
nor ( n60647 , n49850 , n60611 );
and ( n60648 , n60646 , n60647 );
xor ( n60649 , n60646 , n60647 );
xor ( n60650 , n59465 , n59900 );
nor ( n60651 , n48650 , n60611 );
and ( n60652 , n60650 , n60651 );
xor ( n60653 , n60650 , n60651 );
xor ( n60654 , n59469 , n59898 );
nor ( n60655 , n47449 , n60611 );
and ( n60656 , n60654 , n60655 );
xor ( n60657 , n60654 , n60655 );
xor ( n60658 , n59473 , n59896 );
nor ( n60659 , n46248 , n60611 );
and ( n60660 , n60658 , n60659 );
xor ( n60661 , n60658 , n60659 );
xor ( n60662 , n59477 , n59894 );
nor ( n60663 , n45047 , n60611 );
and ( n60664 , n60662 , n60663 );
xor ( n60665 , n60662 , n60663 );
xor ( n60666 , n59481 , n59892 );
nor ( n60667 , n43843 , n60611 );
and ( n60668 , n60666 , n60667 );
xor ( n60669 , n60666 , n60667 );
xor ( n60670 , n59485 , n59890 );
nor ( n60671 , n42641 , n60611 );
and ( n60672 , n60670 , n60671 );
xor ( n60673 , n60670 , n60671 );
xor ( n60674 , n59489 , n59888 );
nor ( n60675 , n41437 , n60611 );
and ( n60676 , n60674 , n60675 );
xor ( n60677 , n60674 , n60675 );
xor ( n60678 , n59493 , n59886 );
nor ( n60679 , n40232 , n60611 );
and ( n60680 , n60678 , n60679 );
xor ( n60681 , n60678 , n60679 );
xor ( n60682 , n59497 , n59884 );
nor ( n60683 , n39027 , n60611 );
and ( n60684 , n60682 , n60683 );
xor ( n60685 , n60682 , n60683 );
xor ( n60686 , n59501 , n59882 );
nor ( n60687 , n37825 , n60611 );
and ( n60688 , n60686 , n60687 );
xor ( n60689 , n60686 , n60687 );
xor ( n60690 , n59505 , n59880 );
nor ( n60691 , n36620 , n60611 );
and ( n60692 , n60690 , n60691 );
xor ( n60693 , n60690 , n60691 );
xor ( n60694 , n59509 , n59878 );
nor ( n60695 , n35419 , n60611 );
and ( n60696 , n60694 , n60695 );
xor ( n60697 , n60694 , n60695 );
xor ( n60698 , n59513 , n59876 );
nor ( n60699 , n34224 , n60611 );
and ( n60700 , n60698 , n60699 );
xor ( n60701 , n60698 , n60699 );
xor ( n60702 , n59517 , n59874 );
nor ( n60703 , n33033 , n60611 );
and ( n60704 , n60702 , n60703 );
xor ( n60705 , n60702 , n60703 );
xor ( n60706 , n59521 , n59872 );
nor ( n60707 , n31867 , n60611 );
and ( n60708 , n60706 , n60707 );
xor ( n60709 , n60706 , n60707 );
xor ( n60710 , n59525 , n59870 );
nor ( n60711 , n30725 , n60611 );
and ( n60712 , n60710 , n60711 );
xor ( n60713 , n60710 , n60711 );
xor ( n60714 , n59529 , n59868 );
nor ( n60715 , n29596 , n60611 );
and ( n60716 , n60714 , n60715 );
xor ( n60717 , n60714 , n60715 );
xor ( n60718 , n59533 , n59866 );
nor ( n60719 , n28487 , n60611 );
and ( n60720 , n60718 , n60719 );
xor ( n60721 , n60718 , n60719 );
xor ( n60722 , n59537 , n59864 );
nor ( n60723 , n27397 , n60611 );
and ( n60724 , n60722 , n60723 );
xor ( n60725 , n60722 , n60723 );
xor ( n60726 , n59541 , n59862 );
nor ( n60727 , n26326 , n60611 );
and ( n60728 , n60726 , n60727 );
xor ( n60729 , n60726 , n60727 );
xor ( n60730 , n59545 , n59860 );
nor ( n60731 , n25272 , n60611 );
and ( n60732 , n60730 , n60731 );
xor ( n60733 , n60730 , n60731 );
xor ( n60734 , n59549 , n59858 );
nor ( n60735 , n24242 , n60611 );
and ( n60736 , n60734 , n60735 );
xor ( n60737 , n60734 , n60735 );
xor ( n60738 , n59553 , n59856 );
nor ( n60739 , n23225 , n60611 );
and ( n60740 , n60738 , n60739 );
xor ( n60741 , n60738 , n60739 );
xor ( n60742 , n59557 , n59854 );
nor ( n60743 , n22231 , n60611 );
and ( n60744 , n60742 , n60743 );
xor ( n60745 , n60742 , n60743 );
xor ( n60746 , n59561 , n59852 );
nor ( n60747 , n21258 , n60611 );
and ( n60748 , n60746 , n60747 );
xor ( n60749 , n60746 , n60747 );
xor ( n60750 , n59565 , n59850 );
nor ( n60751 , n20303 , n60611 );
and ( n60752 , n60750 , n60751 );
xor ( n60753 , n60750 , n60751 );
xor ( n60754 , n59569 , n59848 );
nor ( n60755 , n19365 , n60611 );
and ( n60756 , n60754 , n60755 );
xor ( n60757 , n60754 , n60755 );
xor ( n60758 , n59573 , n59846 );
nor ( n60759 , n18448 , n60611 );
and ( n60760 , n60758 , n60759 );
xor ( n60761 , n60758 , n60759 );
xor ( n60762 , n59577 , n59844 );
nor ( n60763 , n17548 , n60611 );
and ( n60764 , n60762 , n60763 );
xor ( n60765 , n60762 , n60763 );
xor ( n60766 , n59581 , n59842 );
nor ( n60767 , n16669 , n60611 );
and ( n60768 , n60766 , n60767 );
xor ( n60769 , n60766 , n60767 );
xor ( n60770 , n59585 , n59840 );
nor ( n60771 , n15809 , n60611 );
and ( n60772 , n60770 , n60771 );
xor ( n60773 , n60770 , n60771 );
xor ( n60774 , n59589 , n59838 );
nor ( n60775 , n14968 , n60611 );
and ( n60776 , n60774 , n60775 );
xor ( n60777 , n60774 , n60775 );
xor ( n60778 , n59593 , n59836 );
nor ( n60779 , n14147 , n60611 );
and ( n60780 , n60778 , n60779 );
xor ( n60781 , n60778 , n60779 );
xor ( n60782 , n59597 , n59834 );
nor ( n60783 , n13349 , n60611 );
and ( n60784 , n60782 , n60783 );
xor ( n60785 , n60782 , n60783 );
xor ( n60786 , n59601 , n59832 );
nor ( n60787 , n12564 , n60611 );
and ( n60788 , n60786 , n60787 );
xor ( n60789 , n60786 , n60787 );
xor ( n60790 , n59605 , n59830 );
nor ( n60791 , n11799 , n60611 );
and ( n60792 , n60790 , n60791 );
xor ( n60793 , n60790 , n60791 );
xor ( n60794 , n59609 , n59828 );
nor ( n60795 , n11050 , n60611 );
and ( n60796 , n60794 , n60795 );
xor ( n60797 , n60794 , n60795 );
xor ( n60798 , n59613 , n59826 );
nor ( n60799 , n10321 , n60611 );
and ( n60800 , n60798 , n60799 );
xor ( n60801 , n60798 , n60799 );
xor ( n60802 , n59617 , n59824 );
nor ( n60803 , n9429 , n60611 );
and ( n60804 , n60802 , n60803 );
xor ( n60805 , n60802 , n60803 );
xor ( n60806 , n59621 , n59822 );
nor ( n60807 , n8949 , n60611 );
and ( n60808 , n60806 , n60807 );
xor ( n60809 , n60806 , n60807 );
xor ( n60810 , n59625 , n59820 );
nor ( n60811 , n9437 , n60611 );
and ( n60812 , n60810 , n60811 );
xor ( n60813 , n60810 , n60811 );
xor ( n60814 , n59629 , n59818 );
nor ( n60815 , n9446 , n60611 );
and ( n60816 , n60814 , n60815 );
xor ( n60817 , n60814 , n60815 );
xor ( n60818 , n59633 , n59816 );
nor ( n60819 , n9455 , n60611 );
and ( n60820 , n60818 , n60819 );
xor ( n60821 , n60818 , n60819 );
xor ( n60822 , n59637 , n59814 );
nor ( n60823 , n9464 , n60611 );
and ( n60824 , n60822 , n60823 );
xor ( n60825 , n60822 , n60823 );
xor ( n60826 , n59641 , n59812 );
nor ( n60827 , n9473 , n60611 );
and ( n60828 , n60826 , n60827 );
xor ( n60829 , n60826 , n60827 );
xor ( n60830 , n59645 , n59810 );
nor ( n60831 , n9482 , n60611 );
and ( n60832 , n60830 , n60831 );
xor ( n60833 , n60830 , n60831 );
xor ( n60834 , n59649 , n59808 );
nor ( n60835 , n9491 , n60611 );
and ( n60836 , n60834 , n60835 );
xor ( n60837 , n60834 , n60835 );
xor ( n60838 , n59653 , n59806 );
nor ( n60839 , n9500 , n60611 );
and ( n60840 , n60838 , n60839 );
xor ( n60841 , n60838 , n60839 );
xor ( n60842 , n59657 , n59804 );
nor ( n60843 , n9509 , n60611 );
and ( n60844 , n60842 , n60843 );
xor ( n60845 , n60842 , n60843 );
xor ( n60846 , n59661 , n59802 );
nor ( n60847 , n9518 , n60611 );
and ( n60848 , n60846 , n60847 );
xor ( n60849 , n60846 , n60847 );
xor ( n60850 , n59665 , n59800 );
nor ( n60851 , n9527 , n60611 );
and ( n60852 , n60850 , n60851 );
xor ( n60853 , n60850 , n60851 );
xor ( n60854 , n59669 , n59798 );
nor ( n60855 , n9536 , n60611 );
and ( n60856 , n60854 , n60855 );
xor ( n60857 , n60854 , n60855 );
xor ( n60858 , n59673 , n59796 );
nor ( n60859 , n9545 , n60611 );
and ( n60860 , n60858 , n60859 );
xor ( n60861 , n60858 , n60859 );
xor ( n60862 , n59677 , n59794 );
nor ( n60863 , n9554 , n60611 );
and ( n60864 , n60862 , n60863 );
xor ( n60865 , n60862 , n60863 );
xor ( n60866 , n59681 , n59792 );
nor ( n60867 , n9563 , n60611 );
and ( n60868 , n60866 , n60867 );
xor ( n60869 , n60866 , n60867 );
xor ( n60870 , n59685 , n59790 );
nor ( n60871 , n9572 , n60611 );
and ( n60872 , n60870 , n60871 );
xor ( n60873 , n60870 , n60871 );
xor ( n60874 , n59689 , n59788 );
nor ( n60875 , n9581 , n60611 );
and ( n60876 , n60874 , n60875 );
xor ( n60877 , n60874 , n60875 );
xor ( n60878 , n59693 , n59786 );
nor ( n60879 , n9590 , n60611 );
and ( n60880 , n60878 , n60879 );
xor ( n60881 , n60878 , n60879 );
xor ( n60882 , n59697 , n59784 );
nor ( n60883 , n9599 , n60611 );
and ( n60884 , n60882 , n60883 );
xor ( n60885 , n60882 , n60883 );
xor ( n60886 , n59701 , n59782 );
nor ( n60887 , n9608 , n60611 );
and ( n60888 , n60886 , n60887 );
xor ( n60889 , n60886 , n60887 );
xor ( n60890 , n59705 , n59780 );
nor ( n60891 , n9617 , n60611 );
and ( n60892 , n60890 , n60891 );
xor ( n60893 , n60890 , n60891 );
xor ( n60894 , n59709 , n59778 );
nor ( n60895 , n9626 , n60611 );
and ( n60896 , n60894 , n60895 );
xor ( n60897 , n60894 , n60895 );
xor ( n60898 , n59713 , n59776 );
nor ( n60899 , n9635 , n60611 );
and ( n60900 , n60898 , n60899 );
xor ( n60901 , n60898 , n60899 );
xor ( n60902 , n59717 , n59774 );
nor ( n60903 , n9644 , n60611 );
and ( n60904 , n60902 , n60903 );
xor ( n60905 , n60902 , n60903 );
xor ( n60906 , n59721 , n59772 );
nor ( n60907 , n9653 , n60611 );
and ( n60908 , n60906 , n60907 );
xor ( n60909 , n60906 , n60907 );
xor ( n60910 , n59725 , n59770 );
nor ( n60911 , n9662 , n60611 );
and ( n60912 , n60910 , n60911 );
xor ( n60913 , n60910 , n60911 );
xor ( n60914 , n59729 , n59768 );
nor ( n60915 , n9671 , n60611 );
and ( n60916 , n60914 , n60915 );
xor ( n60917 , n60914 , n60915 );
xor ( n60918 , n59733 , n59766 );
nor ( n60919 , n9680 , n60611 );
and ( n60920 , n60918 , n60919 );
xor ( n60921 , n60918 , n60919 );
xor ( n60922 , n59737 , n59764 );
nor ( n60923 , n9689 , n60611 );
and ( n60924 , n60922 , n60923 );
xor ( n60925 , n60922 , n60923 );
xor ( n60926 , n59741 , n59762 );
nor ( n60927 , n9698 , n60611 );
and ( n60928 , n60926 , n60927 );
xor ( n60929 , n60926 , n60927 );
xor ( n60930 , n59745 , n59760 );
nor ( n60931 , n9707 , n60611 );
and ( n60932 , n60930 , n60931 );
xor ( n60933 , n60930 , n60931 );
xor ( n60934 , n59749 , n59758 );
nor ( n60935 , n9716 , n60611 );
and ( n60936 , n60934 , n60935 );
xor ( n60937 , n60934 , n60935 );
xor ( n60938 , n59753 , n59756 );
nor ( n60939 , n9725 , n60611 );
and ( n60940 , n60938 , n60939 );
xor ( n60941 , n60938 , n60939 );
xor ( n60942 , n59754 , n59755 );
nor ( n60943 , n9734 , n60611 );
and ( n60944 , n60942 , n60943 );
xor ( n60945 , n60942 , n60943 );
nor ( n60946 , n9752 , n59423 );
nor ( n60947 , n9743 , n60611 );
and ( n60948 , n60946 , n60947 );
and ( n60949 , n60945 , n60948 );
or ( n60950 , n60944 , n60949 );
and ( n60951 , n60941 , n60950 );
or ( n60952 , n60940 , n60951 );
and ( n60953 , n60937 , n60952 );
or ( n60954 , n60936 , n60953 );
and ( n60955 , n60933 , n60954 );
or ( n60956 , n60932 , n60955 );
and ( n60957 , n60929 , n60956 );
or ( n60958 , n60928 , n60957 );
and ( n60959 , n60925 , n60958 );
or ( n60960 , n60924 , n60959 );
and ( n60961 , n60921 , n60960 );
or ( n60962 , n60920 , n60961 );
and ( n60963 , n60917 , n60962 );
or ( n60964 , n60916 , n60963 );
and ( n60965 , n60913 , n60964 );
or ( n60966 , n60912 , n60965 );
and ( n60967 , n60909 , n60966 );
or ( n60968 , n60908 , n60967 );
and ( n60969 , n60905 , n60968 );
or ( n60970 , n60904 , n60969 );
and ( n60971 , n60901 , n60970 );
or ( n60972 , n60900 , n60971 );
and ( n60973 , n60897 , n60972 );
or ( n60974 , n60896 , n60973 );
and ( n60975 , n60893 , n60974 );
or ( n60976 , n60892 , n60975 );
and ( n60977 , n60889 , n60976 );
or ( n60978 , n60888 , n60977 );
and ( n60979 , n60885 , n60978 );
or ( n60980 , n60884 , n60979 );
and ( n60981 , n60881 , n60980 );
or ( n60982 , n60880 , n60981 );
and ( n60983 , n60877 , n60982 );
or ( n60984 , n60876 , n60983 );
and ( n60985 , n60873 , n60984 );
or ( n60986 , n60872 , n60985 );
and ( n60987 , n60869 , n60986 );
or ( n60988 , n60868 , n60987 );
and ( n60989 , n60865 , n60988 );
or ( n60990 , n60864 , n60989 );
and ( n60991 , n60861 , n60990 );
or ( n60992 , n60860 , n60991 );
and ( n60993 , n60857 , n60992 );
or ( n60994 , n60856 , n60993 );
and ( n60995 , n60853 , n60994 );
or ( n60996 , n60852 , n60995 );
and ( n60997 , n60849 , n60996 );
or ( n60998 , n60848 , n60997 );
and ( n60999 , n60845 , n60998 );
or ( n61000 , n60844 , n60999 );
and ( n61001 , n60841 , n61000 );
or ( n61002 , n60840 , n61001 );
and ( n61003 , n60837 , n61002 );
or ( n61004 , n60836 , n61003 );
and ( n61005 , n60833 , n61004 );
or ( n61006 , n60832 , n61005 );
and ( n61007 , n60829 , n61006 );
or ( n61008 , n60828 , n61007 );
and ( n61009 , n60825 , n61008 );
or ( n61010 , n60824 , n61009 );
and ( n61011 , n60821 , n61010 );
or ( n61012 , n60820 , n61011 );
and ( n61013 , n60817 , n61012 );
or ( n61014 , n60816 , n61013 );
and ( n61015 , n60813 , n61014 );
or ( n61016 , n60812 , n61015 );
and ( n61017 , n60809 , n61016 );
or ( n61018 , n60808 , n61017 );
and ( n61019 , n60805 , n61018 );
or ( n61020 , n60804 , n61019 );
and ( n61021 , n60801 , n61020 );
or ( n61022 , n60800 , n61021 );
and ( n61023 , n60797 , n61022 );
or ( n61024 , n60796 , n61023 );
and ( n61025 , n60793 , n61024 );
or ( n61026 , n60792 , n61025 );
and ( n61027 , n60789 , n61026 );
or ( n61028 , n60788 , n61027 );
and ( n61029 , n60785 , n61028 );
or ( n61030 , n60784 , n61029 );
and ( n61031 , n60781 , n61030 );
or ( n61032 , n60780 , n61031 );
and ( n61033 , n60777 , n61032 );
or ( n61034 , n60776 , n61033 );
and ( n61035 , n60773 , n61034 );
or ( n61036 , n60772 , n61035 );
and ( n61037 , n60769 , n61036 );
or ( n61038 , n60768 , n61037 );
and ( n61039 , n60765 , n61038 );
or ( n61040 , n60764 , n61039 );
and ( n61041 , n60761 , n61040 );
or ( n61042 , n60760 , n61041 );
and ( n61043 , n60757 , n61042 );
or ( n61044 , n60756 , n61043 );
and ( n61045 , n60753 , n61044 );
or ( n61046 , n60752 , n61045 );
and ( n61047 , n60749 , n61046 );
or ( n61048 , n60748 , n61047 );
and ( n61049 , n60745 , n61048 );
or ( n61050 , n60744 , n61049 );
and ( n61051 , n60741 , n61050 );
or ( n61052 , n60740 , n61051 );
and ( n61053 , n60737 , n61052 );
or ( n61054 , n60736 , n61053 );
and ( n61055 , n60733 , n61054 );
or ( n61056 , n60732 , n61055 );
and ( n61057 , n60729 , n61056 );
or ( n61058 , n60728 , n61057 );
and ( n61059 , n60725 , n61058 );
or ( n61060 , n60724 , n61059 );
and ( n61061 , n60721 , n61060 );
or ( n61062 , n60720 , n61061 );
and ( n61063 , n60717 , n61062 );
or ( n61064 , n60716 , n61063 );
and ( n61065 , n60713 , n61064 );
or ( n61066 , n60712 , n61065 );
and ( n61067 , n60709 , n61066 );
or ( n61068 , n60708 , n61067 );
and ( n61069 , n60705 , n61068 );
or ( n61070 , n60704 , n61069 );
and ( n61071 , n60701 , n61070 );
or ( n61072 , n60700 , n61071 );
and ( n61073 , n60697 , n61072 );
or ( n61074 , n60696 , n61073 );
and ( n61075 , n60693 , n61074 );
or ( n61076 , n60692 , n61075 );
and ( n61077 , n60689 , n61076 );
or ( n61078 , n60688 , n61077 );
and ( n61079 , n60685 , n61078 );
or ( n61080 , n60684 , n61079 );
and ( n61081 , n60681 , n61080 );
or ( n61082 , n60680 , n61081 );
and ( n61083 , n60677 , n61082 );
or ( n61084 , n60676 , n61083 );
and ( n61085 , n60673 , n61084 );
or ( n61086 , n60672 , n61085 );
and ( n61087 , n60669 , n61086 );
or ( n61088 , n60668 , n61087 );
and ( n61089 , n60665 , n61088 );
or ( n61090 , n60664 , n61089 );
and ( n61091 , n60661 , n61090 );
or ( n61092 , n60660 , n61091 );
and ( n61093 , n60657 , n61092 );
or ( n61094 , n60656 , n61093 );
and ( n61095 , n60653 , n61094 );
or ( n61096 , n60652 , n61095 );
and ( n61097 , n60649 , n61096 );
or ( n61098 , n60648 , n61097 );
and ( n61099 , n60645 , n61098 );
or ( n61100 , n60644 , n61099 );
and ( n61101 , n60641 , n61100 );
or ( n61102 , n60640 , n61101 );
and ( n61103 , n60637 , n61102 );
or ( n61104 , n60636 , n61103 );
and ( n61105 , n60633 , n61104 );
or ( n61106 , n60632 , n61105 );
and ( n61107 , n60629 , n61106 );
or ( n61108 , n60628 , n61107 );
and ( n61109 , n60625 , n61108 );
or ( n61110 , n60624 , n61109 );
and ( n61111 , n60621 , n61110 );
or ( n61112 , n60620 , n61111 );
and ( n61113 , n60617 , n61112 );
or ( n61114 , n60616 , n61113 );
xor ( n61115 , n60613 , n61114 );
and ( n61116 , n33403 , n3852 );
nor ( n61117 , n3853 , n61116 );
nor ( n61118 , n4151 , n32231 );
xor ( n61119 , n61117 , n61118 );
and ( n61120 , n59923 , n59924 );
and ( n61121 , n59925 , n59928 );
or ( n61122 , n61120 , n61121 );
xor ( n61123 , n61119 , n61122 );
nor ( n61124 , n4458 , n31083 );
xor ( n61125 , n61123 , n61124 );
and ( n61126 , n59929 , n59930 );
and ( n61127 , n59931 , n59934 );
or ( n61128 , n61126 , n61127 );
xor ( n61129 , n61125 , n61128 );
nor ( n61130 , n4786 , n29948 );
xor ( n61131 , n61129 , n61130 );
and ( n61132 , n59935 , n59936 );
and ( n61133 , n59937 , n59940 );
or ( n61134 , n61132 , n61133 );
xor ( n61135 , n61131 , n61134 );
nor ( n61136 , n5126 , n28833 );
xor ( n61137 , n61135 , n61136 );
and ( n61138 , n59941 , n59942 );
and ( n61139 , n59943 , n59946 );
or ( n61140 , n61138 , n61139 );
xor ( n61141 , n61137 , n61140 );
nor ( n61142 , n5477 , n27737 );
xor ( n61143 , n61141 , n61142 );
and ( n61144 , n59947 , n59948 );
and ( n61145 , n59949 , n59952 );
or ( n61146 , n61144 , n61145 );
xor ( n61147 , n61143 , n61146 );
nor ( n61148 , n5838 , n26660 );
xor ( n61149 , n61147 , n61148 );
and ( n61150 , n59953 , n59954 );
and ( n61151 , n59955 , n59958 );
or ( n61152 , n61150 , n61151 );
xor ( n61153 , n61149 , n61152 );
nor ( n61154 , n6212 , n25600 );
xor ( n61155 , n61153 , n61154 );
and ( n61156 , n59959 , n59960 );
and ( n61157 , n59961 , n59964 );
or ( n61158 , n61156 , n61157 );
xor ( n61159 , n61155 , n61158 );
nor ( n61160 , n6596 , n24564 );
xor ( n61161 , n61159 , n61160 );
and ( n61162 , n59965 , n59966 );
and ( n61163 , n59967 , n59970 );
or ( n61164 , n61162 , n61163 );
xor ( n61165 , n61161 , n61164 );
nor ( n61166 , n6997 , n23541 );
xor ( n61167 , n61165 , n61166 );
and ( n61168 , n59971 , n59972 );
and ( n61169 , n59973 , n59976 );
or ( n61170 , n61168 , n61169 );
xor ( n61171 , n61167 , n61170 );
nor ( n61172 , n7413 , n22541 );
xor ( n61173 , n61171 , n61172 );
and ( n61174 , n59977 , n59978 );
and ( n61175 , n59979 , n59982 );
or ( n61176 , n61174 , n61175 );
xor ( n61177 , n61173 , n61176 );
nor ( n61178 , n7841 , n21562 );
xor ( n61179 , n61177 , n61178 );
and ( n61180 , n59983 , n59984 );
and ( n61181 , n59985 , n59988 );
or ( n61182 , n61180 , n61181 );
xor ( n61183 , n61179 , n61182 );
nor ( n61184 , n8281 , n20601 );
xor ( n61185 , n61183 , n61184 );
and ( n61186 , n59989 , n59990 );
and ( n61187 , n59991 , n59994 );
or ( n61188 , n61186 , n61187 );
xor ( n61189 , n61185 , n61188 );
nor ( n61190 , n8737 , n19657 );
xor ( n61191 , n61189 , n61190 );
and ( n61192 , n59995 , n59996 );
and ( n61193 , n59997 , n60000 );
or ( n61194 , n61192 , n61193 );
xor ( n61195 , n61191 , n61194 );
nor ( n61196 , n9420 , n18734 );
xor ( n61197 , n61195 , n61196 );
and ( n61198 , n60001 , n60002 );
and ( n61199 , n60003 , n60006 );
or ( n61200 , n61198 , n61199 );
xor ( n61201 , n61197 , n61200 );
nor ( n61202 , n10312 , n17828 );
xor ( n61203 , n61201 , n61202 );
and ( n61204 , n60007 , n60008 );
and ( n61205 , n60009 , n60012 );
or ( n61206 , n61204 , n61205 );
xor ( n61207 , n61203 , n61206 );
nor ( n61208 , n11041 , n16943 );
xor ( n61209 , n61207 , n61208 );
and ( n61210 , n60013 , n60014 );
and ( n61211 , n60015 , n60018 );
or ( n61212 , n61210 , n61211 );
xor ( n61213 , n61209 , n61212 );
nor ( n61214 , n11790 , n16077 );
xor ( n61215 , n61213 , n61214 );
and ( n61216 , n60019 , n60020 );
and ( n61217 , n60021 , n60024 );
or ( n61218 , n61216 , n61217 );
xor ( n61219 , n61215 , n61218 );
nor ( n61220 , n12555 , n15230 );
xor ( n61221 , n61219 , n61220 );
and ( n61222 , n60025 , n60026 );
and ( n61223 , n60027 , n60030 );
or ( n61224 , n61222 , n61223 );
xor ( n61225 , n61221 , n61224 );
nor ( n61226 , n13340 , n14403 );
xor ( n61227 , n61225 , n61226 );
and ( n61228 , n60031 , n60032 );
and ( n61229 , n60033 , n60036 );
or ( n61230 , n61228 , n61229 );
xor ( n61231 , n61227 , n61230 );
nor ( n61232 , n14138 , n13599 );
xor ( n61233 , n61231 , n61232 );
and ( n61234 , n60037 , n60038 );
and ( n61235 , n60039 , n60042 );
or ( n61236 , n61234 , n61235 );
xor ( n61237 , n61233 , n61236 );
nor ( n61238 , n14959 , n12808 );
xor ( n61239 , n61237 , n61238 );
and ( n61240 , n60043 , n60044 );
and ( n61241 , n60045 , n60048 );
or ( n61242 , n61240 , n61241 );
xor ( n61243 , n61239 , n61242 );
nor ( n61244 , n15800 , n12037 );
xor ( n61245 , n61243 , n61244 );
and ( n61246 , n60049 , n60050 );
and ( n61247 , n60051 , n60054 );
or ( n61248 , n61246 , n61247 );
xor ( n61249 , n61245 , n61248 );
nor ( n61250 , n16660 , n11282 );
xor ( n61251 , n61249 , n61250 );
and ( n61252 , n60055 , n60056 );
and ( n61253 , n60057 , n60060 );
or ( n61254 , n61252 , n61253 );
xor ( n61255 , n61251 , n61254 );
nor ( n61256 , n17539 , n10547 );
xor ( n61257 , n61255 , n61256 );
and ( n61258 , n60061 , n60062 );
and ( n61259 , n60063 , n60066 );
or ( n61260 , n61258 , n61259 );
xor ( n61261 , n61257 , n61260 );
nor ( n61262 , n18439 , n9829 );
xor ( n61263 , n61261 , n61262 );
and ( n61264 , n60067 , n60068 );
and ( n61265 , n60069 , n60072 );
or ( n61266 , n61264 , n61265 );
xor ( n61267 , n61263 , n61266 );
nor ( n61268 , n19356 , n8955 );
xor ( n61269 , n61267 , n61268 );
and ( n61270 , n60073 , n60074 );
and ( n61271 , n60075 , n60078 );
or ( n61272 , n61270 , n61271 );
xor ( n61273 , n61269 , n61272 );
nor ( n61274 , n20294 , n603 );
xor ( n61275 , n61273 , n61274 );
and ( n61276 , n60079 , n60080 );
and ( n61277 , n60081 , n60084 );
or ( n61278 , n61276 , n61277 );
xor ( n61279 , n61275 , n61278 );
nor ( n61280 , n21249 , n652 );
xor ( n61281 , n61279 , n61280 );
and ( n61282 , n60085 , n60086 );
and ( n61283 , n60087 , n60090 );
or ( n61284 , n61282 , n61283 );
xor ( n61285 , n61281 , n61284 );
nor ( n61286 , n22222 , n624 );
xor ( n61287 , n61285 , n61286 );
and ( n61288 , n60091 , n60092 );
and ( n61289 , n60093 , n60096 );
or ( n61290 , n61288 , n61289 );
xor ( n61291 , n61287 , n61290 );
nor ( n61292 , n23216 , n648 );
xor ( n61293 , n61291 , n61292 );
and ( n61294 , n60097 , n60098 );
and ( n61295 , n60099 , n60102 );
or ( n61296 , n61294 , n61295 );
xor ( n61297 , n61293 , n61296 );
nor ( n61298 , n24233 , n686 );
xor ( n61299 , n61297 , n61298 );
and ( n61300 , n60103 , n60104 );
and ( n61301 , n60105 , n60108 );
or ( n61302 , n61300 , n61301 );
xor ( n61303 , n61299 , n61302 );
nor ( n61304 , n25263 , n735 );
xor ( n61305 , n61303 , n61304 );
and ( n61306 , n60109 , n60110 );
and ( n61307 , n60111 , n60114 );
or ( n61308 , n61306 , n61307 );
xor ( n61309 , n61305 , n61308 );
nor ( n61310 , n26317 , n798 );
xor ( n61311 , n61309 , n61310 );
and ( n61312 , n60115 , n60116 );
and ( n61313 , n60117 , n60120 );
or ( n61314 , n61312 , n61313 );
xor ( n61315 , n61311 , n61314 );
nor ( n61316 , n27388 , n870 );
xor ( n61317 , n61315 , n61316 );
and ( n61318 , n60121 , n60122 );
and ( n61319 , n60123 , n60126 );
or ( n61320 , n61318 , n61319 );
xor ( n61321 , n61317 , n61320 );
nor ( n61322 , n28478 , n960 );
xor ( n61323 , n61321 , n61322 );
and ( n61324 , n60127 , n60128 );
and ( n61325 , n60129 , n60132 );
or ( n61326 , n61324 , n61325 );
xor ( n61327 , n61323 , n61326 );
nor ( n61328 , n29587 , n1064 );
xor ( n61329 , n61327 , n61328 );
and ( n61330 , n60133 , n60134 );
and ( n61331 , n60135 , n60138 );
or ( n61332 , n61330 , n61331 );
xor ( n61333 , n61329 , n61332 );
nor ( n61334 , n30716 , n1178 );
xor ( n61335 , n61333 , n61334 );
and ( n61336 , n60139 , n60140 );
and ( n61337 , n60141 , n60144 );
or ( n61338 , n61336 , n61337 );
xor ( n61339 , n61335 , n61338 );
nor ( n61340 , n31858 , n1305 );
xor ( n61341 , n61339 , n61340 );
and ( n61342 , n60145 , n60146 );
and ( n61343 , n60147 , n60150 );
or ( n61344 , n61342 , n61343 );
xor ( n61345 , n61341 , n61344 );
nor ( n61346 , n33024 , n1447 );
xor ( n61347 , n61345 , n61346 );
and ( n61348 , n60151 , n60152 );
and ( n61349 , n60153 , n60156 );
or ( n61350 , n61348 , n61349 );
xor ( n61351 , n61347 , n61350 );
nor ( n61352 , n34215 , n1600 );
xor ( n61353 , n61351 , n61352 );
and ( n61354 , n60157 , n60158 );
and ( n61355 , n60159 , n60162 );
or ( n61356 , n61354 , n61355 );
xor ( n61357 , n61353 , n61356 );
nor ( n61358 , n35410 , n1768 );
xor ( n61359 , n61357 , n61358 );
and ( n61360 , n60163 , n60164 );
and ( n61361 , n60165 , n60168 );
or ( n61362 , n61360 , n61361 );
xor ( n61363 , n61359 , n61362 );
nor ( n61364 , n36611 , n1947 );
xor ( n61365 , n61363 , n61364 );
and ( n61366 , n60169 , n60170 );
and ( n61367 , n60171 , n60174 );
or ( n61368 , n61366 , n61367 );
xor ( n61369 , n61365 , n61368 );
nor ( n61370 , n37816 , n2139 );
xor ( n61371 , n61369 , n61370 );
and ( n61372 , n60175 , n60176 );
and ( n61373 , n60177 , n60180 );
or ( n61374 , n61372 , n61373 );
xor ( n61375 , n61371 , n61374 );
nor ( n61376 , n39018 , n2345 );
xor ( n61377 , n61375 , n61376 );
and ( n61378 , n60181 , n60182 );
and ( n61379 , n60183 , n60186 );
or ( n61380 , n61378 , n61379 );
xor ( n61381 , n61377 , n61380 );
nor ( n61382 , n40223 , n2568 );
xor ( n61383 , n61381 , n61382 );
and ( n61384 , n60187 , n60188 );
and ( n61385 , n60189 , n60192 );
or ( n61386 , n61384 , n61385 );
xor ( n61387 , n61383 , n61386 );
nor ( n61388 , n41428 , n2799 );
xor ( n61389 , n61387 , n61388 );
and ( n61390 , n60193 , n60194 );
and ( n61391 , n60195 , n60198 );
or ( n61392 , n61390 , n61391 );
xor ( n61393 , n61389 , n61392 );
nor ( n61394 , n42632 , n3045 );
xor ( n61395 , n61393 , n61394 );
and ( n61396 , n60199 , n60200 );
and ( n61397 , n60201 , n60204 );
or ( n61398 , n61396 , n61397 );
xor ( n61399 , n61395 , n61398 );
nor ( n61400 , n43834 , n3302 );
xor ( n61401 , n61399 , n61400 );
and ( n61402 , n60205 , n60206 );
and ( n61403 , n60207 , n60210 );
or ( n61404 , n61402 , n61403 );
xor ( n61405 , n61401 , n61404 );
nor ( n61406 , n45038 , n3572 );
xor ( n61407 , n61405 , n61406 );
and ( n61408 , n60211 , n60212 );
and ( n61409 , n60213 , n60216 );
or ( n61410 , n61408 , n61409 );
xor ( n61411 , n61407 , n61410 );
nor ( n61412 , n46239 , n3855 );
xor ( n61413 , n61411 , n61412 );
and ( n61414 , n60217 , n60218 );
and ( n61415 , n60219 , n60222 );
or ( n61416 , n61414 , n61415 );
xor ( n61417 , n61413 , n61416 );
nor ( n61418 , n47440 , n4153 );
xor ( n61419 , n61417 , n61418 );
and ( n61420 , n60223 , n60224 );
and ( n61421 , n60225 , n60228 );
or ( n61422 , n61420 , n61421 );
xor ( n61423 , n61419 , n61422 );
nor ( n61424 , n48641 , n4460 );
xor ( n61425 , n61423 , n61424 );
and ( n61426 , n60229 , n60230 );
and ( n61427 , n60231 , n60234 );
or ( n61428 , n61426 , n61427 );
xor ( n61429 , n61425 , n61428 );
nor ( n61430 , n49841 , n4788 );
xor ( n61431 , n61429 , n61430 );
and ( n61432 , n60235 , n60236 );
and ( n61433 , n60237 , n60240 );
or ( n61434 , n61432 , n61433 );
xor ( n61435 , n61431 , n61434 );
nor ( n61436 , n51040 , n5128 );
xor ( n61437 , n61435 , n61436 );
and ( n61438 , n60241 , n60242 );
and ( n61439 , n60243 , n60246 );
or ( n61440 , n61438 , n61439 );
xor ( n61441 , n61437 , n61440 );
nor ( n61442 , n52238 , n5479 );
xor ( n61443 , n61441 , n61442 );
and ( n61444 , n60247 , n60248 );
and ( n61445 , n60249 , n60252 );
or ( n61446 , n61444 , n61445 );
xor ( n61447 , n61443 , n61446 );
nor ( n61448 , n53432 , n5840 );
xor ( n61449 , n61447 , n61448 );
and ( n61450 , n60253 , n60254 );
and ( n61451 , n60255 , n60258 );
or ( n61452 , n61450 , n61451 );
xor ( n61453 , n61449 , n61452 );
nor ( n61454 , n54629 , n6214 );
xor ( n61455 , n61453 , n61454 );
and ( n61456 , n60259 , n60260 );
and ( n61457 , n60261 , n60264 );
or ( n61458 , n61456 , n61457 );
xor ( n61459 , n61455 , n61458 );
nor ( n61460 , n55826 , n6598 );
xor ( n61461 , n61459 , n61460 );
and ( n61462 , n60265 , n60266 );
and ( n61463 , n60267 , n60270 );
or ( n61464 , n61462 , n61463 );
xor ( n61465 , n61461 , n61464 );
nor ( n61466 , n57022 , n6999 );
xor ( n61467 , n61465 , n61466 );
and ( n61468 , n60271 , n60272 );
and ( n61469 , n60273 , n60276 );
or ( n61470 , n61468 , n61469 );
xor ( n61471 , n61467 , n61470 );
nor ( n61472 , n58217 , n7415 );
xor ( n61473 , n61471 , n61472 );
and ( n61474 , n60277 , n60278 );
and ( n61475 , n60279 , n60282 );
or ( n61476 , n61474 , n61475 );
xor ( n61477 , n61473 , n61476 );
nor ( n61478 , n59412 , n7843 );
xor ( n61479 , n61477 , n61478 );
and ( n61480 , n60283 , n60284 );
and ( n61481 , n60285 , n60288 );
or ( n61482 , n61480 , n61481 );
xor ( n61483 , n61479 , n61482 );
nor ( n61484 , n60600 , n8283 );
xor ( n61485 , n61483 , n61484 );
and ( n61486 , n60289 , n60290 );
and ( n61487 , n60291 , n60294 );
or ( n61488 , n61486 , n61487 );
xor ( n61489 , n61485 , n61488 );
and ( n61490 , n60307 , n60311 );
and ( n61491 , n60311 , n60586 );
and ( n61492 , n60307 , n60586 );
or ( n61493 , n61490 , n61491 , n61492 );
and ( n61494 , n33774 , n3749 );
not ( n61495 , n3749 );
nor ( n61496 , n61494 , n61495 );
xor ( n61497 , n61493 , n61496 );
and ( n61498 , n60320 , n60324 );
and ( n61499 , n60324 , n60392 );
and ( n61500 , n60320 , n60392 );
or ( n61501 , n61498 , n61499 , n61500 );
and ( n61502 , n60316 , n60393 );
and ( n61503 , n60393 , n60585 );
and ( n61504 , n60316 , n60585 );
or ( n61505 , n61502 , n61503 , n61504 );
xor ( n61506 , n61501 , n61505 );
and ( n61507 , n60395 , n60509 );
and ( n61508 , n60509 , n60584 );
and ( n61509 , n60395 , n60584 );
or ( n61510 , n61507 , n61508 , n61509 );
and ( n61511 , n60329 , n60333 );
and ( n61512 , n60333 , n60391 );
and ( n61513 , n60329 , n60391 );
or ( n61514 , n61511 , n61512 , n61513 );
and ( n61515 , n60399 , n60400 );
and ( n61516 , n60400 , n60508 );
and ( n61517 , n60399 , n60508 );
or ( n61518 , n61515 , n61516 , n61517 );
xor ( n61519 , n61514 , n61518 );
and ( n61520 , n60360 , n60364 );
and ( n61521 , n60364 , n60370 );
and ( n61522 , n60360 , n60370 );
or ( n61523 , n61520 , n61521 , n61522 );
and ( n61524 , n60338 , n60342 );
and ( n61525 , n60342 , n60390 );
and ( n61526 , n60338 , n60390 );
or ( n61527 , n61524 , n61525 , n61526 );
xor ( n61528 , n61523 , n61527 );
and ( n61529 , n60347 , n60351 );
and ( n61530 , n60351 , n60389 );
and ( n61531 , n60347 , n60389 );
or ( n61532 , n61529 , n61530 , n61531 );
and ( n61533 , n60409 , n60434 );
and ( n61534 , n60434 , n60469 );
and ( n61535 , n60409 , n60469 );
or ( n61536 , n61533 , n61534 , n61535 );
xor ( n61537 , n61532 , n61536 );
and ( n61538 , n60356 , n60371 );
and ( n61539 , n60371 , n60388 );
and ( n61540 , n60356 , n60388 );
or ( n61541 , n61538 , n61539 , n61540 );
and ( n61542 , n60413 , n60417 );
and ( n61543 , n60417 , n60433 );
and ( n61544 , n60413 , n60433 );
or ( n61545 , n61542 , n61543 , n61544 );
xor ( n61546 , n61541 , n61545 );
and ( n61547 , n60376 , n60381 );
and ( n61548 , n60381 , n60387 );
and ( n61549 , n60376 , n60387 );
or ( n61550 , n61547 , n61548 , n61549 );
and ( n61551 , n60366 , n60367 );
and ( n61552 , n60367 , n60369 );
and ( n61553 , n60366 , n60369 );
or ( n61554 , n61551 , n61552 , n61553 );
and ( n61555 , n60377 , n60378 );
and ( n61556 , n60378 , n60380 );
and ( n61557 , n60377 , n60380 );
or ( n61558 , n61555 , n61556 , n61557 );
xor ( n61559 , n61554 , n61558 );
and ( n61560 , n30695 , n4730 );
and ( n61561 , n31836 , n4403 );
xor ( n61562 , n61560 , n61561 );
and ( n61563 , n32649 , n4102 );
xor ( n61564 , n61562 , n61563 );
xor ( n61565 , n61559 , n61564 );
xor ( n61566 , n61550 , n61565 );
and ( n61567 , n60383 , n60384 );
and ( n61568 , n60384 , n60386 );
and ( n61569 , n60383 , n60386 );
or ( n61570 , n61567 , n61568 , n61569 );
and ( n61571 , n27361 , n5765 );
and ( n61572 , n28456 , n5408 );
xor ( n61573 , n61571 , n61572 );
and ( n61574 , n29559 , n5103 );
xor ( n61575 , n61573 , n61574 );
xor ( n61576 , n61570 , n61575 );
and ( n61577 , n24214 , n6971 );
and ( n61578 , n25243 , n6504 );
xor ( n61579 , n61577 , n61578 );
and ( n61580 , n26296 , n6132 );
xor ( n61581 , n61579 , n61580 );
xor ( n61582 , n61576 , n61581 );
xor ( n61583 , n61566 , n61582 );
xor ( n61584 , n61546 , n61583 );
xor ( n61585 , n61537 , n61584 );
xor ( n61586 , n61528 , n61585 );
xor ( n61587 , n61519 , n61586 );
xor ( n61588 , n61510 , n61587 );
and ( n61589 , n60515 , n60583 );
and ( n61590 , n60405 , n60470 );
and ( n61591 , n60470 , n60507 );
and ( n61592 , n60405 , n60507 );
or ( n61593 , n61590 , n61591 , n61592 );
and ( n61594 , n60519 , n60582 );
xor ( n61595 , n61593 , n61594 );
and ( n61596 , n60475 , n60479 );
and ( n61597 , n60479 , n60506 );
and ( n61598 , n60475 , n60506 );
or ( n61599 , n61596 , n61597 , n61598 );
and ( n61600 , n60439 , n60455 );
and ( n61601 , n60455 , n60468 );
and ( n61602 , n60439 , n60468 );
or ( n61603 , n61600 , n61601 , n61602 );
and ( n61604 , n60422 , n60426 );
and ( n61605 , n60426 , n60432 );
and ( n61606 , n60422 , n60432 );
or ( n61607 , n61604 , n61605 , n61606 );
and ( n61608 , n60443 , n60448 );
and ( n61609 , n60448 , n60454 );
and ( n61610 , n60443 , n60454 );
or ( n61611 , n61608 , n61609 , n61610 );
xor ( n61612 , n61607 , n61611 );
and ( n61613 , n60428 , n60429 );
and ( n61614 , n60429 , n60431 );
and ( n61615 , n60428 , n60431 );
or ( n61616 , n61613 , n61614 , n61615 );
and ( n61617 , n60444 , n60445 );
and ( n61618 , n60445 , n60447 );
and ( n61619 , n60444 , n60447 );
or ( n61620 , n61617 , n61618 , n61619 );
xor ( n61621 , n61616 , n61620 );
and ( n61622 , n21216 , n8243 );
and ( n61623 , n22186 , n7662 );
xor ( n61624 , n61622 , n61623 );
and ( n61625 , n22892 , n7310 );
xor ( n61626 , n61624 , n61625 );
xor ( n61627 , n61621 , n61626 );
xor ( n61628 , n61612 , n61627 );
xor ( n61629 , n61603 , n61628 );
and ( n61630 , n60460 , n60464 );
and ( n61631 , n60464 , n60467 );
and ( n61632 , n60460 , n60467 );
or ( n61633 , n61630 , n61631 , n61632 );
and ( n61634 , n60450 , n60451 );
and ( n61635 , n60451 , n60453 );
and ( n61636 , n60450 , n60453 );
or ( n61637 , n61634 , n61635 , n61636 );
and ( n61638 , n18144 , n10239 );
and ( n61639 , n19324 , n9348 );
xor ( n61640 , n61638 , n61639 );
and ( n61641 , n20233 , n8669 );
xor ( n61642 , n61640 , n61641 );
xor ( n61643 , n61637 , n61642 );
and ( n61644 , n15758 , n12531 );
and ( n61645 , n16637 , n11718 );
xor ( n61646 , n61644 , n61645 );
and ( n61647 , n17512 , n10977 );
xor ( n61648 , n61646 , n61647 );
xor ( n61649 , n61643 , n61648 );
xor ( n61650 , n61633 , n61649 );
and ( n61651 , n13322 , n14044 );
and ( n61652 , n14118 , n13256 );
and ( n61653 , n61651 , n61652 );
and ( n61654 , n61652 , n60466 );
and ( n61655 , n61651 , n60466 );
or ( n61656 , n61653 , n61654 , n61655 );
and ( n61657 , n60494 , n60495 );
and ( n61658 , n60495 , n60497 );
and ( n61659 , n60494 , n60497 );
or ( n61660 , n61657 , n61658 , n61659 );
xor ( n61661 , n61656 , n61660 );
and ( n61662 , n13322 , n14838 );
buf ( n61663 , n14118 );
xor ( n61664 , n61662 , n61663 );
and ( n61665 , n14938 , n13256 );
xor ( n61666 , n61664 , n61665 );
xor ( n61667 , n61661 , n61666 );
xor ( n61668 , n61650 , n61667 );
xor ( n61669 , n61629 , n61668 );
xor ( n61670 , n61599 , n61669 );
and ( n61671 , n60484 , n60488 );
and ( n61672 , n60488 , n60505 );
and ( n61673 , n60484 , n60505 );
or ( n61674 , n61671 , n61672 , n61673 );
and ( n61675 , n60527 , n60542 );
and ( n61676 , n60542 , n60559 );
and ( n61677 , n60527 , n60559 );
or ( n61678 , n61675 , n61676 , n61677 );
xor ( n61679 , n61674 , n61678 );
and ( n61680 , n60493 , n60498 );
and ( n61681 , n60498 , n60504 );
and ( n61682 , n60493 , n60504 );
or ( n61683 , n61680 , n61681 , n61682 );
and ( n61684 , n60531 , n60535 );
and ( n61685 , n60535 , n60541 );
and ( n61686 , n60531 , n60541 );
or ( n61687 , n61684 , n61685 , n61686 );
xor ( n61688 , n61683 , n61687 );
and ( n61689 , n60500 , n60501 );
and ( n61690 , n60501 , n60503 );
and ( n61691 , n60500 , n60503 );
or ( n61692 , n61689 , n61690 , n61691 );
and ( n61693 , n11015 , n17422 );
and ( n61694 , n11769 , n16550 );
xor ( n61695 , n61693 , n61694 );
and ( n61696 , n12320 , n15691 );
xor ( n61697 , n61695 , n61696 );
xor ( n61698 , n61692 , n61697 );
and ( n61699 , n8718 , n20156 );
and ( n61700 , n9400 , n19222 );
xor ( n61701 , n61699 , n61700 );
and ( n61702 , n10291 , n18407 );
xor ( n61703 , n61701 , n61702 );
xor ( n61704 , n61698 , n61703 );
xor ( n61705 , n61688 , n61704 );
xor ( n61706 , n61679 , n61705 );
xor ( n61707 , n61670 , n61706 );
xor ( n61708 , n61595 , n61707 );
xor ( n61709 , n61589 , n61708 );
not ( n61710 , n3801 );
and ( n61711 , n34193 , n3801 );
nor ( n61712 , n61710 , n61711 );
and ( n61713 , n60523 , n60560 );
and ( n61714 , n60560 , n60581 );
and ( n61715 , n60523 , n60581 );
or ( n61716 , n61713 , n61714 , n61715 );
and ( n61717 , n60565 , n60580 );
and ( n61718 , n60547 , n60552 );
and ( n61719 , n60552 , n60558 );
and ( n61720 , n60547 , n60558 );
or ( n61721 , n61718 , n61719 , n61720 );
and ( n61722 , n60537 , n60538 );
and ( n61723 , n60538 , n60540 );
and ( n61724 , n60537 , n60540 );
or ( n61725 , n61722 , n61723 , n61724 );
and ( n61726 , n60548 , n60549 );
and ( n61727 , n60549 , n60551 );
and ( n61728 , n60548 , n60551 );
or ( n61729 , n61726 , n61727 , n61728 );
xor ( n61730 , n61725 , n61729 );
and ( n61731 , n7385 , n23075 );
and ( n61732 , n7808 , n22065 );
xor ( n61733 , n61731 , n61732 );
and ( n61734 , n8079 , n20976 );
xor ( n61735 , n61733 , n61734 );
xor ( n61736 , n61730 , n61735 );
xor ( n61737 , n61721 , n61736 );
and ( n61738 , n60554 , n60555 );
and ( n61739 , n60555 , n60557 );
and ( n61740 , n60554 , n60557 );
or ( n61741 , n61738 , n61739 , n61740 );
and ( n61742 , n6187 , n26216 );
and ( n61743 , n6569 , n25163 );
xor ( n61744 , n61742 , n61743 );
and ( n61745 , n6816 , n24137 );
xor ( n61746 , n61744 , n61745 );
xor ( n61747 , n61741 , n61746 );
and ( n61748 , n4959 , n29508 );
and ( n61749 , n5459 , n28406 );
xor ( n61750 , n61748 , n61749 );
and ( n61751 , n5819 , n27296 );
xor ( n61752 , n61750 , n61751 );
xor ( n61753 , n61747 , n61752 );
xor ( n61754 , n61737 , n61753 );
xor ( n61755 , n61717 , n61754 );
and ( n61756 , n60569 , n60573 );
and ( n61757 , n60573 , n60579 );
and ( n61758 , n60569 , n60579 );
or ( n61759 , n61756 , n61757 , n61758 );
and ( n61760 , n60575 , n60576 );
and ( n61761 , n60576 , n60578 );
and ( n61762 , n60575 , n60578 );
or ( n61763 , n61760 , n61761 , n61762 );
and ( n61764 , n60513 , n60514 );
xor ( n61765 , n61763 , n61764 );
and ( n61766 , n4132 , n32999 );
and ( n61767 , n4438 , n31761 );
xor ( n61768 , n61766 , n61767 );
and ( n61769 , n4766 , n30629 );
xor ( n61770 , n61768 , n61769 );
xor ( n61771 , n61765 , n61770 );
xor ( n61772 , n61759 , n61771 );
xor ( n61773 , n61755 , n61772 );
xor ( n61774 , n61716 , n61773 );
xor ( n61775 , n61712 , n61774 );
xor ( n61776 , n61709 , n61775 );
xor ( n61777 , n61588 , n61776 );
xor ( n61778 , n61506 , n61777 );
xor ( n61779 , n61497 , n61778 );
and ( n61780 , n60299 , n60302 );
and ( n61781 , n60302 , n60587 );
and ( n61782 , n60299 , n60587 );
or ( n61783 , n61780 , n61781 , n61782 );
xor ( n61784 , n61779 , n61783 );
and ( n61785 , n60588 , n60592 );
and ( n61786 , n60593 , n60596 );
or ( n61787 , n61785 , n61786 );
xor ( n61788 , n61784 , n61787 );
buf ( n61789 , n61788 );
buf ( n61790 , n61789 );
not ( n61791 , n61790 );
nor ( n61792 , n61791 , n8739 );
xor ( n61793 , n61489 , n61792 );
and ( n61794 , n60295 , n60601 );
and ( n61795 , n60602 , n60605 );
or ( n61796 , n61794 , n61795 );
xor ( n61797 , n61793 , n61796 );
buf ( n61798 , n61797 );
buf ( n61799 , n61798 );
not ( n61800 , n61799 );
buf ( n61801 , n585 );
not ( n61802 , n61801 );
nor ( n61803 , n61800 , n61802 );
xor ( n61804 , n61115 , n61803 );
xor ( n61805 , n60617 , n61112 );
nor ( n61806 , n60609 , n61802 );
and ( n61807 , n61805 , n61806 );
xor ( n61808 , n61805 , n61806 );
xor ( n61809 , n60621 , n61110 );
nor ( n61810 , n59421 , n61802 );
and ( n61811 , n61809 , n61810 );
xor ( n61812 , n61809 , n61810 );
xor ( n61813 , n60625 , n61108 );
nor ( n61814 , n58226 , n61802 );
and ( n61815 , n61813 , n61814 );
xor ( n61816 , n61813 , n61814 );
xor ( n61817 , n60629 , n61106 );
nor ( n61818 , n57031 , n61802 );
and ( n61819 , n61817 , n61818 );
xor ( n61820 , n61817 , n61818 );
xor ( n61821 , n60633 , n61104 );
nor ( n61822 , n55835 , n61802 );
and ( n61823 , n61821 , n61822 );
xor ( n61824 , n61821 , n61822 );
xor ( n61825 , n60637 , n61102 );
nor ( n61826 , n54638 , n61802 );
and ( n61827 , n61825 , n61826 );
xor ( n61828 , n61825 , n61826 );
xor ( n61829 , n60641 , n61100 );
nor ( n61830 , n53441 , n61802 );
and ( n61831 , n61829 , n61830 );
xor ( n61832 , n61829 , n61830 );
xor ( n61833 , n60645 , n61098 );
nor ( n61834 , n52247 , n61802 );
and ( n61835 , n61833 , n61834 );
xor ( n61836 , n61833 , n61834 );
xor ( n61837 , n60649 , n61096 );
nor ( n61838 , n51049 , n61802 );
and ( n61839 , n61837 , n61838 );
xor ( n61840 , n61837 , n61838 );
xor ( n61841 , n60653 , n61094 );
nor ( n61842 , n49850 , n61802 );
and ( n61843 , n61841 , n61842 );
xor ( n61844 , n61841 , n61842 );
xor ( n61845 , n60657 , n61092 );
nor ( n61846 , n48650 , n61802 );
and ( n61847 , n61845 , n61846 );
xor ( n61848 , n61845 , n61846 );
xor ( n61849 , n60661 , n61090 );
nor ( n61850 , n47449 , n61802 );
and ( n61851 , n61849 , n61850 );
xor ( n61852 , n61849 , n61850 );
xor ( n61853 , n60665 , n61088 );
nor ( n61854 , n46248 , n61802 );
and ( n61855 , n61853 , n61854 );
xor ( n61856 , n61853 , n61854 );
xor ( n61857 , n60669 , n61086 );
nor ( n61858 , n45047 , n61802 );
and ( n61859 , n61857 , n61858 );
xor ( n61860 , n61857 , n61858 );
xor ( n61861 , n60673 , n61084 );
nor ( n61862 , n43843 , n61802 );
and ( n61863 , n61861 , n61862 );
xor ( n61864 , n61861 , n61862 );
xor ( n61865 , n60677 , n61082 );
nor ( n61866 , n42641 , n61802 );
and ( n61867 , n61865 , n61866 );
xor ( n61868 , n61865 , n61866 );
xor ( n61869 , n60681 , n61080 );
nor ( n61870 , n41437 , n61802 );
and ( n61871 , n61869 , n61870 );
xor ( n61872 , n61869 , n61870 );
xor ( n61873 , n60685 , n61078 );
nor ( n61874 , n40232 , n61802 );
and ( n61875 , n61873 , n61874 );
xor ( n61876 , n61873 , n61874 );
xor ( n61877 , n60689 , n61076 );
nor ( n61878 , n39027 , n61802 );
and ( n61879 , n61877 , n61878 );
xor ( n61880 , n61877 , n61878 );
xor ( n61881 , n60693 , n61074 );
nor ( n61882 , n37825 , n61802 );
and ( n61883 , n61881 , n61882 );
xor ( n61884 , n61881 , n61882 );
xor ( n61885 , n60697 , n61072 );
nor ( n61886 , n36620 , n61802 );
and ( n61887 , n61885 , n61886 );
xor ( n61888 , n61885 , n61886 );
xor ( n61889 , n60701 , n61070 );
nor ( n61890 , n35419 , n61802 );
and ( n61891 , n61889 , n61890 );
xor ( n61892 , n61889 , n61890 );
xor ( n61893 , n60705 , n61068 );
nor ( n61894 , n34224 , n61802 );
and ( n61895 , n61893 , n61894 );
xor ( n61896 , n61893 , n61894 );
xor ( n61897 , n60709 , n61066 );
nor ( n61898 , n33033 , n61802 );
and ( n61899 , n61897 , n61898 );
xor ( n61900 , n61897 , n61898 );
xor ( n61901 , n60713 , n61064 );
nor ( n61902 , n31867 , n61802 );
and ( n61903 , n61901 , n61902 );
xor ( n61904 , n61901 , n61902 );
xor ( n61905 , n60717 , n61062 );
nor ( n61906 , n30725 , n61802 );
and ( n61907 , n61905 , n61906 );
xor ( n61908 , n61905 , n61906 );
xor ( n61909 , n60721 , n61060 );
nor ( n61910 , n29596 , n61802 );
and ( n61911 , n61909 , n61910 );
xor ( n61912 , n61909 , n61910 );
xor ( n61913 , n60725 , n61058 );
nor ( n61914 , n28487 , n61802 );
and ( n61915 , n61913 , n61914 );
xor ( n61916 , n61913 , n61914 );
xor ( n61917 , n60729 , n61056 );
nor ( n61918 , n27397 , n61802 );
and ( n61919 , n61917 , n61918 );
xor ( n61920 , n61917 , n61918 );
xor ( n61921 , n60733 , n61054 );
nor ( n61922 , n26326 , n61802 );
and ( n61923 , n61921 , n61922 );
xor ( n61924 , n61921 , n61922 );
xor ( n61925 , n60737 , n61052 );
nor ( n61926 , n25272 , n61802 );
and ( n61927 , n61925 , n61926 );
xor ( n61928 , n61925 , n61926 );
xor ( n61929 , n60741 , n61050 );
nor ( n61930 , n24242 , n61802 );
and ( n61931 , n61929 , n61930 );
xor ( n61932 , n61929 , n61930 );
xor ( n61933 , n60745 , n61048 );
nor ( n61934 , n23225 , n61802 );
and ( n61935 , n61933 , n61934 );
xor ( n61936 , n61933 , n61934 );
xor ( n61937 , n60749 , n61046 );
nor ( n61938 , n22231 , n61802 );
and ( n61939 , n61937 , n61938 );
xor ( n61940 , n61937 , n61938 );
xor ( n61941 , n60753 , n61044 );
nor ( n61942 , n21258 , n61802 );
and ( n61943 , n61941 , n61942 );
xor ( n61944 , n61941 , n61942 );
xor ( n61945 , n60757 , n61042 );
nor ( n61946 , n20303 , n61802 );
and ( n61947 , n61945 , n61946 );
xor ( n61948 , n61945 , n61946 );
xor ( n61949 , n60761 , n61040 );
nor ( n61950 , n19365 , n61802 );
and ( n61951 , n61949 , n61950 );
xor ( n61952 , n61949 , n61950 );
xor ( n61953 , n60765 , n61038 );
nor ( n61954 , n18448 , n61802 );
and ( n61955 , n61953 , n61954 );
xor ( n61956 , n61953 , n61954 );
xor ( n61957 , n60769 , n61036 );
nor ( n61958 , n17548 , n61802 );
and ( n61959 , n61957 , n61958 );
xor ( n61960 , n61957 , n61958 );
xor ( n61961 , n60773 , n61034 );
nor ( n61962 , n16669 , n61802 );
and ( n61963 , n61961 , n61962 );
xor ( n61964 , n61961 , n61962 );
xor ( n61965 , n60777 , n61032 );
nor ( n61966 , n15809 , n61802 );
and ( n61967 , n61965 , n61966 );
xor ( n61968 , n61965 , n61966 );
xor ( n61969 , n60781 , n61030 );
nor ( n61970 , n14968 , n61802 );
and ( n61971 , n61969 , n61970 );
xor ( n61972 , n61969 , n61970 );
xor ( n61973 , n60785 , n61028 );
nor ( n61974 , n14147 , n61802 );
and ( n61975 , n61973 , n61974 );
xor ( n61976 , n61973 , n61974 );
xor ( n61977 , n60789 , n61026 );
nor ( n61978 , n13349 , n61802 );
and ( n61979 , n61977 , n61978 );
xor ( n61980 , n61977 , n61978 );
xor ( n61981 , n60793 , n61024 );
nor ( n61982 , n12564 , n61802 );
and ( n61983 , n61981 , n61982 );
xor ( n61984 , n61981 , n61982 );
xor ( n61985 , n60797 , n61022 );
nor ( n61986 , n11799 , n61802 );
and ( n61987 , n61985 , n61986 );
xor ( n61988 , n61985 , n61986 );
xor ( n61989 , n60801 , n61020 );
nor ( n61990 , n11050 , n61802 );
and ( n61991 , n61989 , n61990 );
xor ( n61992 , n61989 , n61990 );
xor ( n61993 , n60805 , n61018 );
nor ( n61994 , n10321 , n61802 );
and ( n61995 , n61993 , n61994 );
xor ( n61996 , n61993 , n61994 );
xor ( n61997 , n60809 , n61016 );
nor ( n61998 , n9429 , n61802 );
and ( n61999 , n61997 , n61998 );
xor ( n62000 , n61997 , n61998 );
xor ( n62001 , n60813 , n61014 );
nor ( n62002 , n8949 , n61802 );
and ( n62003 , n62001 , n62002 );
xor ( n62004 , n62001 , n62002 );
xor ( n62005 , n60817 , n61012 );
nor ( n62006 , n9437 , n61802 );
and ( n62007 , n62005 , n62006 );
xor ( n62008 , n62005 , n62006 );
xor ( n62009 , n60821 , n61010 );
nor ( n62010 , n9446 , n61802 );
and ( n62011 , n62009 , n62010 );
xor ( n62012 , n62009 , n62010 );
xor ( n62013 , n60825 , n61008 );
nor ( n62014 , n9455 , n61802 );
and ( n62015 , n62013 , n62014 );
xor ( n62016 , n62013 , n62014 );
xor ( n62017 , n60829 , n61006 );
nor ( n62018 , n9464 , n61802 );
and ( n62019 , n62017 , n62018 );
xor ( n62020 , n62017 , n62018 );
xor ( n62021 , n60833 , n61004 );
nor ( n62022 , n9473 , n61802 );
and ( n62023 , n62021 , n62022 );
xor ( n62024 , n62021 , n62022 );
xor ( n62025 , n60837 , n61002 );
nor ( n62026 , n9482 , n61802 );
and ( n62027 , n62025 , n62026 );
xor ( n62028 , n62025 , n62026 );
xor ( n62029 , n60841 , n61000 );
nor ( n62030 , n9491 , n61802 );
and ( n62031 , n62029 , n62030 );
xor ( n62032 , n62029 , n62030 );
xor ( n62033 , n60845 , n60998 );
nor ( n62034 , n9500 , n61802 );
and ( n62035 , n62033 , n62034 );
xor ( n62036 , n62033 , n62034 );
xor ( n62037 , n60849 , n60996 );
nor ( n62038 , n9509 , n61802 );
and ( n62039 , n62037 , n62038 );
xor ( n62040 , n62037 , n62038 );
xor ( n62041 , n60853 , n60994 );
nor ( n62042 , n9518 , n61802 );
and ( n62043 , n62041 , n62042 );
xor ( n62044 , n62041 , n62042 );
xor ( n62045 , n60857 , n60992 );
nor ( n62046 , n9527 , n61802 );
and ( n62047 , n62045 , n62046 );
xor ( n62048 , n62045 , n62046 );
xor ( n62049 , n60861 , n60990 );
nor ( n62050 , n9536 , n61802 );
and ( n62051 , n62049 , n62050 );
xor ( n62052 , n62049 , n62050 );
xor ( n62053 , n60865 , n60988 );
nor ( n62054 , n9545 , n61802 );
and ( n62055 , n62053 , n62054 );
xor ( n62056 , n62053 , n62054 );
xor ( n62057 , n60869 , n60986 );
nor ( n62058 , n9554 , n61802 );
and ( n62059 , n62057 , n62058 );
xor ( n62060 , n62057 , n62058 );
xor ( n62061 , n60873 , n60984 );
nor ( n62062 , n9563 , n61802 );
and ( n62063 , n62061 , n62062 );
xor ( n62064 , n62061 , n62062 );
xor ( n62065 , n60877 , n60982 );
nor ( n62066 , n9572 , n61802 );
and ( n62067 , n62065 , n62066 );
xor ( n62068 , n62065 , n62066 );
xor ( n62069 , n60881 , n60980 );
nor ( n62070 , n9581 , n61802 );
and ( n62071 , n62069 , n62070 );
xor ( n62072 , n62069 , n62070 );
xor ( n62073 , n60885 , n60978 );
nor ( n62074 , n9590 , n61802 );
and ( n62075 , n62073 , n62074 );
xor ( n62076 , n62073 , n62074 );
xor ( n62077 , n60889 , n60976 );
nor ( n62078 , n9599 , n61802 );
and ( n62079 , n62077 , n62078 );
xor ( n62080 , n62077 , n62078 );
xor ( n62081 , n60893 , n60974 );
nor ( n62082 , n9608 , n61802 );
and ( n62083 , n62081 , n62082 );
xor ( n62084 , n62081 , n62082 );
xor ( n62085 , n60897 , n60972 );
nor ( n62086 , n9617 , n61802 );
and ( n62087 , n62085 , n62086 );
xor ( n62088 , n62085 , n62086 );
xor ( n62089 , n60901 , n60970 );
nor ( n62090 , n9626 , n61802 );
and ( n62091 , n62089 , n62090 );
xor ( n62092 , n62089 , n62090 );
xor ( n62093 , n60905 , n60968 );
nor ( n62094 , n9635 , n61802 );
and ( n62095 , n62093 , n62094 );
xor ( n62096 , n62093 , n62094 );
xor ( n62097 , n60909 , n60966 );
nor ( n62098 , n9644 , n61802 );
and ( n62099 , n62097 , n62098 );
xor ( n62100 , n62097 , n62098 );
xor ( n62101 , n60913 , n60964 );
nor ( n62102 , n9653 , n61802 );
and ( n62103 , n62101 , n62102 );
xor ( n62104 , n62101 , n62102 );
xor ( n62105 , n60917 , n60962 );
nor ( n62106 , n9662 , n61802 );
and ( n62107 , n62105 , n62106 );
xor ( n62108 , n62105 , n62106 );
xor ( n62109 , n60921 , n60960 );
nor ( n62110 , n9671 , n61802 );
and ( n62111 , n62109 , n62110 );
xor ( n62112 , n62109 , n62110 );
xor ( n62113 , n60925 , n60958 );
nor ( n62114 , n9680 , n61802 );
and ( n62115 , n62113 , n62114 );
xor ( n62116 , n62113 , n62114 );
xor ( n62117 , n60929 , n60956 );
nor ( n62118 , n9689 , n61802 );
and ( n62119 , n62117 , n62118 );
xor ( n62120 , n62117 , n62118 );
xor ( n62121 , n60933 , n60954 );
nor ( n62122 , n9698 , n61802 );
and ( n62123 , n62121 , n62122 );
xor ( n62124 , n62121 , n62122 );
xor ( n62125 , n60937 , n60952 );
nor ( n62126 , n9707 , n61802 );
and ( n62127 , n62125 , n62126 );
xor ( n62128 , n62125 , n62126 );
xor ( n62129 , n60941 , n60950 );
nor ( n62130 , n9716 , n61802 );
and ( n62131 , n62129 , n62130 );
xor ( n62132 , n62129 , n62130 );
xor ( n62133 , n60945 , n60948 );
nor ( n62134 , n9725 , n61802 );
and ( n62135 , n62133 , n62134 );
xor ( n62136 , n62133 , n62134 );
xor ( n62137 , n60946 , n60947 );
nor ( n62138 , n9734 , n61802 );
and ( n62139 , n62137 , n62138 );
xor ( n62140 , n62137 , n62138 );
nor ( n62141 , n9752 , n60611 );
nor ( n62142 , n9743 , n61802 );
and ( n62143 , n62141 , n62142 );
and ( n62144 , n62140 , n62143 );
or ( n62145 , n62139 , n62144 );
and ( n62146 , n62136 , n62145 );
or ( n62147 , n62135 , n62146 );
and ( n62148 , n62132 , n62147 );
or ( n62149 , n62131 , n62148 );
and ( n62150 , n62128 , n62149 );
or ( n62151 , n62127 , n62150 );
and ( n62152 , n62124 , n62151 );
or ( n62153 , n62123 , n62152 );
and ( n62154 , n62120 , n62153 );
or ( n62155 , n62119 , n62154 );
and ( n62156 , n62116 , n62155 );
or ( n62157 , n62115 , n62156 );
and ( n62158 , n62112 , n62157 );
or ( n62159 , n62111 , n62158 );
and ( n62160 , n62108 , n62159 );
or ( n62161 , n62107 , n62160 );
and ( n62162 , n62104 , n62161 );
or ( n62163 , n62103 , n62162 );
and ( n62164 , n62100 , n62163 );
or ( n62165 , n62099 , n62164 );
and ( n62166 , n62096 , n62165 );
or ( n62167 , n62095 , n62166 );
and ( n62168 , n62092 , n62167 );
or ( n62169 , n62091 , n62168 );
and ( n62170 , n62088 , n62169 );
or ( n62171 , n62087 , n62170 );
and ( n62172 , n62084 , n62171 );
or ( n62173 , n62083 , n62172 );
and ( n62174 , n62080 , n62173 );
or ( n62175 , n62079 , n62174 );
and ( n62176 , n62076 , n62175 );
or ( n62177 , n62075 , n62176 );
and ( n62178 , n62072 , n62177 );
or ( n62179 , n62071 , n62178 );
and ( n62180 , n62068 , n62179 );
or ( n62181 , n62067 , n62180 );
and ( n62182 , n62064 , n62181 );
or ( n62183 , n62063 , n62182 );
and ( n62184 , n62060 , n62183 );
or ( n62185 , n62059 , n62184 );
and ( n62186 , n62056 , n62185 );
or ( n62187 , n62055 , n62186 );
and ( n62188 , n62052 , n62187 );
or ( n62189 , n62051 , n62188 );
and ( n62190 , n62048 , n62189 );
or ( n62191 , n62047 , n62190 );
and ( n62192 , n62044 , n62191 );
or ( n62193 , n62043 , n62192 );
and ( n62194 , n62040 , n62193 );
or ( n62195 , n62039 , n62194 );
and ( n62196 , n62036 , n62195 );
or ( n62197 , n62035 , n62196 );
and ( n62198 , n62032 , n62197 );
or ( n62199 , n62031 , n62198 );
and ( n62200 , n62028 , n62199 );
or ( n62201 , n62027 , n62200 );
and ( n62202 , n62024 , n62201 );
or ( n62203 , n62023 , n62202 );
and ( n62204 , n62020 , n62203 );
or ( n62205 , n62019 , n62204 );
and ( n62206 , n62016 , n62205 );
or ( n62207 , n62015 , n62206 );
and ( n62208 , n62012 , n62207 );
or ( n62209 , n62011 , n62208 );
and ( n62210 , n62008 , n62209 );
or ( n62211 , n62007 , n62210 );
and ( n62212 , n62004 , n62211 );
or ( n62213 , n62003 , n62212 );
and ( n62214 , n62000 , n62213 );
or ( n62215 , n61999 , n62214 );
and ( n62216 , n61996 , n62215 );
or ( n62217 , n61995 , n62216 );
and ( n62218 , n61992 , n62217 );
or ( n62219 , n61991 , n62218 );
and ( n62220 , n61988 , n62219 );
or ( n62221 , n61987 , n62220 );
and ( n62222 , n61984 , n62221 );
or ( n62223 , n61983 , n62222 );
and ( n62224 , n61980 , n62223 );
or ( n62225 , n61979 , n62224 );
and ( n62226 , n61976 , n62225 );
or ( n62227 , n61975 , n62226 );
and ( n62228 , n61972 , n62227 );
or ( n62229 , n61971 , n62228 );
and ( n62230 , n61968 , n62229 );
or ( n62231 , n61967 , n62230 );
and ( n62232 , n61964 , n62231 );
or ( n62233 , n61963 , n62232 );
and ( n62234 , n61960 , n62233 );
or ( n62235 , n61959 , n62234 );
and ( n62236 , n61956 , n62235 );
or ( n62237 , n61955 , n62236 );
and ( n62238 , n61952 , n62237 );
or ( n62239 , n61951 , n62238 );
and ( n62240 , n61948 , n62239 );
or ( n62241 , n61947 , n62240 );
and ( n62242 , n61944 , n62241 );
or ( n62243 , n61943 , n62242 );
and ( n62244 , n61940 , n62243 );
or ( n62245 , n61939 , n62244 );
and ( n62246 , n61936 , n62245 );
or ( n62247 , n61935 , n62246 );
and ( n62248 , n61932 , n62247 );
or ( n62249 , n61931 , n62248 );
and ( n62250 , n61928 , n62249 );
or ( n62251 , n61927 , n62250 );
and ( n62252 , n61924 , n62251 );
or ( n62253 , n61923 , n62252 );
and ( n62254 , n61920 , n62253 );
or ( n62255 , n61919 , n62254 );
and ( n62256 , n61916 , n62255 );
or ( n62257 , n61915 , n62256 );
and ( n62258 , n61912 , n62257 );
or ( n62259 , n61911 , n62258 );
and ( n62260 , n61908 , n62259 );
or ( n62261 , n61907 , n62260 );
and ( n62262 , n61904 , n62261 );
or ( n62263 , n61903 , n62262 );
and ( n62264 , n61900 , n62263 );
or ( n62265 , n61899 , n62264 );
and ( n62266 , n61896 , n62265 );
or ( n62267 , n61895 , n62266 );
and ( n62268 , n61892 , n62267 );
or ( n62269 , n61891 , n62268 );
and ( n62270 , n61888 , n62269 );
or ( n62271 , n61887 , n62270 );
and ( n62272 , n61884 , n62271 );
or ( n62273 , n61883 , n62272 );
and ( n62274 , n61880 , n62273 );
or ( n62275 , n61879 , n62274 );
and ( n62276 , n61876 , n62275 );
or ( n62277 , n61875 , n62276 );
and ( n62278 , n61872 , n62277 );
or ( n62279 , n61871 , n62278 );
and ( n62280 , n61868 , n62279 );
or ( n62281 , n61867 , n62280 );
and ( n62282 , n61864 , n62281 );
or ( n62283 , n61863 , n62282 );
and ( n62284 , n61860 , n62283 );
or ( n62285 , n61859 , n62284 );
and ( n62286 , n61856 , n62285 );
or ( n62287 , n61855 , n62286 );
and ( n62288 , n61852 , n62287 );
or ( n62289 , n61851 , n62288 );
and ( n62290 , n61848 , n62289 );
or ( n62291 , n61847 , n62290 );
and ( n62292 , n61844 , n62291 );
or ( n62293 , n61843 , n62292 );
and ( n62294 , n61840 , n62293 );
or ( n62295 , n61839 , n62294 );
and ( n62296 , n61836 , n62295 );
or ( n62297 , n61835 , n62296 );
and ( n62298 , n61832 , n62297 );
or ( n62299 , n61831 , n62298 );
and ( n62300 , n61828 , n62299 );
or ( n62301 , n61827 , n62300 );
and ( n62302 , n61824 , n62301 );
or ( n62303 , n61823 , n62302 );
and ( n62304 , n61820 , n62303 );
or ( n62305 , n61819 , n62304 );
and ( n62306 , n61816 , n62305 );
or ( n62307 , n61815 , n62306 );
and ( n62308 , n61812 , n62307 );
or ( n62309 , n61811 , n62308 );
and ( n62310 , n61808 , n62309 );
or ( n62311 , n61807 , n62310 );
xor ( n62312 , n61804 , n62311 );
and ( n62313 , n33403 , n4150 );
nor ( n62314 , n4151 , n62313 );
nor ( n62315 , n4458 , n32231 );
xor ( n62316 , n62314 , n62315 );
and ( n62317 , n61117 , n61118 );
and ( n62318 , n61119 , n61122 );
or ( n62319 , n62317 , n62318 );
xor ( n62320 , n62316 , n62319 );
nor ( n62321 , n4786 , n31083 );
xor ( n62322 , n62320 , n62321 );
and ( n62323 , n61123 , n61124 );
and ( n62324 , n61125 , n61128 );
or ( n62325 , n62323 , n62324 );
xor ( n62326 , n62322 , n62325 );
nor ( n62327 , n5126 , n29948 );
xor ( n62328 , n62326 , n62327 );
and ( n62329 , n61129 , n61130 );
and ( n62330 , n61131 , n61134 );
or ( n62331 , n62329 , n62330 );
xor ( n62332 , n62328 , n62331 );
nor ( n62333 , n5477 , n28833 );
xor ( n62334 , n62332 , n62333 );
and ( n62335 , n61135 , n61136 );
and ( n62336 , n61137 , n61140 );
or ( n62337 , n62335 , n62336 );
xor ( n62338 , n62334 , n62337 );
nor ( n62339 , n5838 , n27737 );
xor ( n62340 , n62338 , n62339 );
and ( n62341 , n61141 , n61142 );
and ( n62342 , n61143 , n61146 );
or ( n62343 , n62341 , n62342 );
xor ( n62344 , n62340 , n62343 );
nor ( n62345 , n6212 , n26660 );
xor ( n62346 , n62344 , n62345 );
and ( n62347 , n61147 , n61148 );
and ( n62348 , n61149 , n61152 );
or ( n62349 , n62347 , n62348 );
xor ( n62350 , n62346 , n62349 );
nor ( n62351 , n6596 , n25600 );
xor ( n62352 , n62350 , n62351 );
and ( n62353 , n61153 , n61154 );
and ( n62354 , n61155 , n61158 );
or ( n62355 , n62353 , n62354 );
xor ( n62356 , n62352 , n62355 );
nor ( n62357 , n6997 , n24564 );
xor ( n62358 , n62356 , n62357 );
and ( n62359 , n61159 , n61160 );
and ( n62360 , n61161 , n61164 );
or ( n62361 , n62359 , n62360 );
xor ( n62362 , n62358 , n62361 );
nor ( n62363 , n7413 , n23541 );
xor ( n62364 , n62362 , n62363 );
and ( n62365 , n61165 , n61166 );
and ( n62366 , n61167 , n61170 );
or ( n62367 , n62365 , n62366 );
xor ( n62368 , n62364 , n62367 );
nor ( n62369 , n7841 , n22541 );
xor ( n62370 , n62368 , n62369 );
and ( n62371 , n61171 , n61172 );
and ( n62372 , n61173 , n61176 );
or ( n62373 , n62371 , n62372 );
xor ( n62374 , n62370 , n62373 );
nor ( n62375 , n8281 , n21562 );
xor ( n62376 , n62374 , n62375 );
and ( n62377 , n61177 , n61178 );
and ( n62378 , n61179 , n61182 );
or ( n62379 , n62377 , n62378 );
xor ( n62380 , n62376 , n62379 );
nor ( n62381 , n8737 , n20601 );
xor ( n62382 , n62380 , n62381 );
and ( n62383 , n61183 , n61184 );
and ( n62384 , n61185 , n61188 );
or ( n62385 , n62383 , n62384 );
xor ( n62386 , n62382 , n62385 );
nor ( n62387 , n9420 , n19657 );
xor ( n62388 , n62386 , n62387 );
and ( n62389 , n61189 , n61190 );
and ( n62390 , n61191 , n61194 );
or ( n62391 , n62389 , n62390 );
xor ( n62392 , n62388 , n62391 );
nor ( n62393 , n10312 , n18734 );
xor ( n62394 , n62392 , n62393 );
and ( n62395 , n61195 , n61196 );
and ( n62396 , n61197 , n61200 );
or ( n62397 , n62395 , n62396 );
xor ( n62398 , n62394 , n62397 );
nor ( n62399 , n11041 , n17828 );
xor ( n62400 , n62398 , n62399 );
and ( n62401 , n61201 , n61202 );
and ( n62402 , n61203 , n61206 );
or ( n62403 , n62401 , n62402 );
xor ( n62404 , n62400 , n62403 );
nor ( n62405 , n11790 , n16943 );
xor ( n62406 , n62404 , n62405 );
and ( n62407 , n61207 , n61208 );
and ( n62408 , n61209 , n61212 );
or ( n62409 , n62407 , n62408 );
xor ( n62410 , n62406 , n62409 );
nor ( n62411 , n12555 , n16077 );
xor ( n62412 , n62410 , n62411 );
and ( n62413 , n61213 , n61214 );
and ( n62414 , n61215 , n61218 );
or ( n62415 , n62413 , n62414 );
xor ( n62416 , n62412 , n62415 );
nor ( n62417 , n13340 , n15230 );
xor ( n62418 , n62416 , n62417 );
and ( n62419 , n61219 , n61220 );
and ( n62420 , n61221 , n61224 );
or ( n62421 , n62419 , n62420 );
xor ( n62422 , n62418 , n62421 );
nor ( n62423 , n14138 , n14403 );
xor ( n62424 , n62422 , n62423 );
and ( n62425 , n61225 , n61226 );
and ( n62426 , n61227 , n61230 );
or ( n62427 , n62425 , n62426 );
xor ( n62428 , n62424 , n62427 );
nor ( n62429 , n14959 , n13599 );
xor ( n62430 , n62428 , n62429 );
and ( n62431 , n61231 , n61232 );
and ( n62432 , n61233 , n61236 );
or ( n62433 , n62431 , n62432 );
xor ( n62434 , n62430 , n62433 );
nor ( n62435 , n15800 , n12808 );
xor ( n62436 , n62434 , n62435 );
and ( n62437 , n61237 , n61238 );
and ( n62438 , n61239 , n61242 );
or ( n62439 , n62437 , n62438 );
xor ( n62440 , n62436 , n62439 );
nor ( n62441 , n16660 , n12037 );
xor ( n62442 , n62440 , n62441 );
and ( n62443 , n61243 , n61244 );
and ( n62444 , n61245 , n61248 );
or ( n62445 , n62443 , n62444 );
xor ( n62446 , n62442 , n62445 );
nor ( n62447 , n17539 , n11282 );
xor ( n62448 , n62446 , n62447 );
and ( n62449 , n61249 , n61250 );
and ( n62450 , n61251 , n61254 );
or ( n62451 , n62449 , n62450 );
xor ( n62452 , n62448 , n62451 );
nor ( n62453 , n18439 , n10547 );
xor ( n62454 , n62452 , n62453 );
and ( n62455 , n61255 , n61256 );
and ( n62456 , n61257 , n61260 );
or ( n62457 , n62455 , n62456 );
xor ( n62458 , n62454 , n62457 );
nor ( n62459 , n19356 , n9829 );
xor ( n62460 , n62458 , n62459 );
and ( n62461 , n61261 , n61262 );
and ( n62462 , n61263 , n61266 );
or ( n62463 , n62461 , n62462 );
xor ( n62464 , n62460 , n62463 );
nor ( n62465 , n20294 , n8955 );
xor ( n62466 , n62464 , n62465 );
and ( n62467 , n61267 , n61268 );
and ( n62468 , n61269 , n61272 );
or ( n62469 , n62467 , n62468 );
xor ( n62470 , n62466 , n62469 );
nor ( n62471 , n21249 , n603 );
xor ( n62472 , n62470 , n62471 );
and ( n62473 , n61273 , n61274 );
and ( n62474 , n61275 , n61278 );
or ( n62475 , n62473 , n62474 );
xor ( n62476 , n62472 , n62475 );
nor ( n62477 , n22222 , n652 );
xor ( n62478 , n62476 , n62477 );
and ( n62479 , n61279 , n61280 );
and ( n62480 , n61281 , n61284 );
or ( n62481 , n62479 , n62480 );
xor ( n62482 , n62478 , n62481 );
nor ( n62483 , n23216 , n624 );
xor ( n62484 , n62482 , n62483 );
and ( n62485 , n61285 , n61286 );
and ( n62486 , n61287 , n61290 );
or ( n62487 , n62485 , n62486 );
xor ( n62488 , n62484 , n62487 );
nor ( n62489 , n24233 , n648 );
xor ( n62490 , n62488 , n62489 );
and ( n62491 , n61291 , n61292 );
and ( n62492 , n61293 , n61296 );
or ( n62493 , n62491 , n62492 );
xor ( n62494 , n62490 , n62493 );
nor ( n62495 , n25263 , n686 );
xor ( n62496 , n62494 , n62495 );
and ( n62497 , n61297 , n61298 );
and ( n62498 , n61299 , n61302 );
or ( n62499 , n62497 , n62498 );
xor ( n62500 , n62496 , n62499 );
nor ( n62501 , n26317 , n735 );
xor ( n62502 , n62500 , n62501 );
and ( n62503 , n61303 , n61304 );
and ( n62504 , n61305 , n61308 );
or ( n62505 , n62503 , n62504 );
xor ( n62506 , n62502 , n62505 );
nor ( n62507 , n27388 , n798 );
xor ( n62508 , n62506 , n62507 );
and ( n62509 , n61309 , n61310 );
and ( n62510 , n61311 , n61314 );
or ( n62511 , n62509 , n62510 );
xor ( n62512 , n62508 , n62511 );
nor ( n62513 , n28478 , n870 );
xor ( n62514 , n62512 , n62513 );
and ( n62515 , n61315 , n61316 );
and ( n62516 , n61317 , n61320 );
or ( n62517 , n62515 , n62516 );
xor ( n62518 , n62514 , n62517 );
nor ( n62519 , n29587 , n960 );
xor ( n62520 , n62518 , n62519 );
and ( n62521 , n61321 , n61322 );
and ( n62522 , n61323 , n61326 );
or ( n62523 , n62521 , n62522 );
xor ( n62524 , n62520 , n62523 );
nor ( n62525 , n30716 , n1064 );
xor ( n62526 , n62524 , n62525 );
and ( n62527 , n61327 , n61328 );
and ( n62528 , n61329 , n61332 );
or ( n62529 , n62527 , n62528 );
xor ( n62530 , n62526 , n62529 );
nor ( n62531 , n31858 , n1178 );
xor ( n62532 , n62530 , n62531 );
and ( n62533 , n61333 , n61334 );
and ( n62534 , n61335 , n61338 );
or ( n62535 , n62533 , n62534 );
xor ( n62536 , n62532 , n62535 );
nor ( n62537 , n33024 , n1305 );
xor ( n62538 , n62536 , n62537 );
and ( n62539 , n61339 , n61340 );
and ( n62540 , n61341 , n61344 );
or ( n62541 , n62539 , n62540 );
xor ( n62542 , n62538 , n62541 );
nor ( n62543 , n34215 , n1447 );
xor ( n62544 , n62542 , n62543 );
and ( n62545 , n61345 , n61346 );
and ( n62546 , n61347 , n61350 );
or ( n62547 , n62545 , n62546 );
xor ( n62548 , n62544 , n62547 );
nor ( n62549 , n35410 , n1600 );
xor ( n62550 , n62548 , n62549 );
and ( n62551 , n61351 , n61352 );
and ( n62552 , n61353 , n61356 );
or ( n62553 , n62551 , n62552 );
xor ( n62554 , n62550 , n62553 );
nor ( n62555 , n36611 , n1768 );
xor ( n62556 , n62554 , n62555 );
and ( n62557 , n61357 , n61358 );
and ( n62558 , n61359 , n61362 );
or ( n62559 , n62557 , n62558 );
xor ( n62560 , n62556 , n62559 );
nor ( n62561 , n37816 , n1947 );
xor ( n62562 , n62560 , n62561 );
and ( n62563 , n61363 , n61364 );
and ( n62564 , n61365 , n61368 );
or ( n62565 , n62563 , n62564 );
xor ( n62566 , n62562 , n62565 );
nor ( n62567 , n39018 , n2139 );
xor ( n62568 , n62566 , n62567 );
and ( n62569 , n61369 , n61370 );
and ( n62570 , n61371 , n61374 );
or ( n62571 , n62569 , n62570 );
xor ( n62572 , n62568 , n62571 );
nor ( n62573 , n40223 , n2345 );
xor ( n62574 , n62572 , n62573 );
and ( n62575 , n61375 , n61376 );
and ( n62576 , n61377 , n61380 );
or ( n62577 , n62575 , n62576 );
xor ( n62578 , n62574 , n62577 );
nor ( n62579 , n41428 , n2568 );
xor ( n62580 , n62578 , n62579 );
and ( n62581 , n61381 , n61382 );
and ( n62582 , n61383 , n61386 );
or ( n62583 , n62581 , n62582 );
xor ( n62584 , n62580 , n62583 );
nor ( n62585 , n42632 , n2799 );
xor ( n62586 , n62584 , n62585 );
and ( n62587 , n61387 , n61388 );
and ( n62588 , n61389 , n61392 );
or ( n62589 , n62587 , n62588 );
xor ( n62590 , n62586 , n62589 );
nor ( n62591 , n43834 , n3045 );
xor ( n62592 , n62590 , n62591 );
and ( n62593 , n61393 , n61394 );
and ( n62594 , n61395 , n61398 );
or ( n62595 , n62593 , n62594 );
xor ( n62596 , n62592 , n62595 );
nor ( n62597 , n45038 , n3302 );
xor ( n62598 , n62596 , n62597 );
and ( n62599 , n61399 , n61400 );
and ( n62600 , n61401 , n61404 );
or ( n62601 , n62599 , n62600 );
xor ( n62602 , n62598 , n62601 );
nor ( n62603 , n46239 , n3572 );
xor ( n62604 , n62602 , n62603 );
and ( n62605 , n61405 , n61406 );
and ( n62606 , n61407 , n61410 );
or ( n62607 , n62605 , n62606 );
xor ( n62608 , n62604 , n62607 );
nor ( n62609 , n47440 , n3855 );
xor ( n62610 , n62608 , n62609 );
and ( n62611 , n61411 , n61412 );
and ( n62612 , n61413 , n61416 );
or ( n62613 , n62611 , n62612 );
xor ( n62614 , n62610 , n62613 );
nor ( n62615 , n48641 , n4153 );
xor ( n62616 , n62614 , n62615 );
and ( n62617 , n61417 , n61418 );
and ( n62618 , n61419 , n61422 );
or ( n62619 , n62617 , n62618 );
xor ( n62620 , n62616 , n62619 );
nor ( n62621 , n49841 , n4460 );
xor ( n62622 , n62620 , n62621 );
and ( n62623 , n61423 , n61424 );
and ( n62624 , n61425 , n61428 );
or ( n62625 , n62623 , n62624 );
xor ( n62626 , n62622 , n62625 );
nor ( n62627 , n51040 , n4788 );
xor ( n62628 , n62626 , n62627 );
and ( n62629 , n61429 , n61430 );
and ( n62630 , n61431 , n61434 );
or ( n62631 , n62629 , n62630 );
xor ( n62632 , n62628 , n62631 );
nor ( n62633 , n52238 , n5128 );
xor ( n62634 , n62632 , n62633 );
and ( n62635 , n61435 , n61436 );
and ( n62636 , n61437 , n61440 );
or ( n62637 , n62635 , n62636 );
xor ( n62638 , n62634 , n62637 );
nor ( n62639 , n53432 , n5479 );
xor ( n62640 , n62638 , n62639 );
and ( n62641 , n61441 , n61442 );
and ( n62642 , n61443 , n61446 );
or ( n62643 , n62641 , n62642 );
xor ( n62644 , n62640 , n62643 );
nor ( n62645 , n54629 , n5840 );
xor ( n62646 , n62644 , n62645 );
and ( n62647 , n61447 , n61448 );
and ( n62648 , n61449 , n61452 );
or ( n62649 , n62647 , n62648 );
xor ( n62650 , n62646 , n62649 );
nor ( n62651 , n55826 , n6214 );
xor ( n62652 , n62650 , n62651 );
and ( n62653 , n61453 , n61454 );
and ( n62654 , n61455 , n61458 );
or ( n62655 , n62653 , n62654 );
xor ( n62656 , n62652 , n62655 );
nor ( n62657 , n57022 , n6598 );
xor ( n62658 , n62656 , n62657 );
and ( n62659 , n61459 , n61460 );
and ( n62660 , n61461 , n61464 );
or ( n62661 , n62659 , n62660 );
xor ( n62662 , n62658 , n62661 );
nor ( n62663 , n58217 , n6999 );
xor ( n62664 , n62662 , n62663 );
and ( n62665 , n61465 , n61466 );
and ( n62666 , n61467 , n61470 );
or ( n62667 , n62665 , n62666 );
xor ( n62668 , n62664 , n62667 );
nor ( n62669 , n59412 , n7415 );
xor ( n62670 , n62668 , n62669 );
and ( n62671 , n61471 , n61472 );
and ( n62672 , n61473 , n61476 );
or ( n62673 , n62671 , n62672 );
xor ( n62674 , n62670 , n62673 );
nor ( n62675 , n60600 , n7843 );
xor ( n62676 , n62674 , n62675 );
and ( n62677 , n61477 , n61478 );
and ( n62678 , n61479 , n61482 );
or ( n62679 , n62677 , n62678 );
xor ( n62680 , n62676 , n62679 );
nor ( n62681 , n61791 , n8283 );
xor ( n62682 , n62680 , n62681 );
and ( n62683 , n61483 , n61484 );
and ( n62684 , n61485 , n61488 );
or ( n62685 , n62683 , n62684 );
xor ( n62686 , n62682 , n62685 );
and ( n62687 , n61501 , n61505 );
and ( n62688 , n61505 , n61777 );
and ( n62689 , n61501 , n61777 );
or ( n62690 , n62687 , n62688 , n62689 );
and ( n62691 , n33774 , n4102 );
not ( n62692 , n4102 );
nor ( n62693 , n62691 , n62692 );
xor ( n62694 , n62690 , n62693 );
and ( n62695 , n61514 , n61518 );
and ( n62696 , n61518 , n61586 );
and ( n62697 , n61514 , n61586 );
or ( n62698 , n62695 , n62696 , n62697 );
and ( n62699 , n61510 , n61587 );
and ( n62700 , n61587 , n61776 );
and ( n62701 , n61510 , n61776 );
or ( n62702 , n62699 , n62700 , n62701 );
xor ( n62703 , n62698 , n62702 );
and ( n62704 , n61589 , n61708 );
and ( n62705 , n61708 , n61775 );
and ( n62706 , n61589 , n61775 );
or ( n62707 , n62704 , n62705 , n62706 );
and ( n62708 , n61523 , n61527 );
and ( n62709 , n61527 , n61585 );
and ( n62710 , n61523 , n61585 );
or ( n62711 , n62708 , n62709 , n62710 );
and ( n62712 , n61593 , n61594 );
and ( n62713 , n61594 , n61707 );
and ( n62714 , n61593 , n61707 );
or ( n62715 , n62712 , n62713 , n62714 );
xor ( n62716 , n62711 , n62715 );
and ( n62717 , n61554 , n61558 );
and ( n62718 , n61558 , n61564 );
and ( n62719 , n61554 , n61564 );
or ( n62720 , n62717 , n62718 , n62719 );
and ( n62721 , n61532 , n61536 );
and ( n62722 , n61536 , n61584 );
and ( n62723 , n61532 , n61584 );
or ( n62724 , n62721 , n62722 , n62723 );
xor ( n62725 , n62720 , n62724 );
and ( n62726 , n61541 , n61545 );
and ( n62727 , n61545 , n61583 );
and ( n62728 , n61541 , n61583 );
or ( n62729 , n62726 , n62727 , n62728 );
and ( n62730 , n61603 , n61628 );
and ( n62731 , n61628 , n61668 );
and ( n62732 , n61603 , n61668 );
or ( n62733 , n62730 , n62731 , n62732 );
xor ( n62734 , n62729 , n62733 );
and ( n62735 , n61550 , n61565 );
and ( n62736 , n61565 , n61582 );
and ( n62737 , n61550 , n61582 );
or ( n62738 , n62735 , n62736 , n62737 );
and ( n62739 , n61607 , n61611 );
and ( n62740 , n61611 , n61627 );
and ( n62741 , n61607 , n61627 );
or ( n62742 , n62739 , n62740 , n62741 );
xor ( n62743 , n62738 , n62742 );
and ( n62744 , n61570 , n61575 );
and ( n62745 , n61575 , n61581 );
and ( n62746 , n61570 , n61581 );
or ( n62747 , n62744 , n62745 , n62746 );
and ( n62748 , n61560 , n61561 );
and ( n62749 , n61561 , n61563 );
and ( n62750 , n61560 , n61563 );
or ( n62751 , n62748 , n62749 , n62750 );
and ( n62752 , n61571 , n61572 );
and ( n62753 , n61572 , n61574 );
and ( n62754 , n61571 , n61574 );
or ( n62755 , n62752 , n62753 , n62754 );
xor ( n62756 , n62751 , n62755 );
and ( n62757 , n30695 , n5103 );
and ( n62758 , n31836 , n4730 );
xor ( n62759 , n62757 , n62758 );
and ( n62760 , n32649 , n4403 );
xor ( n62761 , n62759 , n62760 );
xor ( n62762 , n62756 , n62761 );
xor ( n62763 , n62747 , n62762 );
and ( n62764 , n61577 , n61578 );
and ( n62765 , n61578 , n61580 );
and ( n62766 , n61577 , n61580 );
or ( n62767 , n62764 , n62765 , n62766 );
and ( n62768 , n27361 , n6132 );
and ( n62769 , n28456 , n5765 );
xor ( n62770 , n62768 , n62769 );
and ( n62771 , n29559 , n5408 );
xor ( n62772 , n62770 , n62771 );
xor ( n62773 , n62767 , n62772 );
and ( n62774 , n24214 , n7310 );
and ( n62775 , n25243 , n6971 );
xor ( n62776 , n62774 , n62775 );
and ( n62777 , n26296 , n6504 );
xor ( n62778 , n62776 , n62777 );
xor ( n62779 , n62773 , n62778 );
xor ( n62780 , n62763 , n62779 );
xor ( n62781 , n62743 , n62780 );
xor ( n62782 , n62734 , n62781 );
xor ( n62783 , n62725 , n62782 );
xor ( n62784 , n62716 , n62783 );
xor ( n62785 , n62707 , n62784 );
and ( n62786 , n61712 , n61774 );
and ( n62787 , n61599 , n61669 );
and ( n62788 , n61669 , n61706 );
and ( n62789 , n61599 , n61706 );
or ( n62790 , n62787 , n62788 , n62789 );
and ( n62791 , n61716 , n61773 );
xor ( n62792 , n62790 , n62791 );
and ( n62793 , n61674 , n61678 );
and ( n62794 , n61678 , n61705 );
and ( n62795 , n61674 , n61705 );
or ( n62796 , n62793 , n62794 , n62795 );
and ( n62797 , n61633 , n61649 );
and ( n62798 , n61649 , n61667 );
and ( n62799 , n61633 , n61667 );
or ( n62800 , n62797 , n62798 , n62799 );
and ( n62801 , n61616 , n61620 );
and ( n62802 , n61620 , n61626 );
and ( n62803 , n61616 , n61626 );
or ( n62804 , n62801 , n62802 , n62803 );
and ( n62805 , n61637 , n61642 );
and ( n62806 , n61642 , n61648 );
and ( n62807 , n61637 , n61648 );
or ( n62808 , n62805 , n62806 , n62807 );
xor ( n62809 , n62804 , n62808 );
and ( n62810 , n61622 , n61623 );
and ( n62811 , n61623 , n61625 );
and ( n62812 , n61622 , n61625 );
or ( n62813 , n62810 , n62811 , n62812 );
and ( n62814 , n61638 , n61639 );
and ( n62815 , n61639 , n61641 );
and ( n62816 , n61638 , n61641 );
or ( n62817 , n62814 , n62815 , n62816 );
xor ( n62818 , n62813 , n62817 );
and ( n62819 , n21216 , n8669 );
and ( n62820 , n22186 , n8243 );
xor ( n62821 , n62819 , n62820 );
and ( n62822 , n22892 , n7662 );
xor ( n62823 , n62821 , n62822 );
xor ( n62824 , n62818 , n62823 );
xor ( n62825 , n62809 , n62824 );
xor ( n62826 , n62800 , n62825 );
and ( n62827 , n61656 , n61660 );
and ( n62828 , n61660 , n61666 );
and ( n62829 , n61656 , n61666 );
or ( n62830 , n62827 , n62828 , n62829 );
and ( n62831 , n61644 , n61645 );
and ( n62832 , n61645 , n61647 );
and ( n62833 , n61644 , n61647 );
or ( n62834 , n62831 , n62832 , n62833 );
and ( n62835 , n18144 , n10977 );
and ( n62836 , n19324 , n10239 );
xor ( n62837 , n62835 , n62836 );
and ( n62838 , n20233 , n9348 );
xor ( n62839 , n62837 , n62838 );
xor ( n62840 , n62834 , n62839 );
and ( n62841 , n15758 , n13256 );
and ( n62842 , n16637 , n12531 );
xor ( n62843 , n62841 , n62842 );
and ( n62844 , n17512 , n11718 );
xor ( n62845 , n62843 , n62844 );
xor ( n62846 , n62840 , n62845 );
xor ( n62847 , n62830 , n62846 );
and ( n62848 , n61662 , n61663 );
and ( n62849 , n61663 , n61665 );
and ( n62850 , n61662 , n61665 );
or ( n62851 , n62848 , n62849 , n62850 );
and ( n62852 , n61693 , n61694 );
and ( n62853 , n61694 , n61696 );
and ( n62854 , n61693 , n61696 );
or ( n62855 , n62852 , n62853 , n62854 );
xor ( n62856 , n62851 , n62855 );
and ( n62857 , n13322 , n15691 );
and ( n62858 , n14118 , n14838 );
xor ( n62859 , n62857 , n62858 );
and ( n62860 , n14938 , n14044 );
xor ( n62861 , n62859 , n62860 );
xor ( n62862 , n62856 , n62861 );
xor ( n62863 , n62847 , n62862 );
xor ( n62864 , n62826 , n62863 );
xor ( n62865 , n62796 , n62864 );
and ( n62866 , n61683 , n61687 );
and ( n62867 , n61687 , n61704 );
and ( n62868 , n61683 , n61704 );
or ( n62869 , n62866 , n62867 , n62868 );
and ( n62870 , n61721 , n61736 );
and ( n62871 , n61736 , n61753 );
and ( n62872 , n61721 , n61753 );
or ( n62873 , n62870 , n62871 , n62872 );
xor ( n62874 , n62869 , n62873 );
and ( n62875 , n61692 , n61697 );
and ( n62876 , n61697 , n61703 );
and ( n62877 , n61692 , n61703 );
or ( n62878 , n62875 , n62876 , n62877 );
and ( n62879 , n61725 , n61729 );
and ( n62880 , n61729 , n61735 );
and ( n62881 , n61725 , n61735 );
or ( n62882 , n62879 , n62880 , n62881 );
xor ( n62883 , n62878 , n62882 );
and ( n62884 , n61699 , n61700 );
and ( n62885 , n61700 , n61702 );
and ( n62886 , n61699 , n61702 );
or ( n62887 , n62884 , n62885 , n62886 );
and ( n62888 , n11015 , n18407 );
and ( n62889 , n11769 , n17422 );
xor ( n62890 , n62888 , n62889 );
and ( n62891 , n12320 , n16550 );
xor ( n62892 , n62890 , n62891 );
xor ( n62893 , n62887 , n62892 );
and ( n62894 , n8718 , n20976 );
and ( n62895 , n9400 , n20156 );
xor ( n62896 , n62894 , n62895 );
and ( n62897 , n10291 , n19222 );
xor ( n62898 , n62896 , n62897 );
xor ( n62899 , n62893 , n62898 );
xor ( n62900 , n62883 , n62899 );
xor ( n62901 , n62874 , n62900 );
xor ( n62902 , n62865 , n62901 );
xor ( n62903 , n62792 , n62902 );
xor ( n62904 , n62786 , n62903 );
and ( n62905 , n61717 , n61754 );
and ( n62906 , n61754 , n61772 );
and ( n62907 , n61717 , n61772 );
or ( n62908 , n62905 , n62906 , n62907 );
and ( n62909 , n61759 , n61771 );
and ( n62910 , n61741 , n61746 );
and ( n62911 , n61746 , n61752 );
and ( n62912 , n61741 , n61752 );
or ( n62913 , n62910 , n62911 , n62912 );
and ( n62914 , n61731 , n61732 );
and ( n62915 , n61732 , n61734 );
and ( n62916 , n61731 , n61734 );
or ( n62917 , n62914 , n62915 , n62916 );
and ( n62918 , n61742 , n61743 );
and ( n62919 , n61743 , n61745 );
and ( n62920 , n61742 , n61745 );
or ( n62921 , n62918 , n62919 , n62920 );
xor ( n62922 , n62917 , n62921 );
and ( n62923 , n7385 , n24137 );
and ( n62924 , n7808 , n23075 );
xor ( n62925 , n62923 , n62924 );
and ( n62926 , n8079 , n22065 );
xor ( n62927 , n62925 , n62926 );
xor ( n62928 , n62922 , n62927 );
xor ( n62929 , n62913 , n62928 );
and ( n62930 , n61748 , n61749 );
and ( n62931 , n61749 , n61751 );
and ( n62932 , n61748 , n61751 );
or ( n62933 , n62930 , n62931 , n62932 );
and ( n62934 , n6187 , n27296 );
and ( n62935 , n6569 , n26216 );
xor ( n62936 , n62934 , n62935 );
and ( n62937 , n6816 , n25163 );
xor ( n62938 , n62936 , n62937 );
xor ( n62939 , n62933 , n62938 );
and ( n62940 , n4959 , n30629 );
and ( n62941 , n5459 , n29508 );
xor ( n62942 , n62940 , n62941 );
and ( n62943 , n5819 , n28406 );
xor ( n62944 , n62942 , n62943 );
xor ( n62945 , n62939 , n62944 );
xor ( n62946 , n62929 , n62945 );
xor ( n62947 , n62909 , n62946 );
and ( n62948 , n61763 , n61764 );
and ( n62949 , n61764 , n61770 );
and ( n62950 , n61763 , n61770 );
or ( n62951 , n62948 , n62949 , n62950 );
and ( n62952 , n61766 , n61767 );
and ( n62953 , n61767 , n61769 );
and ( n62954 , n61766 , n61769 );
or ( n62955 , n62952 , n62953 , n62954 );
not ( n62956 , n4132 );
and ( n62957 , n34193 , n4132 );
nor ( n62958 , n62956 , n62957 );
and ( n62959 , n4438 , n32999 );
xor ( n62960 , n62958 , n62959 );
and ( n62961 , n4766 , n31761 );
xor ( n62962 , n62960 , n62961 );
xor ( n62963 , n62955 , n62962 );
xor ( n62964 , n62951 , n62963 );
xor ( n62965 , n62947 , n62964 );
xor ( n62966 , n62908 , n62965 );
xor ( n62967 , n62904 , n62966 );
xor ( n62968 , n62785 , n62967 );
xor ( n62969 , n62703 , n62968 );
xor ( n62970 , n62694 , n62969 );
and ( n62971 , n61493 , n61496 );
and ( n62972 , n61496 , n61778 );
and ( n62973 , n61493 , n61778 );
or ( n62974 , n62971 , n62972 , n62973 );
xor ( n62975 , n62970 , n62974 );
and ( n62976 , n61779 , n61783 );
and ( n62977 , n61784 , n61787 );
or ( n62978 , n62976 , n62977 );
xor ( n62979 , n62975 , n62978 );
buf ( n62980 , n62979 );
buf ( n62981 , n62980 );
not ( n62982 , n62981 );
nor ( n62983 , n62982 , n8739 );
xor ( n62984 , n62686 , n62983 );
and ( n62985 , n61489 , n61792 );
and ( n62986 , n61793 , n61796 );
or ( n62987 , n62985 , n62986 );
xor ( n62988 , n62984 , n62987 );
buf ( n62989 , n62988 );
buf ( n62990 , n62989 );
not ( n62991 , n62990 );
buf ( n62992 , n586 );
not ( n62993 , n62992 );
nor ( n62994 , n62991 , n62993 );
xor ( n62995 , n62312 , n62994 );
xor ( n62996 , n61808 , n62309 );
nor ( n62997 , n61800 , n62993 );
and ( n62998 , n62996 , n62997 );
xor ( n62999 , n62996 , n62997 );
xor ( n63000 , n61812 , n62307 );
nor ( n63001 , n60609 , n62993 );
and ( n63002 , n63000 , n63001 );
xor ( n63003 , n63000 , n63001 );
xor ( n63004 , n61816 , n62305 );
nor ( n63005 , n59421 , n62993 );
and ( n63006 , n63004 , n63005 );
xor ( n63007 , n63004 , n63005 );
xor ( n63008 , n61820 , n62303 );
nor ( n63009 , n58226 , n62993 );
and ( n63010 , n63008 , n63009 );
xor ( n63011 , n63008 , n63009 );
xor ( n63012 , n61824 , n62301 );
nor ( n63013 , n57031 , n62993 );
and ( n63014 , n63012 , n63013 );
xor ( n63015 , n63012 , n63013 );
xor ( n63016 , n61828 , n62299 );
nor ( n63017 , n55835 , n62993 );
and ( n63018 , n63016 , n63017 );
xor ( n63019 , n63016 , n63017 );
xor ( n63020 , n61832 , n62297 );
nor ( n63021 , n54638 , n62993 );
and ( n63022 , n63020 , n63021 );
xor ( n63023 , n63020 , n63021 );
xor ( n63024 , n61836 , n62295 );
nor ( n63025 , n53441 , n62993 );
and ( n63026 , n63024 , n63025 );
xor ( n63027 , n63024 , n63025 );
xor ( n63028 , n61840 , n62293 );
nor ( n63029 , n52247 , n62993 );
and ( n63030 , n63028 , n63029 );
xor ( n63031 , n63028 , n63029 );
xor ( n63032 , n61844 , n62291 );
nor ( n63033 , n51049 , n62993 );
and ( n63034 , n63032 , n63033 );
xor ( n63035 , n63032 , n63033 );
xor ( n63036 , n61848 , n62289 );
nor ( n63037 , n49850 , n62993 );
and ( n63038 , n63036 , n63037 );
xor ( n63039 , n63036 , n63037 );
xor ( n63040 , n61852 , n62287 );
nor ( n63041 , n48650 , n62993 );
and ( n63042 , n63040 , n63041 );
xor ( n63043 , n63040 , n63041 );
xor ( n63044 , n61856 , n62285 );
nor ( n63045 , n47449 , n62993 );
and ( n63046 , n63044 , n63045 );
xor ( n63047 , n63044 , n63045 );
xor ( n63048 , n61860 , n62283 );
nor ( n63049 , n46248 , n62993 );
and ( n63050 , n63048 , n63049 );
xor ( n63051 , n63048 , n63049 );
xor ( n63052 , n61864 , n62281 );
nor ( n63053 , n45047 , n62993 );
and ( n63054 , n63052 , n63053 );
xor ( n63055 , n63052 , n63053 );
xor ( n63056 , n61868 , n62279 );
nor ( n63057 , n43843 , n62993 );
and ( n63058 , n63056 , n63057 );
xor ( n63059 , n63056 , n63057 );
xor ( n63060 , n61872 , n62277 );
nor ( n63061 , n42641 , n62993 );
and ( n63062 , n63060 , n63061 );
xor ( n63063 , n63060 , n63061 );
xor ( n63064 , n61876 , n62275 );
nor ( n63065 , n41437 , n62993 );
and ( n63066 , n63064 , n63065 );
xor ( n63067 , n63064 , n63065 );
xor ( n63068 , n61880 , n62273 );
nor ( n63069 , n40232 , n62993 );
and ( n63070 , n63068 , n63069 );
xor ( n63071 , n63068 , n63069 );
xor ( n63072 , n61884 , n62271 );
nor ( n63073 , n39027 , n62993 );
and ( n63074 , n63072 , n63073 );
xor ( n63075 , n63072 , n63073 );
xor ( n63076 , n61888 , n62269 );
nor ( n63077 , n37825 , n62993 );
and ( n63078 , n63076 , n63077 );
xor ( n63079 , n63076 , n63077 );
xor ( n63080 , n61892 , n62267 );
nor ( n63081 , n36620 , n62993 );
and ( n63082 , n63080 , n63081 );
xor ( n63083 , n63080 , n63081 );
xor ( n63084 , n61896 , n62265 );
nor ( n63085 , n35419 , n62993 );
and ( n63086 , n63084 , n63085 );
xor ( n63087 , n63084 , n63085 );
xor ( n63088 , n61900 , n62263 );
nor ( n63089 , n34224 , n62993 );
and ( n63090 , n63088 , n63089 );
xor ( n63091 , n63088 , n63089 );
xor ( n63092 , n61904 , n62261 );
nor ( n63093 , n33033 , n62993 );
and ( n63094 , n63092 , n63093 );
xor ( n63095 , n63092 , n63093 );
xor ( n63096 , n61908 , n62259 );
nor ( n63097 , n31867 , n62993 );
and ( n63098 , n63096 , n63097 );
xor ( n63099 , n63096 , n63097 );
xor ( n63100 , n61912 , n62257 );
nor ( n63101 , n30725 , n62993 );
and ( n63102 , n63100 , n63101 );
xor ( n63103 , n63100 , n63101 );
xor ( n63104 , n61916 , n62255 );
nor ( n63105 , n29596 , n62993 );
and ( n63106 , n63104 , n63105 );
xor ( n63107 , n63104 , n63105 );
xor ( n63108 , n61920 , n62253 );
nor ( n63109 , n28487 , n62993 );
and ( n63110 , n63108 , n63109 );
xor ( n63111 , n63108 , n63109 );
xor ( n63112 , n61924 , n62251 );
nor ( n63113 , n27397 , n62993 );
and ( n63114 , n63112 , n63113 );
xor ( n63115 , n63112 , n63113 );
xor ( n63116 , n61928 , n62249 );
nor ( n63117 , n26326 , n62993 );
and ( n63118 , n63116 , n63117 );
xor ( n63119 , n63116 , n63117 );
xor ( n63120 , n61932 , n62247 );
nor ( n63121 , n25272 , n62993 );
and ( n63122 , n63120 , n63121 );
xor ( n63123 , n63120 , n63121 );
xor ( n63124 , n61936 , n62245 );
nor ( n63125 , n24242 , n62993 );
and ( n63126 , n63124 , n63125 );
xor ( n63127 , n63124 , n63125 );
xor ( n63128 , n61940 , n62243 );
nor ( n63129 , n23225 , n62993 );
and ( n63130 , n63128 , n63129 );
xor ( n63131 , n63128 , n63129 );
xor ( n63132 , n61944 , n62241 );
nor ( n63133 , n22231 , n62993 );
and ( n63134 , n63132 , n63133 );
xor ( n63135 , n63132 , n63133 );
xor ( n63136 , n61948 , n62239 );
nor ( n63137 , n21258 , n62993 );
and ( n63138 , n63136 , n63137 );
xor ( n63139 , n63136 , n63137 );
xor ( n63140 , n61952 , n62237 );
nor ( n63141 , n20303 , n62993 );
and ( n63142 , n63140 , n63141 );
xor ( n63143 , n63140 , n63141 );
xor ( n63144 , n61956 , n62235 );
nor ( n63145 , n19365 , n62993 );
and ( n63146 , n63144 , n63145 );
xor ( n63147 , n63144 , n63145 );
xor ( n63148 , n61960 , n62233 );
nor ( n63149 , n18448 , n62993 );
and ( n63150 , n63148 , n63149 );
xor ( n63151 , n63148 , n63149 );
xor ( n63152 , n61964 , n62231 );
nor ( n63153 , n17548 , n62993 );
and ( n63154 , n63152 , n63153 );
xor ( n63155 , n63152 , n63153 );
xor ( n63156 , n61968 , n62229 );
nor ( n63157 , n16669 , n62993 );
and ( n63158 , n63156 , n63157 );
xor ( n63159 , n63156 , n63157 );
xor ( n63160 , n61972 , n62227 );
nor ( n63161 , n15809 , n62993 );
and ( n63162 , n63160 , n63161 );
xor ( n63163 , n63160 , n63161 );
xor ( n63164 , n61976 , n62225 );
nor ( n63165 , n14968 , n62993 );
and ( n63166 , n63164 , n63165 );
xor ( n63167 , n63164 , n63165 );
xor ( n63168 , n61980 , n62223 );
nor ( n63169 , n14147 , n62993 );
and ( n63170 , n63168 , n63169 );
xor ( n63171 , n63168 , n63169 );
xor ( n63172 , n61984 , n62221 );
nor ( n63173 , n13349 , n62993 );
and ( n63174 , n63172 , n63173 );
xor ( n63175 , n63172 , n63173 );
xor ( n63176 , n61988 , n62219 );
nor ( n63177 , n12564 , n62993 );
and ( n63178 , n63176 , n63177 );
xor ( n63179 , n63176 , n63177 );
xor ( n63180 , n61992 , n62217 );
nor ( n63181 , n11799 , n62993 );
and ( n63182 , n63180 , n63181 );
xor ( n63183 , n63180 , n63181 );
xor ( n63184 , n61996 , n62215 );
nor ( n63185 , n11050 , n62993 );
and ( n63186 , n63184 , n63185 );
xor ( n63187 , n63184 , n63185 );
xor ( n63188 , n62000 , n62213 );
nor ( n63189 , n10321 , n62993 );
and ( n63190 , n63188 , n63189 );
xor ( n63191 , n63188 , n63189 );
xor ( n63192 , n62004 , n62211 );
nor ( n63193 , n9429 , n62993 );
and ( n63194 , n63192 , n63193 );
xor ( n63195 , n63192 , n63193 );
xor ( n63196 , n62008 , n62209 );
nor ( n63197 , n8949 , n62993 );
and ( n63198 , n63196 , n63197 );
xor ( n63199 , n63196 , n63197 );
xor ( n63200 , n62012 , n62207 );
nor ( n63201 , n9437 , n62993 );
and ( n63202 , n63200 , n63201 );
xor ( n63203 , n63200 , n63201 );
xor ( n63204 , n62016 , n62205 );
nor ( n63205 , n9446 , n62993 );
and ( n63206 , n63204 , n63205 );
xor ( n63207 , n63204 , n63205 );
xor ( n63208 , n62020 , n62203 );
nor ( n63209 , n9455 , n62993 );
and ( n63210 , n63208 , n63209 );
xor ( n63211 , n63208 , n63209 );
xor ( n63212 , n62024 , n62201 );
nor ( n63213 , n9464 , n62993 );
and ( n63214 , n63212 , n63213 );
xor ( n63215 , n63212 , n63213 );
xor ( n63216 , n62028 , n62199 );
nor ( n63217 , n9473 , n62993 );
and ( n63218 , n63216 , n63217 );
xor ( n63219 , n63216 , n63217 );
xor ( n63220 , n62032 , n62197 );
nor ( n63221 , n9482 , n62993 );
and ( n63222 , n63220 , n63221 );
xor ( n63223 , n63220 , n63221 );
xor ( n63224 , n62036 , n62195 );
nor ( n63225 , n9491 , n62993 );
and ( n63226 , n63224 , n63225 );
xor ( n63227 , n63224 , n63225 );
xor ( n63228 , n62040 , n62193 );
nor ( n63229 , n9500 , n62993 );
and ( n63230 , n63228 , n63229 );
xor ( n63231 , n63228 , n63229 );
xor ( n63232 , n62044 , n62191 );
nor ( n63233 , n9509 , n62993 );
and ( n63234 , n63232 , n63233 );
xor ( n63235 , n63232 , n63233 );
xor ( n63236 , n62048 , n62189 );
nor ( n63237 , n9518 , n62993 );
and ( n63238 , n63236 , n63237 );
xor ( n63239 , n63236 , n63237 );
xor ( n63240 , n62052 , n62187 );
nor ( n63241 , n9527 , n62993 );
and ( n63242 , n63240 , n63241 );
xor ( n63243 , n63240 , n63241 );
xor ( n63244 , n62056 , n62185 );
nor ( n63245 , n9536 , n62993 );
and ( n63246 , n63244 , n63245 );
xor ( n63247 , n63244 , n63245 );
xor ( n63248 , n62060 , n62183 );
nor ( n63249 , n9545 , n62993 );
and ( n63250 , n63248 , n63249 );
xor ( n63251 , n63248 , n63249 );
xor ( n63252 , n62064 , n62181 );
nor ( n63253 , n9554 , n62993 );
and ( n63254 , n63252 , n63253 );
xor ( n63255 , n63252 , n63253 );
xor ( n63256 , n62068 , n62179 );
nor ( n63257 , n9563 , n62993 );
and ( n63258 , n63256 , n63257 );
xor ( n63259 , n63256 , n63257 );
xor ( n63260 , n62072 , n62177 );
nor ( n63261 , n9572 , n62993 );
and ( n63262 , n63260 , n63261 );
xor ( n63263 , n63260 , n63261 );
xor ( n63264 , n62076 , n62175 );
nor ( n63265 , n9581 , n62993 );
and ( n63266 , n63264 , n63265 );
xor ( n63267 , n63264 , n63265 );
xor ( n63268 , n62080 , n62173 );
nor ( n63269 , n9590 , n62993 );
and ( n63270 , n63268 , n63269 );
xor ( n63271 , n63268 , n63269 );
xor ( n63272 , n62084 , n62171 );
nor ( n63273 , n9599 , n62993 );
and ( n63274 , n63272 , n63273 );
xor ( n63275 , n63272 , n63273 );
xor ( n63276 , n62088 , n62169 );
nor ( n63277 , n9608 , n62993 );
and ( n63278 , n63276 , n63277 );
xor ( n63279 , n63276 , n63277 );
xor ( n63280 , n62092 , n62167 );
nor ( n63281 , n9617 , n62993 );
and ( n63282 , n63280 , n63281 );
xor ( n63283 , n63280 , n63281 );
xor ( n63284 , n62096 , n62165 );
nor ( n63285 , n9626 , n62993 );
and ( n63286 , n63284 , n63285 );
xor ( n63287 , n63284 , n63285 );
xor ( n63288 , n62100 , n62163 );
nor ( n63289 , n9635 , n62993 );
and ( n63290 , n63288 , n63289 );
xor ( n63291 , n63288 , n63289 );
xor ( n63292 , n62104 , n62161 );
nor ( n63293 , n9644 , n62993 );
and ( n63294 , n63292 , n63293 );
xor ( n63295 , n63292 , n63293 );
xor ( n63296 , n62108 , n62159 );
nor ( n63297 , n9653 , n62993 );
and ( n63298 , n63296 , n63297 );
xor ( n63299 , n63296 , n63297 );
xor ( n63300 , n62112 , n62157 );
nor ( n63301 , n9662 , n62993 );
and ( n63302 , n63300 , n63301 );
xor ( n63303 , n63300 , n63301 );
xor ( n63304 , n62116 , n62155 );
nor ( n63305 , n9671 , n62993 );
and ( n63306 , n63304 , n63305 );
xor ( n63307 , n63304 , n63305 );
xor ( n63308 , n62120 , n62153 );
nor ( n63309 , n9680 , n62993 );
and ( n63310 , n63308 , n63309 );
xor ( n63311 , n63308 , n63309 );
xor ( n63312 , n62124 , n62151 );
nor ( n63313 , n9689 , n62993 );
and ( n63314 , n63312 , n63313 );
xor ( n63315 , n63312 , n63313 );
xor ( n63316 , n62128 , n62149 );
nor ( n63317 , n9698 , n62993 );
and ( n63318 , n63316 , n63317 );
xor ( n63319 , n63316 , n63317 );
xor ( n63320 , n62132 , n62147 );
nor ( n63321 , n9707 , n62993 );
and ( n63322 , n63320 , n63321 );
xor ( n63323 , n63320 , n63321 );
xor ( n63324 , n62136 , n62145 );
nor ( n63325 , n9716 , n62993 );
and ( n63326 , n63324 , n63325 );
xor ( n63327 , n63324 , n63325 );
xor ( n63328 , n62140 , n62143 );
nor ( n63329 , n9725 , n62993 );
and ( n63330 , n63328 , n63329 );
xor ( n63331 , n63328 , n63329 );
xor ( n63332 , n62141 , n62142 );
nor ( n63333 , n9734 , n62993 );
and ( n63334 , n63332 , n63333 );
xor ( n63335 , n63332 , n63333 );
nor ( n63336 , n9752 , n61802 );
nor ( n63337 , n9743 , n62993 );
and ( n63338 , n63336 , n63337 );
and ( n63339 , n63335 , n63338 );
or ( n63340 , n63334 , n63339 );
and ( n63341 , n63331 , n63340 );
or ( n63342 , n63330 , n63341 );
and ( n63343 , n63327 , n63342 );
or ( n63344 , n63326 , n63343 );
and ( n63345 , n63323 , n63344 );
or ( n63346 , n63322 , n63345 );
and ( n63347 , n63319 , n63346 );
or ( n63348 , n63318 , n63347 );
and ( n63349 , n63315 , n63348 );
or ( n63350 , n63314 , n63349 );
and ( n63351 , n63311 , n63350 );
or ( n63352 , n63310 , n63351 );
and ( n63353 , n63307 , n63352 );
or ( n63354 , n63306 , n63353 );
and ( n63355 , n63303 , n63354 );
or ( n63356 , n63302 , n63355 );
and ( n63357 , n63299 , n63356 );
or ( n63358 , n63298 , n63357 );
and ( n63359 , n63295 , n63358 );
or ( n63360 , n63294 , n63359 );
and ( n63361 , n63291 , n63360 );
or ( n63362 , n63290 , n63361 );
and ( n63363 , n63287 , n63362 );
or ( n63364 , n63286 , n63363 );
and ( n63365 , n63283 , n63364 );
or ( n63366 , n63282 , n63365 );
and ( n63367 , n63279 , n63366 );
or ( n63368 , n63278 , n63367 );
and ( n63369 , n63275 , n63368 );
or ( n63370 , n63274 , n63369 );
and ( n63371 , n63271 , n63370 );
or ( n63372 , n63270 , n63371 );
and ( n63373 , n63267 , n63372 );
or ( n63374 , n63266 , n63373 );
and ( n63375 , n63263 , n63374 );
or ( n63376 , n63262 , n63375 );
and ( n63377 , n63259 , n63376 );
or ( n63378 , n63258 , n63377 );
and ( n63379 , n63255 , n63378 );
or ( n63380 , n63254 , n63379 );
and ( n63381 , n63251 , n63380 );
or ( n63382 , n63250 , n63381 );
and ( n63383 , n63247 , n63382 );
or ( n63384 , n63246 , n63383 );
and ( n63385 , n63243 , n63384 );
or ( n63386 , n63242 , n63385 );
and ( n63387 , n63239 , n63386 );
or ( n63388 , n63238 , n63387 );
and ( n63389 , n63235 , n63388 );
or ( n63390 , n63234 , n63389 );
and ( n63391 , n63231 , n63390 );
or ( n63392 , n63230 , n63391 );
and ( n63393 , n63227 , n63392 );
or ( n63394 , n63226 , n63393 );
and ( n63395 , n63223 , n63394 );
or ( n63396 , n63222 , n63395 );
and ( n63397 , n63219 , n63396 );
or ( n63398 , n63218 , n63397 );
and ( n63399 , n63215 , n63398 );
or ( n63400 , n63214 , n63399 );
and ( n63401 , n63211 , n63400 );
or ( n63402 , n63210 , n63401 );
and ( n63403 , n63207 , n63402 );
or ( n63404 , n63206 , n63403 );
and ( n63405 , n63203 , n63404 );
or ( n63406 , n63202 , n63405 );
and ( n63407 , n63199 , n63406 );
or ( n63408 , n63198 , n63407 );
and ( n63409 , n63195 , n63408 );
or ( n63410 , n63194 , n63409 );
and ( n63411 , n63191 , n63410 );
or ( n63412 , n63190 , n63411 );
and ( n63413 , n63187 , n63412 );
or ( n63414 , n63186 , n63413 );
and ( n63415 , n63183 , n63414 );
or ( n63416 , n63182 , n63415 );
and ( n63417 , n63179 , n63416 );
or ( n63418 , n63178 , n63417 );
and ( n63419 , n63175 , n63418 );
or ( n63420 , n63174 , n63419 );
and ( n63421 , n63171 , n63420 );
or ( n63422 , n63170 , n63421 );
and ( n63423 , n63167 , n63422 );
or ( n63424 , n63166 , n63423 );
and ( n63425 , n63163 , n63424 );
or ( n63426 , n63162 , n63425 );
and ( n63427 , n63159 , n63426 );
or ( n63428 , n63158 , n63427 );
and ( n63429 , n63155 , n63428 );
or ( n63430 , n63154 , n63429 );
and ( n63431 , n63151 , n63430 );
or ( n63432 , n63150 , n63431 );
and ( n63433 , n63147 , n63432 );
or ( n63434 , n63146 , n63433 );
and ( n63435 , n63143 , n63434 );
or ( n63436 , n63142 , n63435 );
and ( n63437 , n63139 , n63436 );
or ( n63438 , n63138 , n63437 );
and ( n63439 , n63135 , n63438 );
or ( n63440 , n63134 , n63439 );
and ( n63441 , n63131 , n63440 );
or ( n63442 , n63130 , n63441 );
and ( n63443 , n63127 , n63442 );
or ( n63444 , n63126 , n63443 );
and ( n63445 , n63123 , n63444 );
or ( n63446 , n63122 , n63445 );
and ( n63447 , n63119 , n63446 );
or ( n63448 , n63118 , n63447 );
and ( n63449 , n63115 , n63448 );
or ( n63450 , n63114 , n63449 );
and ( n63451 , n63111 , n63450 );
or ( n63452 , n63110 , n63451 );
and ( n63453 , n63107 , n63452 );
or ( n63454 , n63106 , n63453 );
and ( n63455 , n63103 , n63454 );
or ( n63456 , n63102 , n63455 );
and ( n63457 , n63099 , n63456 );
or ( n63458 , n63098 , n63457 );
and ( n63459 , n63095 , n63458 );
or ( n63460 , n63094 , n63459 );
and ( n63461 , n63091 , n63460 );
or ( n63462 , n63090 , n63461 );
and ( n63463 , n63087 , n63462 );
or ( n63464 , n63086 , n63463 );
and ( n63465 , n63083 , n63464 );
or ( n63466 , n63082 , n63465 );
and ( n63467 , n63079 , n63466 );
or ( n63468 , n63078 , n63467 );
and ( n63469 , n63075 , n63468 );
or ( n63470 , n63074 , n63469 );
and ( n63471 , n63071 , n63470 );
or ( n63472 , n63070 , n63471 );
and ( n63473 , n63067 , n63472 );
or ( n63474 , n63066 , n63473 );
and ( n63475 , n63063 , n63474 );
or ( n63476 , n63062 , n63475 );
and ( n63477 , n63059 , n63476 );
or ( n63478 , n63058 , n63477 );
and ( n63479 , n63055 , n63478 );
or ( n63480 , n63054 , n63479 );
and ( n63481 , n63051 , n63480 );
or ( n63482 , n63050 , n63481 );
and ( n63483 , n63047 , n63482 );
or ( n63484 , n63046 , n63483 );
and ( n63485 , n63043 , n63484 );
or ( n63486 , n63042 , n63485 );
and ( n63487 , n63039 , n63486 );
or ( n63488 , n63038 , n63487 );
and ( n63489 , n63035 , n63488 );
or ( n63490 , n63034 , n63489 );
and ( n63491 , n63031 , n63490 );
or ( n63492 , n63030 , n63491 );
and ( n63493 , n63027 , n63492 );
or ( n63494 , n63026 , n63493 );
and ( n63495 , n63023 , n63494 );
or ( n63496 , n63022 , n63495 );
and ( n63497 , n63019 , n63496 );
or ( n63498 , n63018 , n63497 );
and ( n63499 , n63015 , n63498 );
or ( n63500 , n63014 , n63499 );
and ( n63501 , n63011 , n63500 );
or ( n63502 , n63010 , n63501 );
and ( n63503 , n63007 , n63502 );
or ( n63504 , n63006 , n63503 );
and ( n63505 , n63003 , n63504 );
or ( n63506 , n63002 , n63505 );
and ( n63507 , n62999 , n63506 );
or ( n63508 , n62998 , n63507 );
xor ( n63509 , n62995 , n63508 );
and ( n63510 , n33403 , n4457 );
nor ( n63511 , n4458 , n63510 );
nor ( n63512 , n4786 , n32231 );
xor ( n63513 , n63511 , n63512 );
and ( n63514 , n62314 , n62315 );
and ( n63515 , n62316 , n62319 );
or ( n63516 , n63514 , n63515 );
xor ( n63517 , n63513 , n63516 );
nor ( n63518 , n5126 , n31083 );
xor ( n63519 , n63517 , n63518 );
and ( n63520 , n62320 , n62321 );
and ( n63521 , n62322 , n62325 );
or ( n63522 , n63520 , n63521 );
xor ( n63523 , n63519 , n63522 );
nor ( n63524 , n5477 , n29948 );
xor ( n63525 , n63523 , n63524 );
and ( n63526 , n62326 , n62327 );
and ( n63527 , n62328 , n62331 );
or ( n63528 , n63526 , n63527 );
xor ( n63529 , n63525 , n63528 );
nor ( n63530 , n5838 , n28833 );
xor ( n63531 , n63529 , n63530 );
and ( n63532 , n62332 , n62333 );
and ( n63533 , n62334 , n62337 );
or ( n63534 , n63532 , n63533 );
xor ( n63535 , n63531 , n63534 );
nor ( n63536 , n6212 , n27737 );
xor ( n63537 , n63535 , n63536 );
and ( n63538 , n62338 , n62339 );
and ( n63539 , n62340 , n62343 );
or ( n63540 , n63538 , n63539 );
xor ( n63541 , n63537 , n63540 );
nor ( n63542 , n6596 , n26660 );
xor ( n63543 , n63541 , n63542 );
and ( n63544 , n62344 , n62345 );
and ( n63545 , n62346 , n62349 );
or ( n63546 , n63544 , n63545 );
xor ( n63547 , n63543 , n63546 );
nor ( n63548 , n6997 , n25600 );
xor ( n63549 , n63547 , n63548 );
and ( n63550 , n62350 , n62351 );
and ( n63551 , n62352 , n62355 );
or ( n63552 , n63550 , n63551 );
xor ( n63553 , n63549 , n63552 );
nor ( n63554 , n7413 , n24564 );
xor ( n63555 , n63553 , n63554 );
and ( n63556 , n62356 , n62357 );
and ( n63557 , n62358 , n62361 );
or ( n63558 , n63556 , n63557 );
xor ( n63559 , n63555 , n63558 );
nor ( n63560 , n7841 , n23541 );
xor ( n63561 , n63559 , n63560 );
and ( n63562 , n62362 , n62363 );
and ( n63563 , n62364 , n62367 );
or ( n63564 , n63562 , n63563 );
xor ( n63565 , n63561 , n63564 );
nor ( n63566 , n8281 , n22541 );
xor ( n63567 , n63565 , n63566 );
and ( n63568 , n62368 , n62369 );
and ( n63569 , n62370 , n62373 );
or ( n63570 , n63568 , n63569 );
xor ( n63571 , n63567 , n63570 );
nor ( n63572 , n8737 , n21562 );
xor ( n63573 , n63571 , n63572 );
and ( n63574 , n62374 , n62375 );
and ( n63575 , n62376 , n62379 );
or ( n63576 , n63574 , n63575 );
xor ( n63577 , n63573 , n63576 );
nor ( n63578 , n9420 , n20601 );
xor ( n63579 , n63577 , n63578 );
and ( n63580 , n62380 , n62381 );
and ( n63581 , n62382 , n62385 );
or ( n63582 , n63580 , n63581 );
xor ( n63583 , n63579 , n63582 );
nor ( n63584 , n10312 , n19657 );
xor ( n63585 , n63583 , n63584 );
and ( n63586 , n62386 , n62387 );
and ( n63587 , n62388 , n62391 );
or ( n63588 , n63586 , n63587 );
xor ( n63589 , n63585 , n63588 );
nor ( n63590 , n11041 , n18734 );
xor ( n63591 , n63589 , n63590 );
and ( n63592 , n62392 , n62393 );
and ( n63593 , n62394 , n62397 );
or ( n63594 , n63592 , n63593 );
xor ( n63595 , n63591 , n63594 );
nor ( n63596 , n11790 , n17828 );
xor ( n63597 , n63595 , n63596 );
and ( n63598 , n62398 , n62399 );
and ( n63599 , n62400 , n62403 );
or ( n63600 , n63598 , n63599 );
xor ( n63601 , n63597 , n63600 );
nor ( n63602 , n12555 , n16943 );
xor ( n63603 , n63601 , n63602 );
and ( n63604 , n62404 , n62405 );
and ( n63605 , n62406 , n62409 );
or ( n63606 , n63604 , n63605 );
xor ( n63607 , n63603 , n63606 );
nor ( n63608 , n13340 , n16077 );
xor ( n63609 , n63607 , n63608 );
and ( n63610 , n62410 , n62411 );
and ( n63611 , n62412 , n62415 );
or ( n63612 , n63610 , n63611 );
xor ( n63613 , n63609 , n63612 );
nor ( n63614 , n14138 , n15230 );
xor ( n63615 , n63613 , n63614 );
and ( n63616 , n62416 , n62417 );
and ( n63617 , n62418 , n62421 );
or ( n63618 , n63616 , n63617 );
xor ( n63619 , n63615 , n63618 );
nor ( n63620 , n14959 , n14403 );
xor ( n63621 , n63619 , n63620 );
and ( n63622 , n62422 , n62423 );
and ( n63623 , n62424 , n62427 );
or ( n63624 , n63622 , n63623 );
xor ( n63625 , n63621 , n63624 );
nor ( n63626 , n15800 , n13599 );
xor ( n63627 , n63625 , n63626 );
and ( n63628 , n62428 , n62429 );
and ( n63629 , n62430 , n62433 );
or ( n63630 , n63628 , n63629 );
xor ( n63631 , n63627 , n63630 );
nor ( n63632 , n16660 , n12808 );
xor ( n63633 , n63631 , n63632 );
and ( n63634 , n62434 , n62435 );
and ( n63635 , n62436 , n62439 );
or ( n63636 , n63634 , n63635 );
xor ( n63637 , n63633 , n63636 );
nor ( n63638 , n17539 , n12037 );
xor ( n63639 , n63637 , n63638 );
and ( n63640 , n62440 , n62441 );
and ( n63641 , n62442 , n62445 );
or ( n63642 , n63640 , n63641 );
xor ( n63643 , n63639 , n63642 );
nor ( n63644 , n18439 , n11282 );
xor ( n63645 , n63643 , n63644 );
and ( n63646 , n62446 , n62447 );
and ( n63647 , n62448 , n62451 );
or ( n63648 , n63646 , n63647 );
xor ( n63649 , n63645 , n63648 );
nor ( n63650 , n19356 , n10547 );
xor ( n63651 , n63649 , n63650 );
and ( n63652 , n62452 , n62453 );
and ( n63653 , n62454 , n62457 );
or ( n63654 , n63652 , n63653 );
xor ( n63655 , n63651 , n63654 );
nor ( n63656 , n20294 , n9829 );
xor ( n63657 , n63655 , n63656 );
and ( n63658 , n62458 , n62459 );
and ( n63659 , n62460 , n62463 );
or ( n63660 , n63658 , n63659 );
xor ( n63661 , n63657 , n63660 );
nor ( n63662 , n21249 , n8955 );
xor ( n63663 , n63661 , n63662 );
and ( n63664 , n62464 , n62465 );
and ( n63665 , n62466 , n62469 );
or ( n63666 , n63664 , n63665 );
xor ( n63667 , n63663 , n63666 );
nor ( n63668 , n22222 , n603 );
xor ( n63669 , n63667 , n63668 );
and ( n63670 , n62470 , n62471 );
and ( n63671 , n62472 , n62475 );
or ( n63672 , n63670 , n63671 );
xor ( n63673 , n63669 , n63672 );
nor ( n63674 , n23216 , n652 );
xor ( n63675 , n63673 , n63674 );
and ( n63676 , n62476 , n62477 );
and ( n63677 , n62478 , n62481 );
or ( n63678 , n63676 , n63677 );
xor ( n63679 , n63675 , n63678 );
nor ( n63680 , n24233 , n624 );
xor ( n63681 , n63679 , n63680 );
and ( n63682 , n62482 , n62483 );
and ( n63683 , n62484 , n62487 );
or ( n63684 , n63682 , n63683 );
xor ( n63685 , n63681 , n63684 );
nor ( n63686 , n25263 , n648 );
xor ( n63687 , n63685 , n63686 );
and ( n63688 , n62488 , n62489 );
and ( n63689 , n62490 , n62493 );
or ( n63690 , n63688 , n63689 );
xor ( n63691 , n63687 , n63690 );
nor ( n63692 , n26317 , n686 );
xor ( n63693 , n63691 , n63692 );
and ( n63694 , n62494 , n62495 );
and ( n63695 , n62496 , n62499 );
or ( n63696 , n63694 , n63695 );
xor ( n63697 , n63693 , n63696 );
nor ( n63698 , n27388 , n735 );
xor ( n63699 , n63697 , n63698 );
and ( n63700 , n62500 , n62501 );
and ( n63701 , n62502 , n62505 );
or ( n63702 , n63700 , n63701 );
xor ( n63703 , n63699 , n63702 );
nor ( n63704 , n28478 , n798 );
xor ( n63705 , n63703 , n63704 );
and ( n63706 , n62506 , n62507 );
and ( n63707 , n62508 , n62511 );
or ( n63708 , n63706 , n63707 );
xor ( n63709 , n63705 , n63708 );
nor ( n63710 , n29587 , n870 );
xor ( n63711 , n63709 , n63710 );
and ( n63712 , n62512 , n62513 );
and ( n63713 , n62514 , n62517 );
or ( n63714 , n63712 , n63713 );
xor ( n63715 , n63711 , n63714 );
nor ( n63716 , n30716 , n960 );
xor ( n63717 , n63715 , n63716 );
and ( n63718 , n62518 , n62519 );
and ( n63719 , n62520 , n62523 );
or ( n63720 , n63718 , n63719 );
xor ( n63721 , n63717 , n63720 );
nor ( n63722 , n31858 , n1064 );
xor ( n63723 , n63721 , n63722 );
and ( n63724 , n62524 , n62525 );
and ( n63725 , n62526 , n62529 );
or ( n63726 , n63724 , n63725 );
xor ( n63727 , n63723 , n63726 );
nor ( n63728 , n33024 , n1178 );
xor ( n63729 , n63727 , n63728 );
and ( n63730 , n62530 , n62531 );
and ( n63731 , n62532 , n62535 );
or ( n63732 , n63730 , n63731 );
xor ( n63733 , n63729 , n63732 );
nor ( n63734 , n34215 , n1305 );
xor ( n63735 , n63733 , n63734 );
and ( n63736 , n62536 , n62537 );
and ( n63737 , n62538 , n62541 );
or ( n63738 , n63736 , n63737 );
xor ( n63739 , n63735 , n63738 );
nor ( n63740 , n35410 , n1447 );
xor ( n63741 , n63739 , n63740 );
and ( n63742 , n62542 , n62543 );
and ( n63743 , n62544 , n62547 );
or ( n63744 , n63742 , n63743 );
xor ( n63745 , n63741 , n63744 );
nor ( n63746 , n36611 , n1600 );
xor ( n63747 , n63745 , n63746 );
and ( n63748 , n62548 , n62549 );
and ( n63749 , n62550 , n62553 );
or ( n63750 , n63748 , n63749 );
xor ( n63751 , n63747 , n63750 );
nor ( n63752 , n37816 , n1768 );
xor ( n63753 , n63751 , n63752 );
and ( n63754 , n62554 , n62555 );
and ( n63755 , n62556 , n62559 );
or ( n63756 , n63754 , n63755 );
xor ( n63757 , n63753 , n63756 );
nor ( n63758 , n39018 , n1947 );
xor ( n63759 , n63757 , n63758 );
and ( n63760 , n62560 , n62561 );
and ( n63761 , n62562 , n62565 );
or ( n63762 , n63760 , n63761 );
xor ( n63763 , n63759 , n63762 );
nor ( n63764 , n40223 , n2139 );
xor ( n63765 , n63763 , n63764 );
and ( n63766 , n62566 , n62567 );
and ( n63767 , n62568 , n62571 );
or ( n63768 , n63766 , n63767 );
xor ( n63769 , n63765 , n63768 );
nor ( n63770 , n41428 , n2345 );
xor ( n63771 , n63769 , n63770 );
and ( n63772 , n62572 , n62573 );
and ( n63773 , n62574 , n62577 );
or ( n63774 , n63772 , n63773 );
xor ( n63775 , n63771 , n63774 );
nor ( n63776 , n42632 , n2568 );
xor ( n63777 , n63775 , n63776 );
and ( n63778 , n62578 , n62579 );
and ( n63779 , n62580 , n62583 );
or ( n63780 , n63778 , n63779 );
xor ( n63781 , n63777 , n63780 );
nor ( n63782 , n43834 , n2799 );
xor ( n63783 , n63781 , n63782 );
and ( n63784 , n62584 , n62585 );
and ( n63785 , n62586 , n62589 );
or ( n63786 , n63784 , n63785 );
xor ( n63787 , n63783 , n63786 );
nor ( n63788 , n45038 , n3045 );
xor ( n63789 , n63787 , n63788 );
and ( n63790 , n62590 , n62591 );
and ( n63791 , n62592 , n62595 );
or ( n63792 , n63790 , n63791 );
xor ( n63793 , n63789 , n63792 );
nor ( n63794 , n46239 , n3302 );
xor ( n63795 , n63793 , n63794 );
and ( n63796 , n62596 , n62597 );
and ( n63797 , n62598 , n62601 );
or ( n63798 , n63796 , n63797 );
xor ( n63799 , n63795 , n63798 );
nor ( n63800 , n47440 , n3572 );
xor ( n63801 , n63799 , n63800 );
and ( n63802 , n62602 , n62603 );
and ( n63803 , n62604 , n62607 );
or ( n63804 , n63802 , n63803 );
xor ( n63805 , n63801 , n63804 );
nor ( n63806 , n48641 , n3855 );
xor ( n63807 , n63805 , n63806 );
and ( n63808 , n62608 , n62609 );
and ( n63809 , n62610 , n62613 );
or ( n63810 , n63808 , n63809 );
xor ( n63811 , n63807 , n63810 );
nor ( n63812 , n49841 , n4153 );
xor ( n63813 , n63811 , n63812 );
and ( n63814 , n62614 , n62615 );
and ( n63815 , n62616 , n62619 );
or ( n63816 , n63814 , n63815 );
xor ( n63817 , n63813 , n63816 );
nor ( n63818 , n51040 , n4460 );
xor ( n63819 , n63817 , n63818 );
and ( n63820 , n62620 , n62621 );
and ( n63821 , n62622 , n62625 );
or ( n63822 , n63820 , n63821 );
xor ( n63823 , n63819 , n63822 );
nor ( n63824 , n52238 , n4788 );
xor ( n63825 , n63823 , n63824 );
and ( n63826 , n62626 , n62627 );
and ( n63827 , n62628 , n62631 );
or ( n63828 , n63826 , n63827 );
xor ( n63829 , n63825 , n63828 );
nor ( n63830 , n53432 , n5128 );
xor ( n63831 , n63829 , n63830 );
and ( n63832 , n62632 , n62633 );
and ( n63833 , n62634 , n62637 );
or ( n63834 , n63832 , n63833 );
xor ( n63835 , n63831 , n63834 );
nor ( n63836 , n54629 , n5479 );
xor ( n63837 , n63835 , n63836 );
and ( n63838 , n62638 , n62639 );
and ( n63839 , n62640 , n62643 );
or ( n63840 , n63838 , n63839 );
xor ( n63841 , n63837 , n63840 );
nor ( n63842 , n55826 , n5840 );
xor ( n63843 , n63841 , n63842 );
and ( n63844 , n62644 , n62645 );
and ( n63845 , n62646 , n62649 );
or ( n63846 , n63844 , n63845 );
xor ( n63847 , n63843 , n63846 );
nor ( n63848 , n57022 , n6214 );
xor ( n63849 , n63847 , n63848 );
and ( n63850 , n62650 , n62651 );
and ( n63851 , n62652 , n62655 );
or ( n63852 , n63850 , n63851 );
xor ( n63853 , n63849 , n63852 );
nor ( n63854 , n58217 , n6598 );
xor ( n63855 , n63853 , n63854 );
and ( n63856 , n62656 , n62657 );
and ( n63857 , n62658 , n62661 );
or ( n63858 , n63856 , n63857 );
xor ( n63859 , n63855 , n63858 );
nor ( n63860 , n59412 , n6999 );
xor ( n63861 , n63859 , n63860 );
and ( n63862 , n62662 , n62663 );
and ( n63863 , n62664 , n62667 );
or ( n63864 , n63862 , n63863 );
xor ( n63865 , n63861 , n63864 );
nor ( n63866 , n60600 , n7415 );
xor ( n63867 , n63865 , n63866 );
and ( n63868 , n62668 , n62669 );
and ( n63869 , n62670 , n62673 );
or ( n63870 , n63868 , n63869 );
xor ( n63871 , n63867 , n63870 );
nor ( n63872 , n61791 , n7843 );
xor ( n63873 , n63871 , n63872 );
and ( n63874 , n62674 , n62675 );
and ( n63875 , n62676 , n62679 );
or ( n63876 , n63874 , n63875 );
xor ( n63877 , n63873 , n63876 );
nor ( n63878 , n62982 , n8283 );
xor ( n63879 , n63877 , n63878 );
and ( n63880 , n62680 , n62681 );
and ( n63881 , n62682 , n62685 );
or ( n63882 , n63880 , n63881 );
xor ( n63883 , n63879 , n63882 );
and ( n63884 , n62698 , n62702 );
and ( n63885 , n62702 , n62968 );
and ( n63886 , n62698 , n62968 );
or ( n63887 , n63884 , n63885 , n63886 );
and ( n63888 , n33774 , n4403 );
not ( n63889 , n4403 );
nor ( n63890 , n63888 , n63889 );
xor ( n63891 , n63887 , n63890 );
and ( n63892 , n62711 , n62715 );
and ( n63893 , n62715 , n62783 );
and ( n63894 , n62711 , n62783 );
or ( n63895 , n63892 , n63893 , n63894 );
and ( n63896 , n62707 , n62784 );
and ( n63897 , n62784 , n62967 );
and ( n63898 , n62707 , n62967 );
or ( n63899 , n63896 , n63897 , n63898 );
xor ( n63900 , n63895 , n63899 );
and ( n63901 , n62786 , n62903 );
and ( n63902 , n62903 , n62966 );
and ( n63903 , n62786 , n62966 );
or ( n63904 , n63901 , n63902 , n63903 );
and ( n63905 , n62720 , n62724 );
and ( n63906 , n62724 , n62782 );
and ( n63907 , n62720 , n62782 );
or ( n63908 , n63905 , n63906 , n63907 );
and ( n63909 , n62790 , n62791 );
and ( n63910 , n62791 , n62902 );
and ( n63911 , n62790 , n62902 );
or ( n63912 , n63909 , n63910 , n63911 );
xor ( n63913 , n63908 , n63912 );
and ( n63914 , n62751 , n62755 );
and ( n63915 , n62755 , n62761 );
and ( n63916 , n62751 , n62761 );
or ( n63917 , n63914 , n63915 , n63916 );
and ( n63918 , n62729 , n62733 );
and ( n63919 , n62733 , n62781 );
and ( n63920 , n62729 , n62781 );
or ( n63921 , n63918 , n63919 , n63920 );
xor ( n63922 , n63917 , n63921 );
and ( n63923 , n62738 , n62742 );
and ( n63924 , n62742 , n62780 );
and ( n63925 , n62738 , n62780 );
or ( n63926 , n63923 , n63924 , n63925 );
and ( n63927 , n62800 , n62825 );
and ( n63928 , n62825 , n62863 );
and ( n63929 , n62800 , n62863 );
or ( n63930 , n63927 , n63928 , n63929 );
xor ( n63931 , n63926 , n63930 );
and ( n63932 , n62747 , n62762 );
and ( n63933 , n62762 , n62779 );
and ( n63934 , n62747 , n62779 );
or ( n63935 , n63932 , n63933 , n63934 );
and ( n63936 , n62804 , n62808 );
and ( n63937 , n62808 , n62824 );
and ( n63938 , n62804 , n62824 );
or ( n63939 , n63936 , n63937 , n63938 );
xor ( n63940 , n63935 , n63939 );
and ( n63941 , n62767 , n62772 );
and ( n63942 , n62772 , n62778 );
and ( n63943 , n62767 , n62778 );
or ( n63944 , n63941 , n63942 , n63943 );
and ( n63945 , n62757 , n62758 );
and ( n63946 , n62758 , n62760 );
and ( n63947 , n62757 , n62760 );
or ( n63948 , n63945 , n63946 , n63947 );
and ( n63949 , n62768 , n62769 );
and ( n63950 , n62769 , n62771 );
and ( n63951 , n62768 , n62771 );
or ( n63952 , n63949 , n63950 , n63951 );
xor ( n63953 , n63948 , n63952 );
and ( n63954 , n30695 , n5408 );
and ( n63955 , n31836 , n5103 );
xor ( n63956 , n63954 , n63955 );
and ( n63957 , n32649 , n4730 );
xor ( n63958 , n63956 , n63957 );
xor ( n63959 , n63953 , n63958 );
xor ( n63960 , n63944 , n63959 );
and ( n63961 , n62774 , n62775 );
and ( n63962 , n62775 , n62777 );
and ( n63963 , n62774 , n62777 );
or ( n63964 , n63961 , n63962 , n63963 );
and ( n63965 , n27361 , n6504 );
and ( n63966 , n28456 , n6132 );
xor ( n63967 , n63965 , n63966 );
and ( n63968 , n29559 , n5765 );
xor ( n63969 , n63967 , n63968 );
xor ( n63970 , n63964 , n63969 );
and ( n63971 , n24214 , n7662 );
and ( n63972 , n25243 , n7310 );
xor ( n63973 , n63971 , n63972 );
and ( n63974 , n26296 , n6971 );
xor ( n63975 , n63973 , n63974 );
xor ( n63976 , n63970 , n63975 );
xor ( n63977 , n63960 , n63976 );
xor ( n63978 , n63940 , n63977 );
xor ( n63979 , n63931 , n63978 );
xor ( n63980 , n63922 , n63979 );
xor ( n63981 , n63913 , n63980 );
xor ( n63982 , n63904 , n63981 );
and ( n63983 , n62796 , n62864 );
and ( n63984 , n62864 , n62901 );
and ( n63985 , n62796 , n62901 );
or ( n63986 , n63983 , n63984 , n63985 );
and ( n63987 , n62908 , n62965 );
xor ( n63988 , n63986 , n63987 );
and ( n63989 , n62869 , n62873 );
and ( n63990 , n62873 , n62900 );
and ( n63991 , n62869 , n62900 );
or ( n63992 , n63989 , n63990 , n63991 );
and ( n63993 , n62830 , n62846 );
and ( n63994 , n62846 , n62862 );
and ( n63995 , n62830 , n62862 );
or ( n63996 , n63993 , n63994 , n63995 );
and ( n63997 , n62813 , n62817 );
and ( n63998 , n62817 , n62823 );
and ( n63999 , n62813 , n62823 );
or ( n64000 , n63997 , n63998 , n63999 );
and ( n64001 , n62834 , n62839 );
and ( n64002 , n62839 , n62845 );
and ( n64003 , n62834 , n62845 );
or ( n64004 , n64001 , n64002 , n64003 );
xor ( n64005 , n64000 , n64004 );
and ( n64006 , n62819 , n62820 );
and ( n64007 , n62820 , n62822 );
and ( n64008 , n62819 , n62822 );
or ( n64009 , n64006 , n64007 , n64008 );
and ( n64010 , n62835 , n62836 );
and ( n64011 , n62836 , n62838 );
and ( n64012 , n62835 , n62838 );
or ( n64013 , n64010 , n64011 , n64012 );
xor ( n64014 , n64009 , n64013 );
and ( n64015 , n21216 , n9348 );
and ( n64016 , n22186 , n8669 );
xor ( n64017 , n64015 , n64016 );
and ( n64018 , n22892 , n8243 );
xor ( n64019 , n64017 , n64018 );
xor ( n64020 , n64014 , n64019 );
xor ( n64021 , n64005 , n64020 );
xor ( n64022 , n63996 , n64021 );
and ( n64023 , n62851 , n62855 );
and ( n64024 , n62855 , n62861 );
and ( n64025 , n62851 , n62861 );
or ( n64026 , n64023 , n64024 , n64025 );
and ( n64027 , n62841 , n62842 );
and ( n64028 , n62842 , n62844 );
and ( n64029 , n62841 , n62844 );
or ( n64030 , n64027 , n64028 , n64029 );
and ( n64031 , n18144 , n11718 );
and ( n64032 , n19324 , n10977 );
xor ( n64033 , n64031 , n64032 );
and ( n64034 , n20233 , n10239 );
xor ( n64035 , n64033 , n64034 );
xor ( n64036 , n64030 , n64035 );
and ( n64037 , n15758 , n14044 );
and ( n64038 , n16637 , n13256 );
xor ( n64039 , n64037 , n64038 );
and ( n64040 , n17512 , n12531 );
xor ( n64041 , n64039 , n64040 );
xor ( n64042 , n64036 , n64041 );
xor ( n64043 , n64026 , n64042 );
and ( n64044 , n62857 , n62858 );
and ( n64045 , n62858 , n62860 );
and ( n64046 , n62857 , n62860 );
or ( n64047 , n64044 , n64045 , n64046 );
and ( n64048 , n62888 , n62889 );
and ( n64049 , n62889 , n62891 );
and ( n64050 , n62888 , n62891 );
or ( n64051 , n64048 , n64049 , n64050 );
xor ( n64052 , n64047 , n64051 );
and ( n64053 , n13322 , n16550 );
and ( n64054 , n14118 , n15691 );
xor ( n64055 , n64053 , n64054 );
buf ( n64056 , n14938 );
xor ( n64057 , n64055 , n64056 );
xor ( n64058 , n64052 , n64057 );
xor ( n64059 , n64043 , n64058 );
xor ( n64060 , n64022 , n64059 );
xor ( n64061 , n63992 , n64060 );
and ( n64062 , n62878 , n62882 );
and ( n64063 , n62882 , n62899 );
and ( n64064 , n62878 , n62899 );
or ( n64065 , n64062 , n64063 , n64064 );
and ( n64066 , n62913 , n62928 );
and ( n64067 , n62928 , n62945 );
and ( n64068 , n62913 , n62945 );
or ( n64069 , n64066 , n64067 , n64068 );
xor ( n64070 , n64065 , n64069 );
and ( n64071 , n62887 , n62892 );
and ( n64072 , n62892 , n62898 );
and ( n64073 , n62887 , n62898 );
or ( n64074 , n64071 , n64072 , n64073 );
and ( n64075 , n62917 , n62921 );
and ( n64076 , n62921 , n62927 );
and ( n64077 , n62917 , n62927 );
or ( n64078 , n64075 , n64076 , n64077 );
xor ( n64079 , n64074 , n64078 );
and ( n64080 , n62894 , n62895 );
and ( n64081 , n62895 , n62897 );
and ( n64082 , n62894 , n62897 );
or ( n64083 , n64080 , n64081 , n64082 );
and ( n64084 , n8718 , n22065 );
and ( n64085 , n9400 , n20976 );
xor ( n64086 , n64084 , n64085 );
and ( n64087 , n10291 , n20156 );
xor ( n64088 , n64086 , n64087 );
xor ( n64089 , n64083 , n64088 );
and ( n64090 , n11015 , n19222 );
and ( n64091 , n11769 , n18407 );
xor ( n64092 , n64090 , n64091 );
and ( n64093 , n12320 , n17422 );
xor ( n64094 , n64092 , n64093 );
xor ( n64095 , n64089 , n64094 );
xor ( n64096 , n64079 , n64095 );
xor ( n64097 , n64070 , n64096 );
xor ( n64098 , n64061 , n64097 );
xor ( n64099 , n63988 , n64098 );
and ( n64100 , n62909 , n62946 );
and ( n64101 , n62946 , n62964 );
and ( n64102 , n62909 , n62964 );
or ( n64103 , n64100 , n64101 , n64102 );
and ( n64104 , n62951 , n62963 );
and ( n64105 , n62933 , n62938 );
and ( n64106 , n62938 , n62944 );
and ( n64107 , n62933 , n62944 );
or ( n64108 , n64105 , n64106 , n64107 );
and ( n64109 , n62923 , n62924 );
and ( n64110 , n62924 , n62926 );
and ( n64111 , n62923 , n62926 );
or ( n64112 , n64109 , n64110 , n64111 );
and ( n64113 , n62934 , n62935 );
and ( n64114 , n62935 , n62937 );
and ( n64115 , n62934 , n62937 );
or ( n64116 , n64113 , n64114 , n64115 );
xor ( n64117 , n64112 , n64116 );
and ( n64118 , n7385 , n25163 );
and ( n64119 , n7808 , n24137 );
xor ( n64120 , n64118 , n64119 );
and ( n64121 , n8079 , n23075 );
xor ( n64122 , n64120 , n64121 );
xor ( n64123 , n64117 , n64122 );
xor ( n64124 , n64108 , n64123 );
and ( n64125 , n62940 , n62941 );
and ( n64126 , n62941 , n62943 );
and ( n64127 , n62940 , n62943 );
or ( n64128 , n64125 , n64126 , n64127 );
and ( n64129 , n4959 , n31761 );
and ( n64130 , n5459 , n30629 );
xor ( n64131 , n64129 , n64130 );
and ( n64132 , n5819 , n29508 );
xor ( n64133 , n64131 , n64132 );
xor ( n64134 , n64128 , n64133 );
and ( n64135 , n6187 , n28406 );
and ( n64136 , n6569 , n27296 );
xor ( n64137 , n64135 , n64136 );
and ( n64138 , n6816 , n26216 );
xor ( n64139 , n64137 , n64138 );
xor ( n64140 , n64134 , n64139 );
xor ( n64141 , n64124 , n64140 );
xor ( n64142 , n64104 , n64141 );
and ( n64143 , n62955 , n62962 );
and ( n64144 , n62958 , n62959 );
and ( n64145 , n62959 , n62961 );
and ( n64146 , n62958 , n62961 );
or ( n64147 , n64144 , n64145 , n64146 );
not ( n64148 , n4438 );
and ( n64149 , n34193 , n4438 );
nor ( n64150 , n64148 , n64149 );
and ( n64151 , n4766 , n32999 );
xor ( n64152 , n64150 , n64151 );
xor ( n64153 , n64147 , n64152 );
xor ( n64154 , n64143 , n64153 );
xor ( n64155 , n64142 , n64154 );
xor ( n64156 , n64103 , n64155 );
xor ( n64157 , n64099 , n64156 );
xor ( n64158 , n63982 , n64157 );
xor ( n64159 , n63900 , n64158 );
xor ( n64160 , n63891 , n64159 );
and ( n64161 , n62690 , n62693 );
and ( n64162 , n62693 , n62969 );
and ( n64163 , n62690 , n62969 );
or ( n64164 , n64161 , n64162 , n64163 );
xor ( n64165 , n64160 , n64164 );
and ( n64166 , n62970 , n62974 );
and ( n64167 , n62975 , n62978 );
or ( n64168 , n64166 , n64167 );
xor ( n64169 , n64165 , n64168 );
buf ( n64170 , n64169 );
buf ( n64171 , n64170 );
not ( n64172 , n64171 );
nor ( n64173 , n64172 , n8739 );
xor ( n64174 , n63883 , n64173 );
and ( n64175 , n62686 , n62983 );
and ( n64176 , n62984 , n62987 );
or ( n64177 , n64175 , n64176 );
xor ( n64178 , n64174 , n64177 );
buf ( n64179 , n64178 );
buf ( n64180 , n64179 );
not ( n64181 , n64180 );
buf ( n64182 , n587 );
not ( n64183 , n64182 );
nor ( n64184 , n64181 , n64183 );
xor ( n64185 , n63509 , n64184 );
xor ( n64186 , n62999 , n63506 );
nor ( n64187 , n62991 , n64183 );
and ( n64188 , n64186 , n64187 );
xor ( n64189 , n64186 , n64187 );
xor ( n64190 , n63003 , n63504 );
nor ( n64191 , n61800 , n64183 );
and ( n64192 , n64190 , n64191 );
xor ( n64193 , n64190 , n64191 );
xor ( n64194 , n63007 , n63502 );
nor ( n64195 , n60609 , n64183 );
and ( n64196 , n64194 , n64195 );
xor ( n64197 , n64194 , n64195 );
xor ( n64198 , n63011 , n63500 );
nor ( n64199 , n59421 , n64183 );
and ( n64200 , n64198 , n64199 );
xor ( n64201 , n64198 , n64199 );
xor ( n64202 , n63015 , n63498 );
nor ( n64203 , n58226 , n64183 );
and ( n64204 , n64202 , n64203 );
xor ( n64205 , n64202 , n64203 );
xor ( n64206 , n63019 , n63496 );
nor ( n64207 , n57031 , n64183 );
and ( n64208 , n64206 , n64207 );
xor ( n64209 , n64206 , n64207 );
xor ( n64210 , n63023 , n63494 );
nor ( n64211 , n55835 , n64183 );
and ( n64212 , n64210 , n64211 );
xor ( n64213 , n64210 , n64211 );
xor ( n64214 , n63027 , n63492 );
nor ( n64215 , n54638 , n64183 );
and ( n64216 , n64214 , n64215 );
xor ( n64217 , n64214 , n64215 );
xor ( n64218 , n63031 , n63490 );
nor ( n64219 , n53441 , n64183 );
and ( n64220 , n64218 , n64219 );
xor ( n64221 , n64218 , n64219 );
xor ( n64222 , n63035 , n63488 );
nor ( n64223 , n52247 , n64183 );
and ( n64224 , n64222 , n64223 );
xor ( n64225 , n64222 , n64223 );
xor ( n64226 , n63039 , n63486 );
nor ( n64227 , n51049 , n64183 );
and ( n64228 , n64226 , n64227 );
xor ( n64229 , n64226 , n64227 );
xor ( n64230 , n63043 , n63484 );
nor ( n64231 , n49850 , n64183 );
and ( n64232 , n64230 , n64231 );
xor ( n64233 , n64230 , n64231 );
xor ( n64234 , n63047 , n63482 );
nor ( n64235 , n48650 , n64183 );
and ( n64236 , n64234 , n64235 );
xor ( n64237 , n64234 , n64235 );
xor ( n64238 , n63051 , n63480 );
nor ( n64239 , n47449 , n64183 );
and ( n64240 , n64238 , n64239 );
xor ( n64241 , n64238 , n64239 );
xor ( n64242 , n63055 , n63478 );
nor ( n64243 , n46248 , n64183 );
and ( n64244 , n64242 , n64243 );
xor ( n64245 , n64242 , n64243 );
xor ( n64246 , n63059 , n63476 );
nor ( n64247 , n45047 , n64183 );
and ( n64248 , n64246 , n64247 );
xor ( n64249 , n64246 , n64247 );
xor ( n64250 , n63063 , n63474 );
nor ( n64251 , n43843 , n64183 );
and ( n64252 , n64250 , n64251 );
xor ( n64253 , n64250 , n64251 );
xor ( n64254 , n63067 , n63472 );
nor ( n64255 , n42641 , n64183 );
and ( n64256 , n64254 , n64255 );
xor ( n64257 , n64254 , n64255 );
xor ( n64258 , n63071 , n63470 );
nor ( n64259 , n41437 , n64183 );
and ( n64260 , n64258 , n64259 );
xor ( n64261 , n64258 , n64259 );
xor ( n64262 , n63075 , n63468 );
nor ( n64263 , n40232 , n64183 );
and ( n64264 , n64262 , n64263 );
xor ( n64265 , n64262 , n64263 );
xor ( n64266 , n63079 , n63466 );
nor ( n64267 , n39027 , n64183 );
and ( n64268 , n64266 , n64267 );
xor ( n64269 , n64266 , n64267 );
xor ( n64270 , n63083 , n63464 );
nor ( n64271 , n37825 , n64183 );
and ( n64272 , n64270 , n64271 );
xor ( n64273 , n64270 , n64271 );
xor ( n64274 , n63087 , n63462 );
nor ( n64275 , n36620 , n64183 );
and ( n64276 , n64274 , n64275 );
xor ( n64277 , n64274 , n64275 );
xor ( n64278 , n63091 , n63460 );
nor ( n64279 , n35419 , n64183 );
and ( n64280 , n64278 , n64279 );
xor ( n64281 , n64278 , n64279 );
xor ( n64282 , n63095 , n63458 );
nor ( n64283 , n34224 , n64183 );
and ( n64284 , n64282 , n64283 );
xor ( n64285 , n64282 , n64283 );
xor ( n64286 , n63099 , n63456 );
nor ( n64287 , n33033 , n64183 );
and ( n64288 , n64286 , n64287 );
xor ( n64289 , n64286 , n64287 );
xor ( n64290 , n63103 , n63454 );
nor ( n64291 , n31867 , n64183 );
and ( n64292 , n64290 , n64291 );
xor ( n64293 , n64290 , n64291 );
xor ( n64294 , n63107 , n63452 );
nor ( n64295 , n30725 , n64183 );
and ( n64296 , n64294 , n64295 );
xor ( n64297 , n64294 , n64295 );
xor ( n64298 , n63111 , n63450 );
nor ( n64299 , n29596 , n64183 );
and ( n64300 , n64298 , n64299 );
xor ( n64301 , n64298 , n64299 );
xor ( n64302 , n63115 , n63448 );
nor ( n64303 , n28487 , n64183 );
and ( n64304 , n64302 , n64303 );
xor ( n64305 , n64302 , n64303 );
xor ( n64306 , n63119 , n63446 );
nor ( n64307 , n27397 , n64183 );
and ( n64308 , n64306 , n64307 );
xor ( n64309 , n64306 , n64307 );
xor ( n64310 , n63123 , n63444 );
nor ( n64311 , n26326 , n64183 );
and ( n64312 , n64310 , n64311 );
xor ( n64313 , n64310 , n64311 );
xor ( n64314 , n63127 , n63442 );
nor ( n64315 , n25272 , n64183 );
and ( n64316 , n64314 , n64315 );
xor ( n64317 , n64314 , n64315 );
xor ( n64318 , n63131 , n63440 );
nor ( n64319 , n24242 , n64183 );
and ( n64320 , n64318 , n64319 );
xor ( n64321 , n64318 , n64319 );
xor ( n64322 , n63135 , n63438 );
nor ( n64323 , n23225 , n64183 );
and ( n64324 , n64322 , n64323 );
xor ( n64325 , n64322 , n64323 );
xor ( n64326 , n63139 , n63436 );
nor ( n64327 , n22231 , n64183 );
and ( n64328 , n64326 , n64327 );
xor ( n64329 , n64326 , n64327 );
xor ( n64330 , n63143 , n63434 );
nor ( n64331 , n21258 , n64183 );
and ( n64332 , n64330 , n64331 );
xor ( n64333 , n64330 , n64331 );
xor ( n64334 , n63147 , n63432 );
nor ( n64335 , n20303 , n64183 );
and ( n64336 , n64334 , n64335 );
xor ( n64337 , n64334 , n64335 );
xor ( n64338 , n63151 , n63430 );
nor ( n64339 , n19365 , n64183 );
and ( n64340 , n64338 , n64339 );
xor ( n64341 , n64338 , n64339 );
xor ( n64342 , n63155 , n63428 );
nor ( n64343 , n18448 , n64183 );
and ( n64344 , n64342 , n64343 );
xor ( n64345 , n64342 , n64343 );
xor ( n64346 , n63159 , n63426 );
nor ( n64347 , n17548 , n64183 );
and ( n64348 , n64346 , n64347 );
xor ( n64349 , n64346 , n64347 );
xor ( n64350 , n63163 , n63424 );
nor ( n64351 , n16669 , n64183 );
and ( n64352 , n64350 , n64351 );
xor ( n64353 , n64350 , n64351 );
xor ( n64354 , n63167 , n63422 );
nor ( n64355 , n15809 , n64183 );
and ( n64356 , n64354 , n64355 );
xor ( n64357 , n64354 , n64355 );
xor ( n64358 , n63171 , n63420 );
nor ( n64359 , n14968 , n64183 );
and ( n64360 , n64358 , n64359 );
xor ( n64361 , n64358 , n64359 );
xor ( n64362 , n63175 , n63418 );
nor ( n64363 , n14147 , n64183 );
and ( n64364 , n64362 , n64363 );
xor ( n64365 , n64362 , n64363 );
xor ( n64366 , n63179 , n63416 );
nor ( n64367 , n13349 , n64183 );
and ( n64368 , n64366 , n64367 );
xor ( n64369 , n64366 , n64367 );
xor ( n64370 , n63183 , n63414 );
nor ( n64371 , n12564 , n64183 );
and ( n64372 , n64370 , n64371 );
xor ( n64373 , n64370 , n64371 );
xor ( n64374 , n63187 , n63412 );
nor ( n64375 , n11799 , n64183 );
and ( n64376 , n64374 , n64375 );
xor ( n64377 , n64374 , n64375 );
xor ( n64378 , n63191 , n63410 );
nor ( n64379 , n11050 , n64183 );
and ( n64380 , n64378 , n64379 );
xor ( n64381 , n64378 , n64379 );
xor ( n64382 , n63195 , n63408 );
nor ( n64383 , n10321 , n64183 );
and ( n64384 , n64382 , n64383 );
xor ( n64385 , n64382 , n64383 );
xor ( n64386 , n63199 , n63406 );
nor ( n64387 , n9429 , n64183 );
and ( n64388 , n64386 , n64387 );
xor ( n64389 , n64386 , n64387 );
xor ( n64390 , n63203 , n63404 );
nor ( n64391 , n8949 , n64183 );
and ( n64392 , n64390 , n64391 );
xor ( n64393 , n64390 , n64391 );
xor ( n64394 , n63207 , n63402 );
nor ( n64395 , n9437 , n64183 );
and ( n64396 , n64394 , n64395 );
xor ( n64397 , n64394 , n64395 );
xor ( n64398 , n63211 , n63400 );
nor ( n64399 , n9446 , n64183 );
and ( n64400 , n64398 , n64399 );
xor ( n64401 , n64398 , n64399 );
xor ( n64402 , n63215 , n63398 );
nor ( n64403 , n9455 , n64183 );
and ( n64404 , n64402 , n64403 );
xor ( n64405 , n64402 , n64403 );
xor ( n64406 , n63219 , n63396 );
nor ( n64407 , n9464 , n64183 );
and ( n64408 , n64406 , n64407 );
xor ( n64409 , n64406 , n64407 );
xor ( n64410 , n63223 , n63394 );
nor ( n64411 , n9473 , n64183 );
and ( n64412 , n64410 , n64411 );
xor ( n64413 , n64410 , n64411 );
xor ( n64414 , n63227 , n63392 );
nor ( n64415 , n9482 , n64183 );
and ( n64416 , n64414 , n64415 );
xor ( n64417 , n64414 , n64415 );
xor ( n64418 , n63231 , n63390 );
nor ( n64419 , n9491 , n64183 );
and ( n64420 , n64418 , n64419 );
xor ( n64421 , n64418 , n64419 );
xor ( n64422 , n63235 , n63388 );
nor ( n64423 , n9500 , n64183 );
and ( n64424 , n64422 , n64423 );
xor ( n64425 , n64422 , n64423 );
xor ( n64426 , n63239 , n63386 );
nor ( n64427 , n9509 , n64183 );
and ( n64428 , n64426 , n64427 );
xor ( n64429 , n64426 , n64427 );
xor ( n64430 , n63243 , n63384 );
nor ( n64431 , n9518 , n64183 );
and ( n64432 , n64430 , n64431 );
xor ( n64433 , n64430 , n64431 );
xor ( n64434 , n63247 , n63382 );
nor ( n64435 , n9527 , n64183 );
and ( n64436 , n64434 , n64435 );
xor ( n64437 , n64434 , n64435 );
xor ( n64438 , n63251 , n63380 );
nor ( n64439 , n9536 , n64183 );
and ( n64440 , n64438 , n64439 );
xor ( n64441 , n64438 , n64439 );
xor ( n64442 , n63255 , n63378 );
nor ( n64443 , n9545 , n64183 );
and ( n64444 , n64442 , n64443 );
xor ( n64445 , n64442 , n64443 );
xor ( n64446 , n63259 , n63376 );
nor ( n64447 , n9554 , n64183 );
and ( n64448 , n64446 , n64447 );
xor ( n64449 , n64446 , n64447 );
xor ( n64450 , n63263 , n63374 );
nor ( n64451 , n9563 , n64183 );
and ( n64452 , n64450 , n64451 );
xor ( n64453 , n64450 , n64451 );
xor ( n64454 , n63267 , n63372 );
nor ( n64455 , n9572 , n64183 );
and ( n64456 , n64454 , n64455 );
xor ( n64457 , n64454 , n64455 );
xor ( n64458 , n63271 , n63370 );
nor ( n64459 , n9581 , n64183 );
and ( n64460 , n64458 , n64459 );
xor ( n64461 , n64458 , n64459 );
xor ( n64462 , n63275 , n63368 );
nor ( n64463 , n9590 , n64183 );
and ( n64464 , n64462 , n64463 );
xor ( n64465 , n64462 , n64463 );
xor ( n64466 , n63279 , n63366 );
nor ( n64467 , n9599 , n64183 );
and ( n64468 , n64466 , n64467 );
xor ( n64469 , n64466 , n64467 );
xor ( n64470 , n63283 , n63364 );
nor ( n64471 , n9608 , n64183 );
and ( n64472 , n64470 , n64471 );
xor ( n64473 , n64470 , n64471 );
xor ( n64474 , n63287 , n63362 );
nor ( n64475 , n9617 , n64183 );
and ( n64476 , n64474 , n64475 );
xor ( n64477 , n64474 , n64475 );
xor ( n64478 , n63291 , n63360 );
nor ( n64479 , n9626 , n64183 );
and ( n64480 , n64478 , n64479 );
xor ( n64481 , n64478 , n64479 );
xor ( n64482 , n63295 , n63358 );
nor ( n64483 , n9635 , n64183 );
and ( n64484 , n64482 , n64483 );
xor ( n64485 , n64482 , n64483 );
xor ( n64486 , n63299 , n63356 );
nor ( n64487 , n9644 , n64183 );
and ( n64488 , n64486 , n64487 );
xor ( n64489 , n64486 , n64487 );
xor ( n64490 , n63303 , n63354 );
nor ( n64491 , n9653 , n64183 );
and ( n64492 , n64490 , n64491 );
xor ( n64493 , n64490 , n64491 );
xor ( n64494 , n63307 , n63352 );
nor ( n64495 , n9662 , n64183 );
and ( n64496 , n64494 , n64495 );
xor ( n64497 , n64494 , n64495 );
xor ( n64498 , n63311 , n63350 );
nor ( n64499 , n9671 , n64183 );
and ( n64500 , n64498 , n64499 );
xor ( n64501 , n64498 , n64499 );
xor ( n64502 , n63315 , n63348 );
nor ( n64503 , n9680 , n64183 );
and ( n64504 , n64502 , n64503 );
xor ( n64505 , n64502 , n64503 );
xor ( n64506 , n63319 , n63346 );
nor ( n64507 , n9689 , n64183 );
and ( n64508 , n64506 , n64507 );
xor ( n64509 , n64506 , n64507 );
xor ( n64510 , n63323 , n63344 );
nor ( n64511 , n9698 , n64183 );
and ( n64512 , n64510 , n64511 );
xor ( n64513 , n64510 , n64511 );
xor ( n64514 , n63327 , n63342 );
nor ( n64515 , n9707 , n64183 );
and ( n64516 , n64514 , n64515 );
xor ( n64517 , n64514 , n64515 );
xor ( n64518 , n63331 , n63340 );
nor ( n64519 , n9716 , n64183 );
and ( n64520 , n64518 , n64519 );
xor ( n64521 , n64518 , n64519 );
xor ( n64522 , n63335 , n63338 );
nor ( n64523 , n9725 , n64183 );
and ( n64524 , n64522 , n64523 );
xor ( n64525 , n64522 , n64523 );
xor ( n64526 , n63336 , n63337 );
nor ( n64527 , n9734 , n64183 );
and ( n64528 , n64526 , n64527 );
xor ( n64529 , n64526 , n64527 );
nor ( n64530 , n9752 , n62993 );
nor ( n64531 , n9743 , n64183 );
and ( n64532 , n64530 , n64531 );
and ( n64533 , n64529 , n64532 );
or ( n64534 , n64528 , n64533 );
and ( n64535 , n64525 , n64534 );
or ( n64536 , n64524 , n64535 );
and ( n64537 , n64521 , n64536 );
or ( n64538 , n64520 , n64537 );
and ( n64539 , n64517 , n64538 );
or ( n64540 , n64516 , n64539 );
and ( n64541 , n64513 , n64540 );
or ( n64542 , n64512 , n64541 );
and ( n64543 , n64509 , n64542 );
or ( n64544 , n64508 , n64543 );
and ( n64545 , n64505 , n64544 );
or ( n64546 , n64504 , n64545 );
and ( n64547 , n64501 , n64546 );
or ( n64548 , n64500 , n64547 );
and ( n64549 , n64497 , n64548 );
or ( n64550 , n64496 , n64549 );
and ( n64551 , n64493 , n64550 );
or ( n64552 , n64492 , n64551 );
and ( n64553 , n64489 , n64552 );
or ( n64554 , n64488 , n64553 );
and ( n64555 , n64485 , n64554 );
or ( n64556 , n64484 , n64555 );
and ( n64557 , n64481 , n64556 );
or ( n64558 , n64480 , n64557 );
and ( n64559 , n64477 , n64558 );
or ( n64560 , n64476 , n64559 );
and ( n64561 , n64473 , n64560 );
or ( n64562 , n64472 , n64561 );
and ( n64563 , n64469 , n64562 );
or ( n64564 , n64468 , n64563 );
and ( n64565 , n64465 , n64564 );
or ( n64566 , n64464 , n64565 );
and ( n64567 , n64461 , n64566 );
or ( n64568 , n64460 , n64567 );
and ( n64569 , n64457 , n64568 );
or ( n64570 , n64456 , n64569 );
and ( n64571 , n64453 , n64570 );
or ( n64572 , n64452 , n64571 );
and ( n64573 , n64449 , n64572 );
or ( n64574 , n64448 , n64573 );
and ( n64575 , n64445 , n64574 );
or ( n64576 , n64444 , n64575 );
and ( n64577 , n64441 , n64576 );
or ( n64578 , n64440 , n64577 );
and ( n64579 , n64437 , n64578 );
or ( n64580 , n64436 , n64579 );
and ( n64581 , n64433 , n64580 );
or ( n64582 , n64432 , n64581 );
and ( n64583 , n64429 , n64582 );
or ( n64584 , n64428 , n64583 );
and ( n64585 , n64425 , n64584 );
or ( n64586 , n64424 , n64585 );
and ( n64587 , n64421 , n64586 );
or ( n64588 , n64420 , n64587 );
and ( n64589 , n64417 , n64588 );
or ( n64590 , n64416 , n64589 );
and ( n64591 , n64413 , n64590 );
or ( n64592 , n64412 , n64591 );
and ( n64593 , n64409 , n64592 );
or ( n64594 , n64408 , n64593 );
and ( n64595 , n64405 , n64594 );
or ( n64596 , n64404 , n64595 );
and ( n64597 , n64401 , n64596 );
or ( n64598 , n64400 , n64597 );
and ( n64599 , n64397 , n64598 );
or ( n64600 , n64396 , n64599 );
and ( n64601 , n64393 , n64600 );
or ( n64602 , n64392 , n64601 );
and ( n64603 , n64389 , n64602 );
or ( n64604 , n64388 , n64603 );
and ( n64605 , n64385 , n64604 );
or ( n64606 , n64384 , n64605 );
and ( n64607 , n64381 , n64606 );
or ( n64608 , n64380 , n64607 );
and ( n64609 , n64377 , n64608 );
or ( n64610 , n64376 , n64609 );
and ( n64611 , n64373 , n64610 );
or ( n64612 , n64372 , n64611 );
and ( n64613 , n64369 , n64612 );
or ( n64614 , n64368 , n64613 );
and ( n64615 , n64365 , n64614 );
or ( n64616 , n64364 , n64615 );
and ( n64617 , n64361 , n64616 );
or ( n64618 , n64360 , n64617 );
and ( n64619 , n64357 , n64618 );
or ( n64620 , n64356 , n64619 );
and ( n64621 , n64353 , n64620 );
or ( n64622 , n64352 , n64621 );
and ( n64623 , n64349 , n64622 );
or ( n64624 , n64348 , n64623 );
and ( n64625 , n64345 , n64624 );
or ( n64626 , n64344 , n64625 );
and ( n64627 , n64341 , n64626 );
or ( n64628 , n64340 , n64627 );
and ( n64629 , n64337 , n64628 );
or ( n64630 , n64336 , n64629 );
and ( n64631 , n64333 , n64630 );
or ( n64632 , n64332 , n64631 );
and ( n64633 , n64329 , n64632 );
or ( n64634 , n64328 , n64633 );
and ( n64635 , n64325 , n64634 );
or ( n64636 , n64324 , n64635 );
and ( n64637 , n64321 , n64636 );
or ( n64638 , n64320 , n64637 );
and ( n64639 , n64317 , n64638 );
or ( n64640 , n64316 , n64639 );
and ( n64641 , n64313 , n64640 );
or ( n64642 , n64312 , n64641 );
and ( n64643 , n64309 , n64642 );
or ( n64644 , n64308 , n64643 );
and ( n64645 , n64305 , n64644 );
or ( n64646 , n64304 , n64645 );
and ( n64647 , n64301 , n64646 );
or ( n64648 , n64300 , n64647 );
and ( n64649 , n64297 , n64648 );
or ( n64650 , n64296 , n64649 );
and ( n64651 , n64293 , n64650 );
or ( n64652 , n64292 , n64651 );
and ( n64653 , n64289 , n64652 );
or ( n64654 , n64288 , n64653 );
and ( n64655 , n64285 , n64654 );
or ( n64656 , n64284 , n64655 );
and ( n64657 , n64281 , n64656 );
or ( n64658 , n64280 , n64657 );
and ( n64659 , n64277 , n64658 );
or ( n64660 , n64276 , n64659 );
and ( n64661 , n64273 , n64660 );
or ( n64662 , n64272 , n64661 );
and ( n64663 , n64269 , n64662 );
or ( n64664 , n64268 , n64663 );
and ( n64665 , n64265 , n64664 );
or ( n64666 , n64264 , n64665 );
and ( n64667 , n64261 , n64666 );
or ( n64668 , n64260 , n64667 );
and ( n64669 , n64257 , n64668 );
or ( n64670 , n64256 , n64669 );
and ( n64671 , n64253 , n64670 );
or ( n64672 , n64252 , n64671 );
and ( n64673 , n64249 , n64672 );
or ( n64674 , n64248 , n64673 );
and ( n64675 , n64245 , n64674 );
or ( n64676 , n64244 , n64675 );
and ( n64677 , n64241 , n64676 );
or ( n64678 , n64240 , n64677 );
and ( n64679 , n64237 , n64678 );
or ( n64680 , n64236 , n64679 );
and ( n64681 , n64233 , n64680 );
or ( n64682 , n64232 , n64681 );
and ( n64683 , n64229 , n64682 );
or ( n64684 , n64228 , n64683 );
and ( n64685 , n64225 , n64684 );
or ( n64686 , n64224 , n64685 );
and ( n64687 , n64221 , n64686 );
or ( n64688 , n64220 , n64687 );
and ( n64689 , n64217 , n64688 );
or ( n64690 , n64216 , n64689 );
and ( n64691 , n64213 , n64690 );
or ( n64692 , n64212 , n64691 );
and ( n64693 , n64209 , n64692 );
or ( n64694 , n64208 , n64693 );
and ( n64695 , n64205 , n64694 );
or ( n64696 , n64204 , n64695 );
and ( n64697 , n64201 , n64696 );
or ( n64698 , n64200 , n64697 );
and ( n64699 , n64197 , n64698 );
or ( n64700 , n64196 , n64699 );
and ( n64701 , n64193 , n64700 );
or ( n64702 , n64192 , n64701 );
and ( n64703 , n64189 , n64702 );
or ( n64704 , n64188 , n64703 );
xor ( n64705 , n64185 , n64704 );
and ( n64706 , n33403 , n4785 );
nor ( n64707 , n4786 , n64706 );
nor ( n64708 , n5126 , n32231 );
xor ( n64709 , n64707 , n64708 );
and ( n64710 , n63511 , n63512 );
and ( n64711 , n63513 , n63516 );
or ( n64712 , n64710 , n64711 );
xor ( n64713 , n64709 , n64712 );
nor ( n64714 , n5477 , n31083 );
xor ( n64715 , n64713 , n64714 );
and ( n64716 , n63517 , n63518 );
and ( n64717 , n63519 , n63522 );
or ( n64718 , n64716 , n64717 );
xor ( n64719 , n64715 , n64718 );
nor ( n64720 , n5838 , n29948 );
xor ( n64721 , n64719 , n64720 );
and ( n64722 , n63523 , n63524 );
and ( n64723 , n63525 , n63528 );
or ( n64724 , n64722 , n64723 );
xor ( n64725 , n64721 , n64724 );
nor ( n64726 , n6212 , n28833 );
xor ( n64727 , n64725 , n64726 );
and ( n64728 , n63529 , n63530 );
and ( n64729 , n63531 , n63534 );
or ( n64730 , n64728 , n64729 );
xor ( n64731 , n64727 , n64730 );
nor ( n64732 , n6596 , n27737 );
xor ( n64733 , n64731 , n64732 );
and ( n64734 , n63535 , n63536 );
and ( n64735 , n63537 , n63540 );
or ( n64736 , n64734 , n64735 );
xor ( n64737 , n64733 , n64736 );
nor ( n64738 , n6997 , n26660 );
xor ( n64739 , n64737 , n64738 );
and ( n64740 , n63541 , n63542 );
and ( n64741 , n63543 , n63546 );
or ( n64742 , n64740 , n64741 );
xor ( n64743 , n64739 , n64742 );
nor ( n64744 , n7413 , n25600 );
xor ( n64745 , n64743 , n64744 );
and ( n64746 , n63547 , n63548 );
and ( n64747 , n63549 , n63552 );
or ( n64748 , n64746 , n64747 );
xor ( n64749 , n64745 , n64748 );
nor ( n64750 , n7841 , n24564 );
xor ( n64751 , n64749 , n64750 );
and ( n64752 , n63553 , n63554 );
and ( n64753 , n63555 , n63558 );
or ( n64754 , n64752 , n64753 );
xor ( n64755 , n64751 , n64754 );
nor ( n64756 , n8281 , n23541 );
xor ( n64757 , n64755 , n64756 );
and ( n64758 , n63559 , n63560 );
and ( n64759 , n63561 , n63564 );
or ( n64760 , n64758 , n64759 );
xor ( n64761 , n64757 , n64760 );
nor ( n64762 , n8737 , n22541 );
xor ( n64763 , n64761 , n64762 );
and ( n64764 , n63565 , n63566 );
and ( n64765 , n63567 , n63570 );
or ( n64766 , n64764 , n64765 );
xor ( n64767 , n64763 , n64766 );
nor ( n64768 , n9420 , n21562 );
xor ( n64769 , n64767 , n64768 );
and ( n64770 , n63571 , n63572 );
and ( n64771 , n63573 , n63576 );
or ( n64772 , n64770 , n64771 );
xor ( n64773 , n64769 , n64772 );
nor ( n64774 , n10312 , n20601 );
xor ( n64775 , n64773 , n64774 );
and ( n64776 , n63577 , n63578 );
and ( n64777 , n63579 , n63582 );
or ( n64778 , n64776 , n64777 );
xor ( n64779 , n64775 , n64778 );
nor ( n64780 , n11041 , n19657 );
xor ( n64781 , n64779 , n64780 );
and ( n64782 , n63583 , n63584 );
and ( n64783 , n63585 , n63588 );
or ( n64784 , n64782 , n64783 );
xor ( n64785 , n64781 , n64784 );
nor ( n64786 , n11790 , n18734 );
xor ( n64787 , n64785 , n64786 );
and ( n64788 , n63589 , n63590 );
and ( n64789 , n63591 , n63594 );
or ( n64790 , n64788 , n64789 );
xor ( n64791 , n64787 , n64790 );
nor ( n64792 , n12555 , n17828 );
xor ( n64793 , n64791 , n64792 );
and ( n64794 , n63595 , n63596 );
and ( n64795 , n63597 , n63600 );
or ( n64796 , n64794 , n64795 );
xor ( n64797 , n64793 , n64796 );
nor ( n64798 , n13340 , n16943 );
xor ( n64799 , n64797 , n64798 );
and ( n64800 , n63601 , n63602 );
and ( n64801 , n63603 , n63606 );
or ( n64802 , n64800 , n64801 );
xor ( n64803 , n64799 , n64802 );
nor ( n64804 , n14138 , n16077 );
xor ( n64805 , n64803 , n64804 );
and ( n64806 , n63607 , n63608 );
and ( n64807 , n63609 , n63612 );
or ( n64808 , n64806 , n64807 );
xor ( n64809 , n64805 , n64808 );
nor ( n64810 , n14959 , n15230 );
xor ( n64811 , n64809 , n64810 );
and ( n64812 , n63613 , n63614 );
and ( n64813 , n63615 , n63618 );
or ( n64814 , n64812 , n64813 );
xor ( n64815 , n64811 , n64814 );
nor ( n64816 , n15800 , n14403 );
xor ( n64817 , n64815 , n64816 );
and ( n64818 , n63619 , n63620 );
and ( n64819 , n63621 , n63624 );
or ( n64820 , n64818 , n64819 );
xor ( n64821 , n64817 , n64820 );
nor ( n64822 , n16660 , n13599 );
xor ( n64823 , n64821 , n64822 );
and ( n64824 , n63625 , n63626 );
and ( n64825 , n63627 , n63630 );
or ( n64826 , n64824 , n64825 );
xor ( n64827 , n64823 , n64826 );
nor ( n64828 , n17539 , n12808 );
xor ( n64829 , n64827 , n64828 );
and ( n64830 , n63631 , n63632 );
and ( n64831 , n63633 , n63636 );
or ( n64832 , n64830 , n64831 );
xor ( n64833 , n64829 , n64832 );
nor ( n64834 , n18439 , n12037 );
xor ( n64835 , n64833 , n64834 );
and ( n64836 , n63637 , n63638 );
and ( n64837 , n63639 , n63642 );
or ( n64838 , n64836 , n64837 );
xor ( n64839 , n64835 , n64838 );
nor ( n64840 , n19356 , n11282 );
xor ( n64841 , n64839 , n64840 );
and ( n64842 , n63643 , n63644 );
and ( n64843 , n63645 , n63648 );
or ( n64844 , n64842 , n64843 );
xor ( n64845 , n64841 , n64844 );
nor ( n64846 , n20294 , n10547 );
xor ( n64847 , n64845 , n64846 );
and ( n64848 , n63649 , n63650 );
and ( n64849 , n63651 , n63654 );
or ( n64850 , n64848 , n64849 );
xor ( n64851 , n64847 , n64850 );
nor ( n64852 , n21249 , n9829 );
xor ( n64853 , n64851 , n64852 );
and ( n64854 , n63655 , n63656 );
and ( n64855 , n63657 , n63660 );
or ( n64856 , n64854 , n64855 );
xor ( n64857 , n64853 , n64856 );
nor ( n64858 , n22222 , n8955 );
xor ( n64859 , n64857 , n64858 );
and ( n64860 , n63661 , n63662 );
and ( n64861 , n63663 , n63666 );
or ( n64862 , n64860 , n64861 );
xor ( n64863 , n64859 , n64862 );
nor ( n64864 , n23216 , n603 );
xor ( n64865 , n64863 , n64864 );
and ( n64866 , n63667 , n63668 );
and ( n64867 , n63669 , n63672 );
or ( n64868 , n64866 , n64867 );
xor ( n64869 , n64865 , n64868 );
nor ( n64870 , n24233 , n652 );
xor ( n64871 , n64869 , n64870 );
and ( n64872 , n63673 , n63674 );
and ( n64873 , n63675 , n63678 );
or ( n64874 , n64872 , n64873 );
xor ( n64875 , n64871 , n64874 );
nor ( n64876 , n25263 , n624 );
xor ( n64877 , n64875 , n64876 );
and ( n64878 , n63679 , n63680 );
and ( n64879 , n63681 , n63684 );
or ( n64880 , n64878 , n64879 );
xor ( n64881 , n64877 , n64880 );
nor ( n64882 , n26317 , n648 );
xor ( n64883 , n64881 , n64882 );
and ( n64884 , n63685 , n63686 );
and ( n64885 , n63687 , n63690 );
or ( n64886 , n64884 , n64885 );
xor ( n64887 , n64883 , n64886 );
nor ( n64888 , n27388 , n686 );
xor ( n64889 , n64887 , n64888 );
and ( n64890 , n63691 , n63692 );
and ( n64891 , n63693 , n63696 );
or ( n64892 , n64890 , n64891 );
xor ( n64893 , n64889 , n64892 );
nor ( n64894 , n28478 , n735 );
xor ( n64895 , n64893 , n64894 );
and ( n64896 , n63697 , n63698 );
and ( n64897 , n63699 , n63702 );
or ( n64898 , n64896 , n64897 );
xor ( n64899 , n64895 , n64898 );
nor ( n64900 , n29587 , n798 );
xor ( n64901 , n64899 , n64900 );
and ( n64902 , n63703 , n63704 );
and ( n64903 , n63705 , n63708 );
or ( n64904 , n64902 , n64903 );
xor ( n64905 , n64901 , n64904 );
nor ( n64906 , n30716 , n870 );
xor ( n64907 , n64905 , n64906 );
and ( n64908 , n63709 , n63710 );
and ( n64909 , n63711 , n63714 );
or ( n64910 , n64908 , n64909 );
xor ( n64911 , n64907 , n64910 );
nor ( n64912 , n31858 , n960 );
xor ( n64913 , n64911 , n64912 );
and ( n64914 , n63715 , n63716 );
and ( n64915 , n63717 , n63720 );
or ( n64916 , n64914 , n64915 );
xor ( n64917 , n64913 , n64916 );
nor ( n64918 , n33024 , n1064 );
xor ( n64919 , n64917 , n64918 );
and ( n64920 , n63721 , n63722 );
and ( n64921 , n63723 , n63726 );
or ( n64922 , n64920 , n64921 );
xor ( n64923 , n64919 , n64922 );
nor ( n64924 , n34215 , n1178 );
xor ( n64925 , n64923 , n64924 );
and ( n64926 , n63727 , n63728 );
and ( n64927 , n63729 , n63732 );
or ( n64928 , n64926 , n64927 );
xor ( n64929 , n64925 , n64928 );
nor ( n64930 , n35410 , n1305 );
xor ( n64931 , n64929 , n64930 );
and ( n64932 , n63733 , n63734 );
and ( n64933 , n63735 , n63738 );
or ( n64934 , n64932 , n64933 );
xor ( n64935 , n64931 , n64934 );
nor ( n64936 , n36611 , n1447 );
xor ( n64937 , n64935 , n64936 );
and ( n64938 , n63739 , n63740 );
and ( n64939 , n63741 , n63744 );
or ( n64940 , n64938 , n64939 );
xor ( n64941 , n64937 , n64940 );
nor ( n64942 , n37816 , n1600 );
xor ( n64943 , n64941 , n64942 );
and ( n64944 , n63745 , n63746 );
and ( n64945 , n63747 , n63750 );
or ( n64946 , n64944 , n64945 );
xor ( n64947 , n64943 , n64946 );
nor ( n64948 , n39018 , n1768 );
xor ( n64949 , n64947 , n64948 );
and ( n64950 , n63751 , n63752 );
and ( n64951 , n63753 , n63756 );
or ( n64952 , n64950 , n64951 );
xor ( n64953 , n64949 , n64952 );
nor ( n64954 , n40223 , n1947 );
xor ( n64955 , n64953 , n64954 );
and ( n64956 , n63757 , n63758 );
and ( n64957 , n63759 , n63762 );
or ( n64958 , n64956 , n64957 );
xor ( n64959 , n64955 , n64958 );
nor ( n64960 , n41428 , n2139 );
xor ( n64961 , n64959 , n64960 );
and ( n64962 , n63763 , n63764 );
and ( n64963 , n63765 , n63768 );
or ( n64964 , n64962 , n64963 );
xor ( n64965 , n64961 , n64964 );
nor ( n64966 , n42632 , n2345 );
xor ( n64967 , n64965 , n64966 );
and ( n64968 , n63769 , n63770 );
and ( n64969 , n63771 , n63774 );
or ( n64970 , n64968 , n64969 );
xor ( n64971 , n64967 , n64970 );
nor ( n64972 , n43834 , n2568 );
xor ( n64973 , n64971 , n64972 );
and ( n64974 , n63775 , n63776 );
and ( n64975 , n63777 , n63780 );
or ( n64976 , n64974 , n64975 );
xor ( n64977 , n64973 , n64976 );
nor ( n64978 , n45038 , n2799 );
xor ( n64979 , n64977 , n64978 );
and ( n64980 , n63781 , n63782 );
and ( n64981 , n63783 , n63786 );
or ( n64982 , n64980 , n64981 );
xor ( n64983 , n64979 , n64982 );
nor ( n64984 , n46239 , n3045 );
xor ( n64985 , n64983 , n64984 );
and ( n64986 , n63787 , n63788 );
and ( n64987 , n63789 , n63792 );
or ( n64988 , n64986 , n64987 );
xor ( n64989 , n64985 , n64988 );
nor ( n64990 , n47440 , n3302 );
xor ( n64991 , n64989 , n64990 );
and ( n64992 , n63793 , n63794 );
and ( n64993 , n63795 , n63798 );
or ( n64994 , n64992 , n64993 );
xor ( n64995 , n64991 , n64994 );
nor ( n64996 , n48641 , n3572 );
xor ( n64997 , n64995 , n64996 );
and ( n64998 , n63799 , n63800 );
and ( n64999 , n63801 , n63804 );
or ( n65000 , n64998 , n64999 );
xor ( n65001 , n64997 , n65000 );
nor ( n65002 , n49841 , n3855 );
xor ( n65003 , n65001 , n65002 );
and ( n65004 , n63805 , n63806 );
and ( n65005 , n63807 , n63810 );
or ( n65006 , n65004 , n65005 );
xor ( n65007 , n65003 , n65006 );
nor ( n65008 , n51040 , n4153 );
xor ( n65009 , n65007 , n65008 );
and ( n65010 , n63811 , n63812 );
and ( n65011 , n63813 , n63816 );
or ( n65012 , n65010 , n65011 );
xor ( n65013 , n65009 , n65012 );
nor ( n65014 , n52238 , n4460 );
xor ( n65015 , n65013 , n65014 );
and ( n65016 , n63817 , n63818 );
and ( n65017 , n63819 , n63822 );
or ( n65018 , n65016 , n65017 );
xor ( n65019 , n65015 , n65018 );
nor ( n65020 , n53432 , n4788 );
xor ( n65021 , n65019 , n65020 );
and ( n65022 , n63823 , n63824 );
and ( n65023 , n63825 , n63828 );
or ( n65024 , n65022 , n65023 );
xor ( n65025 , n65021 , n65024 );
nor ( n65026 , n54629 , n5128 );
xor ( n65027 , n65025 , n65026 );
and ( n65028 , n63829 , n63830 );
and ( n65029 , n63831 , n63834 );
or ( n65030 , n65028 , n65029 );
xor ( n65031 , n65027 , n65030 );
nor ( n65032 , n55826 , n5479 );
xor ( n65033 , n65031 , n65032 );
and ( n65034 , n63835 , n63836 );
and ( n65035 , n63837 , n63840 );
or ( n65036 , n65034 , n65035 );
xor ( n65037 , n65033 , n65036 );
nor ( n65038 , n57022 , n5840 );
xor ( n65039 , n65037 , n65038 );
and ( n65040 , n63841 , n63842 );
and ( n65041 , n63843 , n63846 );
or ( n65042 , n65040 , n65041 );
xor ( n65043 , n65039 , n65042 );
nor ( n65044 , n58217 , n6214 );
xor ( n65045 , n65043 , n65044 );
and ( n65046 , n63847 , n63848 );
and ( n65047 , n63849 , n63852 );
or ( n65048 , n65046 , n65047 );
xor ( n65049 , n65045 , n65048 );
nor ( n65050 , n59412 , n6598 );
xor ( n65051 , n65049 , n65050 );
and ( n65052 , n63853 , n63854 );
and ( n65053 , n63855 , n63858 );
or ( n65054 , n65052 , n65053 );
xor ( n65055 , n65051 , n65054 );
nor ( n65056 , n60600 , n6999 );
xor ( n65057 , n65055 , n65056 );
and ( n65058 , n63859 , n63860 );
and ( n65059 , n63861 , n63864 );
or ( n65060 , n65058 , n65059 );
xor ( n65061 , n65057 , n65060 );
nor ( n65062 , n61791 , n7415 );
xor ( n65063 , n65061 , n65062 );
and ( n65064 , n63865 , n63866 );
and ( n65065 , n63867 , n63870 );
or ( n65066 , n65064 , n65065 );
xor ( n65067 , n65063 , n65066 );
nor ( n65068 , n62982 , n7843 );
xor ( n65069 , n65067 , n65068 );
and ( n65070 , n63871 , n63872 );
and ( n65071 , n63873 , n63876 );
or ( n65072 , n65070 , n65071 );
xor ( n65073 , n65069 , n65072 );
nor ( n65074 , n64172 , n8283 );
xor ( n65075 , n65073 , n65074 );
and ( n65076 , n63877 , n63878 );
and ( n65077 , n63879 , n63882 );
or ( n65078 , n65076 , n65077 );
xor ( n65079 , n65075 , n65078 );
and ( n65080 , n63895 , n63899 );
and ( n65081 , n63899 , n64158 );
and ( n65082 , n63895 , n64158 );
or ( n65083 , n65080 , n65081 , n65082 );
and ( n65084 , n33774 , n4730 );
not ( n65085 , n4730 );
nor ( n65086 , n65084 , n65085 );
xor ( n65087 , n65083 , n65086 );
and ( n65088 , n63908 , n63912 );
and ( n65089 , n63912 , n63980 );
and ( n65090 , n63908 , n63980 );
or ( n65091 , n65088 , n65089 , n65090 );
and ( n65092 , n63904 , n63981 );
and ( n65093 , n63981 , n64157 );
and ( n65094 , n63904 , n64157 );
or ( n65095 , n65092 , n65093 , n65094 );
xor ( n65096 , n65091 , n65095 );
and ( n65097 , n64099 , n64156 );
and ( n65098 , n63986 , n63987 );
and ( n65099 , n63987 , n64098 );
and ( n65100 , n63986 , n64098 );
or ( n65101 , n65098 , n65099 , n65100 );
and ( n65102 , n63917 , n63921 );
and ( n65103 , n63921 , n63979 );
and ( n65104 , n63917 , n63979 );
or ( n65105 , n65102 , n65103 , n65104 );
xor ( n65106 , n65101 , n65105 );
and ( n65107 , n63948 , n63952 );
and ( n65108 , n63952 , n63958 );
and ( n65109 , n63948 , n63958 );
or ( n65110 , n65107 , n65108 , n65109 );
and ( n65111 , n63926 , n63930 );
and ( n65112 , n63930 , n63978 );
and ( n65113 , n63926 , n63978 );
or ( n65114 , n65111 , n65112 , n65113 );
xor ( n65115 , n65110 , n65114 );
and ( n65116 , n63935 , n63939 );
and ( n65117 , n63939 , n63977 );
and ( n65118 , n63935 , n63977 );
or ( n65119 , n65116 , n65117 , n65118 );
and ( n65120 , n63996 , n64021 );
and ( n65121 , n64021 , n64059 );
and ( n65122 , n63996 , n64059 );
or ( n65123 , n65120 , n65121 , n65122 );
xor ( n65124 , n65119 , n65123 );
and ( n65125 , n63944 , n63959 );
and ( n65126 , n63959 , n63976 );
and ( n65127 , n63944 , n63976 );
or ( n65128 , n65125 , n65126 , n65127 );
and ( n65129 , n64000 , n64004 );
and ( n65130 , n64004 , n64020 );
and ( n65131 , n64000 , n64020 );
or ( n65132 , n65129 , n65130 , n65131 );
xor ( n65133 , n65128 , n65132 );
and ( n65134 , n63964 , n63969 );
and ( n65135 , n63969 , n63975 );
and ( n65136 , n63964 , n63975 );
or ( n65137 , n65134 , n65135 , n65136 );
and ( n65138 , n63954 , n63955 );
and ( n65139 , n63955 , n63957 );
and ( n65140 , n63954 , n63957 );
or ( n65141 , n65138 , n65139 , n65140 );
and ( n65142 , n63965 , n63966 );
and ( n65143 , n63966 , n63968 );
and ( n65144 , n63965 , n63968 );
or ( n65145 , n65142 , n65143 , n65144 );
xor ( n65146 , n65141 , n65145 );
and ( n65147 , n30695 , n5765 );
and ( n65148 , n31836 , n5408 );
xor ( n65149 , n65147 , n65148 );
and ( n65150 , n32649 , n5103 );
xor ( n65151 , n65149 , n65150 );
xor ( n65152 , n65146 , n65151 );
xor ( n65153 , n65137 , n65152 );
and ( n65154 , n63971 , n63972 );
and ( n65155 , n63972 , n63974 );
and ( n65156 , n63971 , n63974 );
or ( n65157 , n65154 , n65155 , n65156 );
and ( n65158 , n27361 , n6971 );
and ( n65159 , n28456 , n6504 );
xor ( n65160 , n65158 , n65159 );
and ( n65161 , n29559 , n6132 );
xor ( n65162 , n65160 , n65161 );
xor ( n65163 , n65157 , n65162 );
and ( n65164 , n24214 , n8243 );
and ( n65165 , n25243 , n7662 );
xor ( n65166 , n65164 , n65165 );
and ( n65167 , n26296 , n7310 );
xor ( n65168 , n65166 , n65167 );
xor ( n65169 , n65163 , n65168 );
xor ( n65170 , n65153 , n65169 );
xor ( n65171 , n65133 , n65170 );
xor ( n65172 , n65124 , n65171 );
xor ( n65173 , n65115 , n65172 );
xor ( n65174 , n65106 , n65173 );
xor ( n65175 , n65097 , n65174 );
and ( n65176 , n63992 , n64060 );
and ( n65177 , n64060 , n64097 );
and ( n65178 , n63992 , n64097 );
or ( n65179 , n65176 , n65177 , n65178 );
and ( n65180 , n64103 , n64155 );
xor ( n65181 , n65179 , n65180 );
and ( n65182 , n64065 , n64069 );
and ( n65183 , n64069 , n64096 );
and ( n65184 , n64065 , n64096 );
or ( n65185 , n65182 , n65183 , n65184 );
and ( n65186 , n64026 , n64042 );
and ( n65187 , n64042 , n64058 );
and ( n65188 , n64026 , n64058 );
or ( n65189 , n65186 , n65187 , n65188 );
and ( n65190 , n64009 , n64013 );
and ( n65191 , n64013 , n64019 );
and ( n65192 , n64009 , n64019 );
or ( n65193 , n65190 , n65191 , n65192 );
and ( n65194 , n64030 , n64035 );
and ( n65195 , n64035 , n64041 );
and ( n65196 , n64030 , n64041 );
or ( n65197 , n65194 , n65195 , n65196 );
xor ( n65198 , n65193 , n65197 );
and ( n65199 , n64015 , n64016 );
and ( n65200 , n64016 , n64018 );
and ( n65201 , n64015 , n64018 );
or ( n65202 , n65199 , n65200 , n65201 );
and ( n65203 , n64031 , n64032 );
and ( n65204 , n64032 , n64034 );
and ( n65205 , n64031 , n64034 );
or ( n65206 , n65203 , n65204 , n65205 );
xor ( n65207 , n65202 , n65206 );
and ( n65208 , n21216 , n10239 );
and ( n65209 , n22186 , n9348 );
xor ( n65210 , n65208 , n65209 );
and ( n65211 , n22892 , n8669 );
xor ( n65212 , n65210 , n65211 );
xor ( n65213 , n65207 , n65212 );
xor ( n65214 , n65198 , n65213 );
xor ( n65215 , n65189 , n65214 );
and ( n65216 , n64047 , n64051 );
and ( n65217 , n64051 , n64057 );
and ( n65218 , n64047 , n64057 );
or ( n65219 , n65216 , n65217 , n65218 );
and ( n65220 , n64037 , n64038 );
and ( n65221 , n64038 , n64040 );
and ( n65222 , n64037 , n64040 );
or ( n65223 , n65220 , n65221 , n65222 );
and ( n65224 , n18144 , n12531 );
and ( n65225 , n19324 , n11718 );
xor ( n65226 , n65224 , n65225 );
and ( n65227 , n20233 , n10977 );
xor ( n65228 , n65226 , n65227 );
xor ( n65229 , n65223 , n65228 );
and ( n65230 , n15758 , n14838 );
and ( n65231 , n16637 , n14044 );
xor ( n65232 , n65230 , n65231 );
and ( n65233 , n17512 , n13256 );
xor ( n65234 , n65232 , n65233 );
xor ( n65235 , n65229 , n65234 );
xor ( n65236 , n65219 , n65235 );
and ( n65237 , n64090 , n64091 );
and ( n65238 , n64091 , n64093 );
and ( n65239 , n64090 , n64093 );
or ( n65240 , n65237 , n65238 , n65239 );
and ( n65241 , n64053 , n64054 );
and ( n65242 , n64054 , n64056 );
and ( n65243 , n64053 , n64056 );
or ( n65244 , n65241 , n65242 , n65243 );
xor ( n65245 , n65240 , n65244 );
and ( n65246 , n13322 , n17422 );
and ( n65247 , n14118 , n16550 );
xor ( n65248 , n65246 , n65247 );
and ( n65249 , n14938 , n15691 );
xor ( n65250 , n65248 , n65249 );
xor ( n65251 , n65245 , n65250 );
xor ( n65252 , n65236 , n65251 );
xor ( n65253 , n65215 , n65252 );
xor ( n65254 , n65185 , n65253 );
and ( n65255 , n64074 , n64078 );
and ( n65256 , n64078 , n64095 );
and ( n65257 , n64074 , n64095 );
or ( n65258 , n65255 , n65256 , n65257 );
and ( n65259 , n64108 , n64123 );
and ( n65260 , n64123 , n64140 );
and ( n65261 , n64108 , n64140 );
or ( n65262 , n65259 , n65260 , n65261 );
xor ( n65263 , n65258 , n65262 );
and ( n65264 , n64083 , n64088 );
and ( n65265 , n64088 , n64094 );
and ( n65266 , n64083 , n64094 );
or ( n65267 , n65264 , n65265 , n65266 );
and ( n65268 , n64112 , n64116 );
and ( n65269 , n64116 , n64122 );
and ( n65270 , n64112 , n64122 );
or ( n65271 , n65268 , n65269 , n65270 );
xor ( n65272 , n65267 , n65271 );
and ( n65273 , n64084 , n64085 );
and ( n65274 , n64085 , n64087 );
and ( n65275 , n64084 , n64087 );
or ( n65276 , n65273 , n65274 , n65275 );
and ( n65277 , n11015 , n20156 );
and ( n65278 , n11769 , n19222 );
xor ( n65279 , n65277 , n65278 );
and ( n65280 , n12320 , n18407 );
xor ( n65281 , n65279 , n65280 );
xor ( n65282 , n65276 , n65281 );
and ( n65283 , n8718 , n23075 );
and ( n65284 , n9400 , n22065 );
xor ( n65285 , n65283 , n65284 );
and ( n65286 , n10291 , n20976 );
xor ( n65287 , n65285 , n65286 );
xor ( n65288 , n65282 , n65287 );
xor ( n65289 , n65272 , n65288 );
xor ( n65290 , n65263 , n65289 );
xor ( n65291 , n65254 , n65290 );
xor ( n65292 , n65181 , n65291 );
and ( n65293 , n64104 , n64141 );
and ( n65294 , n64141 , n64154 );
and ( n65295 , n64104 , n64154 );
or ( n65296 , n65293 , n65294 , n65295 );
and ( n65297 , n64143 , n64153 );
and ( n65298 , n64128 , n64133 );
and ( n65299 , n64133 , n64139 );
and ( n65300 , n64128 , n64139 );
or ( n65301 , n65298 , n65299 , n65300 );
and ( n65302 , n64135 , n64136 );
and ( n65303 , n64136 , n64138 );
and ( n65304 , n64135 , n64138 );
or ( n65305 , n65302 , n65303 , n65304 );
and ( n65306 , n64118 , n64119 );
and ( n65307 , n64119 , n64121 );
and ( n65308 , n64118 , n64121 );
or ( n65309 , n65306 , n65307 , n65308 );
xor ( n65310 , n65305 , n65309 );
and ( n65311 , n7385 , n26216 );
and ( n65312 , n7808 , n25163 );
xor ( n65313 , n65311 , n65312 );
and ( n65314 , n8079 , n24137 );
xor ( n65315 , n65313 , n65314 );
xor ( n65316 , n65310 , n65315 );
xor ( n65317 , n65301 , n65316 );
and ( n65318 , n64129 , n64130 );
and ( n65319 , n64130 , n64132 );
and ( n65320 , n64129 , n64132 );
or ( n65321 , n65318 , n65319 , n65320 );
and ( n65322 , n6187 , n29508 );
and ( n65323 , n6569 , n28406 );
xor ( n65324 , n65322 , n65323 );
and ( n65325 , n6816 , n27296 );
xor ( n65326 , n65324 , n65325 );
xor ( n65327 , n65321 , n65326 );
and ( n65328 , n4959 , n32999 );
and ( n65329 , n5459 , n31761 );
xor ( n65330 , n65328 , n65329 );
and ( n65331 , n5819 , n30629 );
xor ( n65332 , n65330 , n65331 );
xor ( n65333 , n65327 , n65332 );
xor ( n65334 , n65317 , n65333 );
xor ( n65335 , n65297 , n65334 );
and ( n65336 , n64147 , n64152 );
and ( n65337 , n64150 , n64151 );
not ( n65338 , n4766 );
and ( n65339 , n34193 , n4766 );
nor ( n65340 , n65338 , n65339 );
xor ( n65341 , n65337 , n65340 );
xor ( n65342 , n65336 , n65341 );
xor ( n65343 , n65335 , n65342 );
xor ( n65344 , n65296 , n65343 );
xor ( n65345 , n65292 , n65344 );
xor ( n65346 , n65175 , n65345 );
xor ( n65347 , n65096 , n65346 );
xor ( n65348 , n65087 , n65347 );
and ( n65349 , n63887 , n63890 );
and ( n65350 , n63890 , n64159 );
and ( n65351 , n63887 , n64159 );
or ( n65352 , n65349 , n65350 , n65351 );
xor ( n65353 , n65348 , n65352 );
and ( n65354 , n64160 , n64164 );
and ( n65355 , n64165 , n64168 );
or ( n65356 , n65354 , n65355 );
xor ( n65357 , n65353 , n65356 );
buf ( n65358 , n65357 );
buf ( n65359 , n65358 );
not ( n65360 , n65359 );
nor ( n65361 , n65360 , n8739 );
xor ( n65362 , n65079 , n65361 );
and ( n65363 , n63883 , n64173 );
and ( n65364 , n64174 , n64177 );
or ( n65365 , n65363 , n65364 );
xor ( n65366 , n65362 , n65365 );
buf ( n65367 , n65366 );
buf ( n65368 , n65367 );
not ( n65369 , n65368 );
buf ( n65370 , n588 );
not ( n65371 , n65370 );
nor ( n65372 , n65369 , n65371 );
xor ( n65373 , n64705 , n65372 );
xor ( n65374 , n64189 , n64702 );
nor ( n65375 , n64181 , n65371 );
and ( n65376 , n65374 , n65375 );
xor ( n65377 , n65374 , n65375 );
xor ( n65378 , n64193 , n64700 );
nor ( n65379 , n62991 , n65371 );
and ( n65380 , n65378 , n65379 );
xor ( n65381 , n65378 , n65379 );
xor ( n65382 , n64197 , n64698 );
nor ( n65383 , n61800 , n65371 );
and ( n65384 , n65382 , n65383 );
xor ( n65385 , n65382 , n65383 );
xor ( n65386 , n64201 , n64696 );
nor ( n65387 , n60609 , n65371 );
and ( n65388 , n65386 , n65387 );
xor ( n65389 , n65386 , n65387 );
xor ( n65390 , n64205 , n64694 );
nor ( n65391 , n59421 , n65371 );
and ( n65392 , n65390 , n65391 );
xor ( n65393 , n65390 , n65391 );
xor ( n65394 , n64209 , n64692 );
nor ( n65395 , n58226 , n65371 );
and ( n65396 , n65394 , n65395 );
xor ( n65397 , n65394 , n65395 );
xor ( n65398 , n64213 , n64690 );
nor ( n65399 , n57031 , n65371 );
and ( n65400 , n65398 , n65399 );
xor ( n65401 , n65398 , n65399 );
xor ( n65402 , n64217 , n64688 );
nor ( n65403 , n55835 , n65371 );
and ( n65404 , n65402 , n65403 );
xor ( n65405 , n65402 , n65403 );
xor ( n65406 , n64221 , n64686 );
nor ( n65407 , n54638 , n65371 );
and ( n65408 , n65406 , n65407 );
xor ( n65409 , n65406 , n65407 );
xor ( n65410 , n64225 , n64684 );
nor ( n65411 , n53441 , n65371 );
and ( n65412 , n65410 , n65411 );
xor ( n65413 , n65410 , n65411 );
xor ( n65414 , n64229 , n64682 );
nor ( n65415 , n52247 , n65371 );
and ( n65416 , n65414 , n65415 );
xor ( n65417 , n65414 , n65415 );
xor ( n65418 , n64233 , n64680 );
nor ( n65419 , n51049 , n65371 );
and ( n65420 , n65418 , n65419 );
xor ( n65421 , n65418 , n65419 );
xor ( n65422 , n64237 , n64678 );
nor ( n65423 , n49850 , n65371 );
and ( n65424 , n65422 , n65423 );
xor ( n65425 , n65422 , n65423 );
xor ( n65426 , n64241 , n64676 );
nor ( n65427 , n48650 , n65371 );
and ( n65428 , n65426 , n65427 );
xor ( n65429 , n65426 , n65427 );
xor ( n65430 , n64245 , n64674 );
nor ( n65431 , n47449 , n65371 );
and ( n65432 , n65430 , n65431 );
xor ( n65433 , n65430 , n65431 );
xor ( n65434 , n64249 , n64672 );
nor ( n65435 , n46248 , n65371 );
and ( n65436 , n65434 , n65435 );
xor ( n65437 , n65434 , n65435 );
xor ( n65438 , n64253 , n64670 );
nor ( n65439 , n45047 , n65371 );
and ( n65440 , n65438 , n65439 );
xor ( n65441 , n65438 , n65439 );
xor ( n65442 , n64257 , n64668 );
nor ( n65443 , n43843 , n65371 );
and ( n65444 , n65442 , n65443 );
xor ( n65445 , n65442 , n65443 );
xor ( n65446 , n64261 , n64666 );
nor ( n65447 , n42641 , n65371 );
and ( n65448 , n65446 , n65447 );
xor ( n65449 , n65446 , n65447 );
xor ( n65450 , n64265 , n64664 );
nor ( n65451 , n41437 , n65371 );
and ( n65452 , n65450 , n65451 );
xor ( n65453 , n65450 , n65451 );
xor ( n65454 , n64269 , n64662 );
nor ( n65455 , n40232 , n65371 );
and ( n65456 , n65454 , n65455 );
xor ( n65457 , n65454 , n65455 );
xor ( n65458 , n64273 , n64660 );
nor ( n65459 , n39027 , n65371 );
and ( n65460 , n65458 , n65459 );
xor ( n65461 , n65458 , n65459 );
xor ( n65462 , n64277 , n64658 );
nor ( n65463 , n37825 , n65371 );
and ( n65464 , n65462 , n65463 );
xor ( n65465 , n65462 , n65463 );
xor ( n65466 , n64281 , n64656 );
nor ( n65467 , n36620 , n65371 );
and ( n65468 , n65466 , n65467 );
xor ( n65469 , n65466 , n65467 );
xor ( n65470 , n64285 , n64654 );
nor ( n65471 , n35419 , n65371 );
and ( n65472 , n65470 , n65471 );
xor ( n65473 , n65470 , n65471 );
xor ( n65474 , n64289 , n64652 );
nor ( n65475 , n34224 , n65371 );
and ( n65476 , n65474 , n65475 );
xor ( n65477 , n65474 , n65475 );
xor ( n65478 , n64293 , n64650 );
nor ( n65479 , n33033 , n65371 );
and ( n65480 , n65478 , n65479 );
xor ( n65481 , n65478 , n65479 );
xor ( n65482 , n64297 , n64648 );
nor ( n65483 , n31867 , n65371 );
and ( n65484 , n65482 , n65483 );
xor ( n65485 , n65482 , n65483 );
xor ( n65486 , n64301 , n64646 );
nor ( n65487 , n30725 , n65371 );
and ( n65488 , n65486 , n65487 );
xor ( n65489 , n65486 , n65487 );
xor ( n65490 , n64305 , n64644 );
nor ( n65491 , n29596 , n65371 );
and ( n65492 , n65490 , n65491 );
xor ( n65493 , n65490 , n65491 );
xor ( n65494 , n64309 , n64642 );
nor ( n65495 , n28487 , n65371 );
and ( n65496 , n65494 , n65495 );
xor ( n65497 , n65494 , n65495 );
xor ( n65498 , n64313 , n64640 );
nor ( n65499 , n27397 , n65371 );
and ( n65500 , n65498 , n65499 );
xor ( n65501 , n65498 , n65499 );
xor ( n65502 , n64317 , n64638 );
nor ( n65503 , n26326 , n65371 );
and ( n65504 , n65502 , n65503 );
xor ( n65505 , n65502 , n65503 );
xor ( n65506 , n64321 , n64636 );
nor ( n65507 , n25272 , n65371 );
and ( n65508 , n65506 , n65507 );
xor ( n65509 , n65506 , n65507 );
xor ( n65510 , n64325 , n64634 );
nor ( n65511 , n24242 , n65371 );
and ( n65512 , n65510 , n65511 );
xor ( n65513 , n65510 , n65511 );
xor ( n65514 , n64329 , n64632 );
nor ( n65515 , n23225 , n65371 );
and ( n65516 , n65514 , n65515 );
xor ( n65517 , n65514 , n65515 );
xor ( n65518 , n64333 , n64630 );
nor ( n65519 , n22231 , n65371 );
and ( n65520 , n65518 , n65519 );
xor ( n65521 , n65518 , n65519 );
xor ( n65522 , n64337 , n64628 );
nor ( n65523 , n21258 , n65371 );
and ( n65524 , n65522 , n65523 );
xor ( n65525 , n65522 , n65523 );
xor ( n65526 , n64341 , n64626 );
nor ( n65527 , n20303 , n65371 );
and ( n65528 , n65526 , n65527 );
xor ( n65529 , n65526 , n65527 );
xor ( n65530 , n64345 , n64624 );
nor ( n65531 , n19365 , n65371 );
and ( n65532 , n65530 , n65531 );
xor ( n65533 , n65530 , n65531 );
xor ( n65534 , n64349 , n64622 );
nor ( n65535 , n18448 , n65371 );
and ( n65536 , n65534 , n65535 );
xor ( n65537 , n65534 , n65535 );
xor ( n65538 , n64353 , n64620 );
nor ( n65539 , n17548 , n65371 );
and ( n65540 , n65538 , n65539 );
xor ( n65541 , n65538 , n65539 );
xor ( n65542 , n64357 , n64618 );
nor ( n65543 , n16669 , n65371 );
and ( n65544 , n65542 , n65543 );
xor ( n65545 , n65542 , n65543 );
xor ( n65546 , n64361 , n64616 );
nor ( n65547 , n15809 , n65371 );
and ( n65548 , n65546 , n65547 );
xor ( n65549 , n65546 , n65547 );
xor ( n65550 , n64365 , n64614 );
nor ( n65551 , n14968 , n65371 );
and ( n65552 , n65550 , n65551 );
xor ( n65553 , n65550 , n65551 );
xor ( n65554 , n64369 , n64612 );
nor ( n65555 , n14147 , n65371 );
and ( n65556 , n65554 , n65555 );
xor ( n65557 , n65554 , n65555 );
xor ( n65558 , n64373 , n64610 );
nor ( n65559 , n13349 , n65371 );
and ( n65560 , n65558 , n65559 );
xor ( n65561 , n65558 , n65559 );
xor ( n65562 , n64377 , n64608 );
nor ( n65563 , n12564 , n65371 );
and ( n65564 , n65562 , n65563 );
xor ( n65565 , n65562 , n65563 );
xor ( n65566 , n64381 , n64606 );
nor ( n65567 , n11799 , n65371 );
and ( n65568 , n65566 , n65567 );
xor ( n65569 , n65566 , n65567 );
xor ( n65570 , n64385 , n64604 );
nor ( n65571 , n11050 , n65371 );
and ( n65572 , n65570 , n65571 );
xor ( n65573 , n65570 , n65571 );
xor ( n65574 , n64389 , n64602 );
nor ( n65575 , n10321 , n65371 );
and ( n65576 , n65574 , n65575 );
xor ( n65577 , n65574 , n65575 );
xor ( n65578 , n64393 , n64600 );
nor ( n65579 , n9429 , n65371 );
and ( n65580 , n65578 , n65579 );
xor ( n65581 , n65578 , n65579 );
xor ( n65582 , n64397 , n64598 );
nor ( n65583 , n8949 , n65371 );
and ( n65584 , n65582 , n65583 );
xor ( n65585 , n65582 , n65583 );
xor ( n65586 , n64401 , n64596 );
nor ( n65587 , n9437 , n65371 );
and ( n65588 , n65586 , n65587 );
xor ( n65589 , n65586 , n65587 );
xor ( n65590 , n64405 , n64594 );
nor ( n65591 , n9446 , n65371 );
and ( n65592 , n65590 , n65591 );
xor ( n65593 , n65590 , n65591 );
xor ( n65594 , n64409 , n64592 );
nor ( n65595 , n9455 , n65371 );
and ( n65596 , n65594 , n65595 );
xor ( n65597 , n65594 , n65595 );
xor ( n65598 , n64413 , n64590 );
nor ( n65599 , n9464 , n65371 );
and ( n65600 , n65598 , n65599 );
xor ( n65601 , n65598 , n65599 );
xor ( n65602 , n64417 , n64588 );
nor ( n65603 , n9473 , n65371 );
and ( n65604 , n65602 , n65603 );
xor ( n65605 , n65602 , n65603 );
xor ( n65606 , n64421 , n64586 );
nor ( n65607 , n9482 , n65371 );
and ( n65608 , n65606 , n65607 );
xor ( n65609 , n65606 , n65607 );
xor ( n65610 , n64425 , n64584 );
nor ( n65611 , n9491 , n65371 );
and ( n65612 , n65610 , n65611 );
xor ( n65613 , n65610 , n65611 );
xor ( n65614 , n64429 , n64582 );
nor ( n65615 , n9500 , n65371 );
and ( n65616 , n65614 , n65615 );
xor ( n65617 , n65614 , n65615 );
xor ( n65618 , n64433 , n64580 );
nor ( n65619 , n9509 , n65371 );
and ( n65620 , n65618 , n65619 );
xor ( n65621 , n65618 , n65619 );
xor ( n65622 , n64437 , n64578 );
nor ( n65623 , n9518 , n65371 );
and ( n65624 , n65622 , n65623 );
xor ( n65625 , n65622 , n65623 );
xor ( n65626 , n64441 , n64576 );
nor ( n65627 , n9527 , n65371 );
and ( n65628 , n65626 , n65627 );
xor ( n65629 , n65626 , n65627 );
xor ( n65630 , n64445 , n64574 );
nor ( n65631 , n9536 , n65371 );
and ( n65632 , n65630 , n65631 );
xor ( n65633 , n65630 , n65631 );
xor ( n65634 , n64449 , n64572 );
nor ( n65635 , n9545 , n65371 );
and ( n65636 , n65634 , n65635 );
xor ( n65637 , n65634 , n65635 );
xor ( n65638 , n64453 , n64570 );
nor ( n65639 , n9554 , n65371 );
and ( n65640 , n65638 , n65639 );
xor ( n65641 , n65638 , n65639 );
xor ( n65642 , n64457 , n64568 );
nor ( n65643 , n9563 , n65371 );
and ( n65644 , n65642 , n65643 );
xor ( n65645 , n65642 , n65643 );
xor ( n65646 , n64461 , n64566 );
nor ( n65647 , n9572 , n65371 );
and ( n65648 , n65646 , n65647 );
xor ( n65649 , n65646 , n65647 );
xor ( n65650 , n64465 , n64564 );
nor ( n65651 , n9581 , n65371 );
and ( n65652 , n65650 , n65651 );
xor ( n65653 , n65650 , n65651 );
xor ( n65654 , n64469 , n64562 );
nor ( n65655 , n9590 , n65371 );
and ( n65656 , n65654 , n65655 );
xor ( n65657 , n65654 , n65655 );
xor ( n65658 , n64473 , n64560 );
nor ( n65659 , n9599 , n65371 );
and ( n65660 , n65658 , n65659 );
xor ( n65661 , n65658 , n65659 );
xor ( n65662 , n64477 , n64558 );
nor ( n65663 , n9608 , n65371 );
and ( n65664 , n65662 , n65663 );
xor ( n65665 , n65662 , n65663 );
xor ( n65666 , n64481 , n64556 );
nor ( n65667 , n9617 , n65371 );
and ( n65668 , n65666 , n65667 );
xor ( n65669 , n65666 , n65667 );
xor ( n65670 , n64485 , n64554 );
nor ( n65671 , n9626 , n65371 );
and ( n65672 , n65670 , n65671 );
xor ( n65673 , n65670 , n65671 );
xor ( n65674 , n64489 , n64552 );
nor ( n65675 , n9635 , n65371 );
and ( n65676 , n65674 , n65675 );
xor ( n65677 , n65674 , n65675 );
xor ( n65678 , n64493 , n64550 );
nor ( n65679 , n9644 , n65371 );
and ( n65680 , n65678 , n65679 );
xor ( n65681 , n65678 , n65679 );
xor ( n65682 , n64497 , n64548 );
nor ( n65683 , n9653 , n65371 );
and ( n65684 , n65682 , n65683 );
xor ( n65685 , n65682 , n65683 );
xor ( n65686 , n64501 , n64546 );
nor ( n65687 , n9662 , n65371 );
and ( n65688 , n65686 , n65687 );
xor ( n65689 , n65686 , n65687 );
xor ( n65690 , n64505 , n64544 );
nor ( n65691 , n9671 , n65371 );
and ( n65692 , n65690 , n65691 );
xor ( n65693 , n65690 , n65691 );
xor ( n65694 , n64509 , n64542 );
nor ( n65695 , n9680 , n65371 );
and ( n65696 , n65694 , n65695 );
xor ( n65697 , n65694 , n65695 );
xor ( n65698 , n64513 , n64540 );
nor ( n65699 , n9689 , n65371 );
and ( n65700 , n65698 , n65699 );
xor ( n65701 , n65698 , n65699 );
xor ( n65702 , n64517 , n64538 );
nor ( n65703 , n9698 , n65371 );
and ( n65704 , n65702 , n65703 );
xor ( n65705 , n65702 , n65703 );
xor ( n65706 , n64521 , n64536 );
nor ( n65707 , n9707 , n65371 );
and ( n65708 , n65706 , n65707 );
xor ( n65709 , n65706 , n65707 );
xor ( n65710 , n64525 , n64534 );
nor ( n65711 , n9716 , n65371 );
and ( n65712 , n65710 , n65711 );
xor ( n65713 , n65710 , n65711 );
xor ( n65714 , n64529 , n64532 );
nor ( n65715 , n9725 , n65371 );
and ( n65716 , n65714 , n65715 );
xor ( n65717 , n65714 , n65715 );
xor ( n65718 , n64530 , n64531 );
nor ( n65719 , n9734 , n65371 );
and ( n65720 , n65718 , n65719 );
xor ( n65721 , n65718 , n65719 );
nor ( n65722 , n9752 , n64183 );
nor ( n65723 , n9743 , n65371 );
and ( n65724 , n65722 , n65723 );
and ( n65725 , n65721 , n65724 );
or ( n65726 , n65720 , n65725 );
and ( n65727 , n65717 , n65726 );
or ( n65728 , n65716 , n65727 );
and ( n65729 , n65713 , n65728 );
or ( n65730 , n65712 , n65729 );
and ( n65731 , n65709 , n65730 );
or ( n65732 , n65708 , n65731 );
and ( n65733 , n65705 , n65732 );
or ( n65734 , n65704 , n65733 );
and ( n65735 , n65701 , n65734 );
or ( n65736 , n65700 , n65735 );
and ( n65737 , n65697 , n65736 );
or ( n65738 , n65696 , n65737 );
and ( n65739 , n65693 , n65738 );
or ( n65740 , n65692 , n65739 );
and ( n65741 , n65689 , n65740 );
or ( n65742 , n65688 , n65741 );
and ( n65743 , n65685 , n65742 );
or ( n65744 , n65684 , n65743 );
and ( n65745 , n65681 , n65744 );
or ( n65746 , n65680 , n65745 );
and ( n65747 , n65677 , n65746 );
or ( n65748 , n65676 , n65747 );
and ( n65749 , n65673 , n65748 );
or ( n65750 , n65672 , n65749 );
and ( n65751 , n65669 , n65750 );
or ( n65752 , n65668 , n65751 );
and ( n65753 , n65665 , n65752 );
or ( n65754 , n65664 , n65753 );
and ( n65755 , n65661 , n65754 );
or ( n65756 , n65660 , n65755 );
and ( n65757 , n65657 , n65756 );
or ( n65758 , n65656 , n65757 );
and ( n65759 , n65653 , n65758 );
or ( n65760 , n65652 , n65759 );
and ( n65761 , n65649 , n65760 );
or ( n65762 , n65648 , n65761 );
and ( n65763 , n65645 , n65762 );
or ( n65764 , n65644 , n65763 );
and ( n65765 , n65641 , n65764 );
or ( n65766 , n65640 , n65765 );
and ( n65767 , n65637 , n65766 );
or ( n65768 , n65636 , n65767 );
and ( n65769 , n65633 , n65768 );
or ( n65770 , n65632 , n65769 );
and ( n65771 , n65629 , n65770 );
or ( n65772 , n65628 , n65771 );
and ( n65773 , n65625 , n65772 );
or ( n65774 , n65624 , n65773 );
and ( n65775 , n65621 , n65774 );
or ( n65776 , n65620 , n65775 );
and ( n65777 , n65617 , n65776 );
or ( n65778 , n65616 , n65777 );
and ( n65779 , n65613 , n65778 );
or ( n65780 , n65612 , n65779 );
and ( n65781 , n65609 , n65780 );
or ( n65782 , n65608 , n65781 );
and ( n65783 , n65605 , n65782 );
or ( n65784 , n65604 , n65783 );
and ( n65785 , n65601 , n65784 );
or ( n65786 , n65600 , n65785 );
and ( n65787 , n65597 , n65786 );
or ( n65788 , n65596 , n65787 );
and ( n65789 , n65593 , n65788 );
or ( n65790 , n65592 , n65789 );
and ( n65791 , n65589 , n65790 );
or ( n65792 , n65588 , n65791 );
and ( n65793 , n65585 , n65792 );
or ( n65794 , n65584 , n65793 );
and ( n65795 , n65581 , n65794 );
or ( n65796 , n65580 , n65795 );
and ( n65797 , n65577 , n65796 );
or ( n65798 , n65576 , n65797 );
and ( n65799 , n65573 , n65798 );
or ( n65800 , n65572 , n65799 );
and ( n65801 , n65569 , n65800 );
or ( n65802 , n65568 , n65801 );
and ( n65803 , n65565 , n65802 );
or ( n65804 , n65564 , n65803 );
and ( n65805 , n65561 , n65804 );
or ( n65806 , n65560 , n65805 );
and ( n65807 , n65557 , n65806 );
or ( n65808 , n65556 , n65807 );
and ( n65809 , n65553 , n65808 );
or ( n65810 , n65552 , n65809 );
and ( n65811 , n65549 , n65810 );
or ( n65812 , n65548 , n65811 );
and ( n65813 , n65545 , n65812 );
or ( n65814 , n65544 , n65813 );
and ( n65815 , n65541 , n65814 );
or ( n65816 , n65540 , n65815 );
and ( n65817 , n65537 , n65816 );
or ( n65818 , n65536 , n65817 );
and ( n65819 , n65533 , n65818 );
or ( n65820 , n65532 , n65819 );
and ( n65821 , n65529 , n65820 );
or ( n65822 , n65528 , n65821 );
and ( n65823 , n65525 , n65822 );
or ( n65824 , n65524 , n65823 );
and ( n65825 , n65521 , n65824 );
or ( n65826 , n65520 , n65825 );
and ( n65827 , n65517 , n65826 );
or ( n65828 , n65516 , n65827 );
and ( n65829 , n65513 , n65828 );
or ( n65830 , n65512 , n65829 );
and ( n65831 , n65509 , n65830 );
or ( n65832 , n65508 , n65831 );
and ( n65833 , n65505 , n65832 );
or ( n65834 , n65504 , n65833 );
and ( n65835 , n65501 , n65834 );
or ( n65836 , n65500 , n65835 );
and ( n65837 , n65497 , n65836 );
or ( n65838 , n65496 , n65837 );
and ( n65839 , n65493 , n65838 );
or ( n65840 , n65492 , n65839 );
and ( n65841 , n65489 , n65840 );
or ( n65842 , n65488 , n65841 );
and ( n65843 , n65485 , n65842 );
or ( n65844 , n65484 , n65843 );
and ( n65845 , n65481 , n65844 );
or ( n65846 , n65480 , n65845 );
and ( n65847 , n65477 , n65846 );
or ( n65848 , n65476 , n65847 );
and ( n65849 , n65473 , n65848 );
or ( n65850 , n65472 , n65849 );
and ( n65851 , n65469 , n65850 );
or ( n65852 , n65468 , n65851 );
and ( n65853 , n65465 , n65852 );
or ( n65854 , n65464 , n65853 );
and ( n65855 , n65461 , n65854 );
or ( n65856 , n65460 , n65855 );
and ( n65857 , n65457 , n65856 );
or ( n65858 , n65456 , n65857 );
and ( n65859 , n65453 , n65858 );
or ( n65860 , n65452 , n65859 );
and ( n65861 , n65449 , n65860 );
or ( n65862 , n65448 , n65861 );
and ( n65863 , n65445 , n65862 );
or ( n65864 , n65444 , n65863 );
and ( n65865 , n65441 , n65864 );
or ( n65866 , n65440 , n65865 );
and ( n65867 , n65437 , n65866 );
or ( n65868 , n65436 , n65867 );
and ( n65869 , n65433 , n65868 );
or ( n65870 , n65432 , n65869 );
and ( n65871 , n65429 , n65870 );
or ( n65872 , n65428 , n65871 );
and ( n65873 , n65425 , n65872 );
or ( n65874 , n65424 , n65873 );
and ( n65875 , n65421 , n65874 );
or ( n65876 , n65420 , n65875 );
and ( n65877 , n65417 , n65876 );
or ( n65878 , n65416 , n65877 );
and ( n65879 , n65413 , n65878 );
or ( n65880 , n65412 , n65879 );
and ( n65881 , n65409 , n65880 );
or ( n65882 , n65408 , n65881 );
and ( n65883 , n65405 , n65882 );
or ( n65884 , n65404 , n65883 );
and ( n65885 , n65401 , n65884 );
or ( n65886 , n65400 , n65885 );
and ( n65887 , n65397 , n65886 );
or ( n65888 , n65396 , n65887 );
and ( n65889 , n65393 , n65888 );
or ( n65890 , n65392 , n65889 );
and ( n65891 , n65389 , n65890 );
or ( n65892 , n65388 , n65891 );
and ( n65893 , n65385 , n65892 );
or ( n65894 , n65384 , n65893 );
and ( n65895 , n65381 , n65894 );
or ( n65896 , n65380 , n65895 );
and ( n65897 , n65377 , n65896 );
or ( n65898 , n65376 , n65897 );
xor ( n65899 , n65373 , n65898 );
and ( n65900 , n33403 , n5125 );
nor ( n65901 , n5126 , n65900 );
nor ( n65902 , n5477 , n32231 );
xor ( n65903 , n65901 , n65902 );
and ( n65904 , n64707 , n64708 );
and ( n65905 , n64709 , n64712 );
or ( n65906 , n65904 , n65905 );
xor ( n65907 , n65903 , n65906 );
nor ( n65908 , n5838 , n31083 );
xor ( n65909 , n65907 , n65908 );
and ( n65910 , n64713 , n64714 );
and ( n65911 , n64715 , n64718 );
or ( n65912 , n65910 , n65911 );
xor ( n65913 , n65909 , n65912 );
nor ( n65914 , n6212 , n29948 );
xor ( n65915 , n65913 , n65914 );
and ( n65916 , n64719 , n64720 );
and ( n65917 , n64721 , n64724 );
or ( n65918 , n65916 , n65917 );
xor ( n65919 , n65915 , n65918 );
nor ( n65920 , n6596 , n28833 );
xor ( n65921 , n65919 , n65920 );
and ( n65922 , n64725 , n64726 );
and ( n65923 , n64727 , n64730 );
or ( n65924 , n65922 , n65923 );
xor ( n65925 , n65921 , n65924 );
nor ( n65926 , n6997 , n27737 );
xor ( n65927 , n65925 , n65926 );
and ( n65928 , n64731 , n64732 );
and ( n65929 , n64733 , n64736 );
or ( n65930 , n65928 , n65929 );
xor ( n65931 , n65927 , n65930 );
nor ( n65932 , n7413 , n26660 );
xor ( n65933 , n65931 , n65932 );
and ( n65934 , n64737 , n64738 );
and ( n65935 , n64739 , n64742 );
or ( n65936 , n65934 , n65935 );
xor ( n65937 , n65933 , n65936 );
nor ( n65938 , n7841 , n25600 );
xor ( n65939 , n65937 , n65938 );
and ( n65940 , n64743 , n64744 );
and ( n65941 , n64745 , n64748 );
or ( n65942 , n65940 , n65941 );
xor ( n65943 , n65939 , n65942 );
nor ( n65944 , n8281 , n24564 );
xor ( n65945 , n65943 , n65944 );
and ( n65946 , n64749 , n64750 );
and ( n65947 , n64751 , n64754 );
or ( n65948 , n65946 , n65947 );
xor ( n65949 , n65945 , n65948 );
nor ( n65950 , n8737 , n23541 );
xor ( n65951 , n65949 , n65950 );
and ( n65952 , n64755 , n64756 );
and ( n65953 , n64757 , n64760 );
or ( n65954 , n65952 , n65953 );
xor ( n65955 , n65951 , n65954 );
nor ( n65956 , n9420 , n22541 );
xor ( n65957 , n65955 , n65956 );
and ( n65958 , n64761 , n64762 );
and ( n65959 , n64763 , n64766 );
or ( n65960 , n65958 , n65959 );
xor ( n65961 , n65957 , n65960 );
nor ( n65962 , n10312 , n21562 );
xor ( n65963 , n65961 , n65962 );
and ( n65964 , n64767 , n64768 );
and ( n65965 , n64769 , n64772 );
or ( n65966 , n65964 , n65965 );
xor ( n65967 , n65963 , n65966 );
nor ( n65968 , n11041 , n20601 );
xor ( n65969 , n65967 , n65968 );
and ( n65970 , n64773 , n64774 );
and ( n65971 , n64775 , n64778 );
or ( n65972 , n65970 , n65971 );
xor ( n65973 , n65969 , n65972 );
nor ( n65974 , n11790 , n19657 );
xor ( n65975 , n65973 , n65974 );
and ( n65976 , n64779 , n64780 );
and ( n65977 , n64781 , n64784 );
or ( n65978 , n65976 , n65977 );
xor ( n65979 , n65975 , n65978 );
nor ( n65980 , n12555 , n18734 );
xor ( n65981 , n65979 , n65980 );
and ( n65982 , n64785 , n64786 );
and ( n65983 , n64787 , n64790 );
or ( n65984 , n65982 , n65983 );
xor ( n65985 , n65981 , n65984 );
nor ( n65986 , n13340 , n17828 );
xor ( n65987 , n65985 , n65986 );
and ( n65988 , n64791 , n64792 );
and ( n65989 , n64793 , n64796 );
or ( n65990 , n65988 , n65989 );
xor ( n65991 , n65987 , n65990 );
nor ( n65992 , n14138 , n16943 );
xor ( n65993 , n65991 , n65992 );
and ( n65994 , n64797 , n64798 );
and ( n65995 , n64799 , n64802 );
or ( n65996 , n65994 , n65995 );
xor ( n65997 , n65993 , n65996 );
nor ( n65998 , n14959 , n16077 );
xor ( n65999 , n65997 , n65998 );
and ( n66000 , n64803 , n64804 );
and ( n66001 , n64805 , n64808 );
or ( n66002 , n66000 , n66001 );
xor ( n66003 , n65999 , n66002 );
nor ( n66004 , n15800 , n15230 );
xor ( n66005 , n66003 , n66004 );
and ( n66006 , n64809 , n64810 );
and ( n66007 , n64811 , n64814 );
or ( n66008 , n66006 , n66007 );
xor ( n66009 , n66005 , n66008 );
nor ( n66010 , n16660 , n14403 );
xor ( n66011 , n66009 , n66010 );
and ( n66012 , n64815 , n64816 );
and ( n66013 , n64817 , n64820 );
or ( n66014 , n66012 , n66013 );
xor ( n66015 , n66011 , n66014 );
nor ( n66016 , n17539 , n13599 );
xor ( n66017 , n66015 , n66016 );
and ( n66018 , n64821 , n64822 );
and ( n66019 , n64823 , n64826 );
or ( n66020 , n66018 , n66019 );
xor ( n66021 , n66017 , n66020 );
nor ( n66022 , n18439 , n12808 );
xor ( n66023 , n66021 , n66022 );
and ( n66024 , n64827 , n64828 );
and ( n66025 , n64829 , n64832 );
or ( n66026 , n66024 , n66025 );
xor ( n66027 , n66023 , n66026 );
nor ( n66028 , n19356 , n12037 );
xor ( n66029 , n66027 , n66028 );
and ( n66030 , n64833 , n64834 );
and ( n66031 , n64835 , n64838 );
or ( n66032 , n66030 , n66031 );
xor ( n66033 , n66029 , n66032 );
nor ( n66034 , n20294 , n11282 );
xor ( n66035 , n66033 , n66034 );
and ( n66036 , n64839 , n64840 );
and ( n66037 , n64841 , n64844 );
or ( n66038 , n66036 , n66037 );
xor ( n66039 , n66035 , n66038 );
nor ( n66040 , n21249 , n10547 );
xor ( n66041 , n66039 , n66040 );
and ( n66042 , n64845 , n64846 );
and ( n66043 , n64847 , n64850 );
or ( n66044 , n66042 , n66043 );
xor ( n66045 , n66041 , n66044 );
nor ( n66046 , n22222 , n9829 );
xor ( n66047 , n66045 , n66046 );
and ( n66048 , n64851 , n64852 );
and ( n66049 , n64853 , n64856 );
or ( n66050 , n66048 , n66049 );
xor ( n66051 , n66047 , n66050 );
nor ( n66052 , n23216 , n8955 );
xor ( n66053 , n66051 , n66052 );
and ( n66054 , n64857 , n64858 );
and ( n66055 , n64859 , n64862 );
or ( n66056 , n66054 , n66055 );
xor ( n66057 , n66053 , n66056 );
nor ( n66058 , n24233 , n603 );
xor ( n66059 , n66057 , n66058 );
and ( n66060 , n64863 , n64864 );
and ( n66061 , n64865 , n64868 );
or ( n66062 , n66060 , n66061 );
xor ( n66063 , n66059 , n66062 );
nor ( n66064 , n25263 , n652 );
xor ( n66065 , n66063 , n66064 );
and ( n66066 , n64869 , n64870 );
and ( n66067 , n64871 , n64874 );
or ( n66068 , n66066 , n66067 );
xor ( n66069 , n66065 , n66068 );
nor ( n66070 , n26317 , n624 );
xor ( n66071 , n66069 , n66070 );
and ( n66072 , n64875 , n64876 );
and ( n66073 , n64877 , n64880 );
or ( n66074 , n66072 , n66073 );
xor ( n66075 , n66071 , n66074 );
nor ( n66076 , n27388 , n648 );
xor ( n66077 , n66075 , n66076 );
and ( n66078 , n64881 , n64882 );
and ( n66079 , n64883 , n64886 );
or ( n66080 , n66078 , n66079 );
xor ( n66081 , n66077 , n66080 );
nor ( n66082 , n28478 , n686 );
xor ( n66083 , n66081 , n66082 );
and ( n66084 , n64887 , n64888 );
and ( n66085 , n64889 , n64892 );
or ( n66086 , n66084 , n66085 );
xor ( n66087 , n66083 , n66086 );
nor ( n66088 , n29587 , n735 );
xor ( n66089 , n66087 , n66088 );
and ( n66090 , n64893 , n64894 );
and ( n66091 , n64895 , n64898 );
or ( n66092 , n66090 , n66091 );
xor ( n66093 , n66089 , n66092 );
nor ( n66094 , n30716 , n798 );
xor ( n66095 , n66093 , n66094 );
and ( n66096 , n64899 , n64900 );
and ( n66097 , n64901 , n64904 );
or ( n66098 , n66096 , n66097 );
xor ( n66099 , n66095 , n66098 );
nor ( n66100 , n31858 , n870 );
xor ( n66101 , n66099 , n66100 );
and ( n66102 , n64905 , n64906 );
and ( n66103 , n64907 , n64910 );
or ( n66104 , n66102 , n66103 );
xor ( n66105 , n66101 , n66104 );
nor ( n66106 , n33024 , n960 );
xor ( n66107 , n66105 , n66106 );
and ( n66108 , n64911 , n64912 );
and ( n66109 , n64913 , n64916 );
or ( n66110 , n66108 , n66109 );
xor ( n66111 , n66107 , n66110 );
nor ( n66112 , n34215 , n1064 );
xor ( n66113 , n66111 , n66112 );
and ( n66114 , n64917 , n64918 );
and ( n66115 , n64919 , n64922 );
or ( n66116 , n66114 , n66115 );
xor ( n66117 , n66113 , n66116 );
nor ( n66118 , n35410 , n1178 );
xor ( n66119 , n66117 , n66118 );
and ( n66120 , n64923 , n64924 );
and ( n66121 , n64925 , n64928 );
or ( n66122 , n66120 , n66121 );
xor ( n66123 , n66119 , n66122 );
nor ( n66124 , n36611 , n1305 );
xor ( n66125 , n66123 , n66124 );
and ( n66126 , n64929 , n64930 );
and ( n66127 , n64931 , n64934 );
or ( n66128 , n66126 , n66127 );
xor ( n66129 , n66125 , n66128 );
nor ( n66130 , n37816 , n1447 );
xor ( n66131 , n66129 , n66130 );
and ( n66132 , n64935 , n64936 );
and ( n66133 , n64937 , n64940 );
or ( n66134 , n66132 , n66133 );
xor ( n66135 , n66131 , n66134 );
nor ( n66136 , n39018 , n1600 );
xor ( n66137 , n66135 , n66136 );
and ( n66138 , n64941 , n64942 );
and ( n66139 , n64943 , n64946 );
or ( n66140 , n66138 , n66139 );
xor ( n66141 , n66137 , n66140 );
nor ( n66142 , n40223 , n1768 );
xor ( n66143 , n66141 , n66142 );
and ( n66144 , n64947 , n64948 );
and ( n66145 , n64949 , n64952 );
or ( n66146 , n66144 , n66145 );
xor ( n66147 , n66143 , n66146 );
nor ( n66148 , n41428 , n1947 );
xor ( n66149 , n66147 , n66148 );
and ( n66150 , n64953 , n64954 );
and ( n66151 , n64955 , n64958 );
or ( n66152 , n66150 , n66151 );
xor ( n66153 , n66149 , n66152 );
nor ( n66154 , n42632 , n2139 );
xor ( n66155 , n66153 , n66154 );
and ( n66156 , n64959 , n64960 );
and ( n66157 , n64961 , n64964 );
or ( n66158 , n66156 , n66157 );
xor ( n66159 , n66155 , n66158 );
nor ( n66160 , n43834 , n2345 );
xor ( n66161 , n66159 , n66160 );
and ( n66162 , n64965 , n64966 );
and ( n66163 , n64967 , n64970 );
or ( n66164 , n66162 , n66163 );
xor ( n66165 , n66161 , n66164 );
nor ( n66166 , n45038 , n2568 );
xor ( n66167 , n66165 , n66166 );
and ( n66168 , n64971 , n64972 );
and ( n66169 , n64973 , n64976 );
or ( n66170 , n66168 , n66169 );
xor ( n66171 , n66167 , n66170 );
nor ( n66172 , n46239 , n2799 );
xor ( n66173 , n66171 , n66172 );
and ( n66174 , n64977 , n64978 );
and ( n66175 , n64979 , n64982 );
or ( n66176 , n66174 , n66175 );
xor ( n66177 , n66173 , n66176 );
nor ( n66178 , n47440 , n3045 );
xor ( n66179 , n66177 , n66178 );
and ( n66180 , n64983 , n64984 );
and ( n66181 , n64985 , n64988 );
or ( n66182 , n66180 , n66181 );
xor ( n66183 , n66179 , n66182 );
nor ( n66184 , n48641 , n3302 );
xor ( n66185 , n66183 , n66184 );
and ( n66186 , n64989 , n64990 );
and ( n66187 , n64991 , n64994 );
or ( n66188 , n66186 , n66187 );
xor ( n66189 , n66185 , n66188 );
nor ( n66190 , n49841 , n3572 );
xor ( n66191 , n66189 , n66190 );
and ( n66192 , n64995 , n64996 );
and ( n66193 , n64997 , n65000 );
or ( n66194 , n66192 , n66193 );
xor ( n66195 , n66191 , n66194 );
nor ( n66196 , n51040 , n3855 );
xor ( n66197 , n66195 , n66196 );
and ( n66198 , n65001 , n65002 );
and ( n66199 , n65003 , n65006 );
or ( n66200 , n66198 , n66199 );
xor ( n66201 , n66197 , n66200 );
nor ( n66202 , n52238 , n4153 );
xor ( n66203 , n66201 , n66202 );
and ( n66204 , n65007 , n65008 );
and ( n66205 , n65009 , n65012 );
or ( n66206 , n66204 , n66205 );
xor ( n66207 , n66203 , n66206 );
nor ( n66208 , n53432 , n4460 );
xor ( n66209 , n66207 , n66208 );
and ( n66210 , n65013 , n65014 );
and ( n66211 , n65015 , n65018 );
or ( n66212 , n66210 , n66211 );
xor ( n66213 , n66209 , n66212 );
nor ( n66214 , n54629 , n4788 );
xor ( n66215 , n66213 , n66214 );
and ( n66216 , n65019 , n65020 );
and ( n66217 , n65021 , n65024 );
or ( n66218 , n66216 , n66217 );
xor ( n66219 , n66215 , n66218 );
nor ( n66220 , n55826 , n5128 );
xor ( n66221 , n66219 , n66220 );
and ( n66222 , n65025 , n65026 );
and ( n66223 , n65027 , n65030 );
or ( n66224 , n66222 , n66223 );
xor ( n66225 , n66221 , n66224 );
nor ( n66226 , n57022 , n5479 );
xor ( n66227 , n66225 , n66226 );
and ( n66228 , n65031 , n65032 );
and ( n66229 , n65033 , n65036 );
or ( n66230 , n66228 , n66229 );
xor ( n66231 , n66227 , n66230 );
nor ( n66232 , n58217 , n5840 );
xor ( n66233 , n66231 , n66232 );
and ( n66234 , n65037 , n65038 );
and ( n66235 , n65039 , n65042 );
or ( n66236 , n66234 , n66235 );
xor ( n66237 , n66233 , n66236 );
nor ( n66238 , n59412 , n6214 );
xor ( n66239 , n66237 , n66238 );
and ( n66240 , n65043 , n65044 );
and ( n66241 , n65045 , n65048 );
or ( n66242 , n66240 , n66241 );
xor ( n66243 , n66239 , n66242 );
nor ( n66244 , n60600 , n6598 );
xor ( n66245 , n66243 , n66244 );
and ( n66246 , n65049 , n65050 );
and ( n66247 , n65051 , n65054 );
or ( n66248 , n66246 , n66247 );
xor ( n66249 , n66245 , n66248 );
nor ( n66250 , n61791 , n6999 );
xor ( n66251 , n66249 , n66250 );
and ( n66252 , n65055 , n65056 );
and ( n66253 , n65057 , n65060 );
or ( n66254 , n66252 , n66253 );
xor ( n66255 , n66251 , n66254 );
nor ( n66256 , n62982 , n7415 );
xor ( n66257 , n66255 , n66256 );
and ( n66258 , n65061 , n65062 );
and ( n66259 , n65063 , n65066 );
or ( n66260 , n66258 , n66259 );
xor ( n66261 , n66257 , n66260 );
nor ( n66262 , n64172 , n7843 );
xor ( n66263 , n66261 , n66262 );
and ( n66264 , n65067 , n65068 );
and ( n66265 , n65069 , n65072 );
or ( n66266 , n66264 , n66265 );
xor ( n66267 , n66263 , n66266 );
nor ( n66268 , n65360 , n8283 );
xor ( n66269 , n66267 , n66268 );
and ( n66270 , n65073 , n65074 );
and ( n66271 , n65075 , n65078 );
or ( n66272 , n66270 , n66271 );
xor ( n66273 , n66269 , n66272 );
and ( n66274 , n65091 , n65095 );
and ( n66275 , n65095 , n65346 );
and ( n66276 , n65091 , n65346 );
or ( n66277 , n66274 , n66275 , n66276 );
and ( n66278 , n33774 , n5103 );
not ( n66279 , n5103 );
nor ( n66280 , n66278 , n66279 );
xor ( n66281 , n66277 , n66280 );
and ( n66282 , n65101 , n65105 );
and ( n66283 , n65105 , n65173 );
and ( n66284 , n65101 , n65173 );
or ( n66285 , n66282 , n66283 , n66284 );
and ( n66286 , n65097 , n65174 );
and ( n66287 , n65174 , n65345 );
and ( n66288 , n65097 , n65345 );
or ( n66289 , n66286 , n66287 , n66288 );
xor ( n66290 , n66285 , n66289 );
and ( n66291 , n65292 , n65344 );
and ( n66292 , n65179 , n65180 );
and ( n66293 , n65180 , n65291 );
and ( n66294 , n65179 , n65291 );
or ( n66295 , n66292 , n66293 , n66294 );
and ( n66296 , n65110 , n65114 );
and ( n66297 , n65114 , n65172 );
and ( n66298 , n65110 , n65172 );
or ( n66299 , n66296 , n66297 , n66298 );
xor ( n66300 , n66295 , n66299 );
and ( n66301 , n65141 , n65145 );
and ( n66302 , n65145 , n65151 );
and ( n66303 , n65141 , n65151 );
or ( n66304 , n66301 , n66302 , n66303 );
and ( n66305 , n65119 , n65123 );
and ( n66306 , n65123 , n65171 );
and ( n66307 , n65119 , n65171 );
or ( n66308 , n66305 , n66306 , n66307 );
xor ( n66309 , n66304 , n66308 );
and ( n66310 , n65128 , n65132 );
and ( n66311 , n65132 , n65170 );
and ( n66312 , n65128 , n65170 );
or ( n66313 , n66310 , n66311 , n66312 );
and ( n66314 , n65189 , n65214 );
and ( n66315 , n65214 , n65252 );
and ( n66316 , n65189 , n65252 );
or ( n66317 , n66314 , n66315 , n66316 );
xor ( n66318 , n66313 , n66317 );
and ( n66319 , n65137 , n65152 );
and ( n66320 , n65152 , n65169 );
and ( n66321 , n65137 , n65169 );
or ( n66322 , n66319 , n66320 , n66321 );
and ( n66323 , n65193 , n65197 );
and ( n66324 , n65197 , n65213 );
and ( n66325 , n65193 , n65213 );
or ( n66326 , n66323 , n66324 , n66325 );
xor ( n66327 , n66322 , n66326 );
and ( n66328 , n65157 , n65162 );
and ( n66329 , n65162 , n65168 );
and ( n66330 , n65157 , n65168 );
or ( n66331 , n66328 , n66329 , n66330 );
and ( n66332 , n65147 , n65148 );
and ( n66333 , n65148 , n65150 );
and ( n66334 , n65147 , n65150 );
or ( n66335 , n66332 , n66333 , n66334 );
and ( n66336 , n65158 , n65159 );
and ( n66337 , n65159 , n65161 );
and ( n66338 , n65158 , n65161 );
or ( n66339 , n66336 , n66337 , n66338 );
xor ( n66340 , n66335 , n66339 );
and ( n66341 , n30695 , n6132 );
and ( n66342 , n31836 , n5765 );
xor ( n66343 , n66341 , n66342 );
and ( n66344 , n32649 , n5408 );
xor ( n66345 , n66343 , n66344 );
xor ( n66346 , n66340 , n66345 );
xor ( n66347 , n66331 , n66346 );
and ( n66348 , n65164 , n65165 );
and ( n66349 , n65165 , n65167 );
and ( n66350 , n65164 , n65167 );
or ( n66351 , n66348 , n66349 , n66350 );
and ( n66352 , n27361 , n7310 );
and ( n66353 , n28456 , n6971 );
xor ( n66354 , n66352 , n66353 );
and ( n66355 , n29559 , n6504 );
xor ( n66356 , n66354 , n66355 );
xor ( n66357 , n66351 , n66356 );
and ( n66358 , n24214 , n8669 );
and ( n66359 , n25243 , n8243 );
xor ( n66360 , n66358 , n66359 );
and ( n66361 , n26296 , n7662 );
xor ( n66362 , n66360 , n66361 );
xor ( n66363 , n66357 , n66362 );
xor ( n66364 , n66347 , n66363 );
xor ( n66365 , n66327 , n66364 );
xor ( n66366 , n66318 , n66365 );
xor ( n66367 , n66309 , n66366 );
xor ( n66368 , n66300 , n66367 );
xor ( n66369 , n66291 , n66368 );
and ( n66370 , n65185 , n65253 );
and ( n66371 , n65253 , n65290 );
and ( n66372 , n65185 , n65290 );
or ( n66373 , n66370 , n66371 , n66372 );
and ( n66374 , n65296 , n65343 );
xor ( n66375 , n66373 , n66374 );
and ( n66376 , n65258 , n65262 );
and ( n66377 , n65262 , n65289 );
and ( n66378 , n65258 , n65289 );
or ( n66379 , n66376 , n66377 , n66378 );
and ( n66380 , n65219 , n65235 );
and ( n66381 , n65235 , n65251 );
and ( n66382 , n65219 , n65251 );
or ( n66383 , n66380 , n66381 , n66382 );
and ( n66384 , n65202 , n65206 );
and ( n66385 , n65206 , n65212 );
and ( n66386 , n65202 , n65212 );
or ( n66387 , n66384 , n66385 , n66386 );
and ( n66388 , n65223 , n65228 );
and ( n66389 , n65228 , n65234 );
and ( n66390 , n65223 , n65234 );
or ( n66391 , n66388 , n66389 , n66390 );
xor ( n66392 , n66387 , n66391 );
and ( n66393 , n65208 , n65209 );
and ( n66394 , n65209 , n65211 );
and ( n66395 , n65208 , n65211 );
or ( n66396 , n66393 , n66394 , n66395 );
and ( n66397 , n65224 , n65225 );
and ( n66398 , n65225 , n65227 );
and ( n66399 , n65224 , n65227 );
or ( n66400 , n66397 , n66398 , n66399 );
xor ( n66401 , n66396 , n66400 );
and ( n66402 , n21216 , n10977 );
and ( n66403 , n22186 , n10239 );
xor ( n66404 , n66402 , n66403 );
and ( n66405 , n22892 , n9348 );
xor ( n66406 , n66404 , n66405 );
xor ( n66407 , n66401 , n66406 );
xor ( n66408 , n66392 , n66407 );
xor ( n66409 , n66383 , n66408 );
and ( n66410 , n65240 , n65244 );
and ( n66411 , n65244 , n65250 );
and ( n66412 , n65240 , n65250 );
or ( n66413 , n66410 , n66411 , n66412 );
and ( n66414 , n65230 , n65231 );
and ( n66415 , n65231 , n65233 );
and ( n66416 , n65230 , n65233 );
or ( n66417 , n66414 , n66415 , n66416 );
and ( n66418 , n18144 , n13256 );
and ( n66419 , n19324 , n12531 );
xor ( n66420 , n66418 , n66419 );
and ( n66421 , n20233 , n11718 );
xor ( n66422 , n66420 , n66421 );
xor ( n66423 , n66417 , n66422 );
buf ( n66424 , n15758 );
and ( n66425 , n16637 , n14838 );
xor ( n66426 , n66424 , n66425 );
and ( n66427 , n17512 , n14044 );
xor ( n66428 , n66426 , n66427 );
xor ( n66429 , n66423 , n66428 );
xor ( n66430 , n66413 , n66429 );
and ( n66431 , n65246 , n65247 );
and ( n66432 , n65247 , n65249 );
and ( n66433 , n65246 , n65249 );
or ( n66434 , n66431 , n66432 , n66433 );
and ( n66435 , n65277 , n65278 );
and ( n66436 , n65278 , n65280 );
and ( n66437 , n65277 , n65280 );
or ( n66438 , n66435 , n66436 , n66437 );
xor ( n66439 , n66434 , n66438 );
and ( n66440 , n13322 , n18407 );
and ( n66441 , n14118 , n17422 );
xor ( n66442 , n66440 , n66441 );
and ( n66443 , n14938 , n16550 );
xor ( n66444 , n66442 , n66443 );
xor ( n66445 , n66439 , n66444 );
xor ( n66446 , n66430 , n66445 );
xor ( n66447 , n66409 , n66446 );
xor ( n66448 , n66379 , n66447 );
and ( n66449 , n65267 , n65271 );
and ( n66450 , n65271 , n65288 );
and ( n66451 , n65267 , n65288 );
or ( n66452 , n66449 , n66450 , n66451 );
and ( n66453 , n65301 , n65316 );
and ( n66454 , n65316 , n65333 );
and ( n66455 , n65301 , n65333 );
or ( n66456 , n66453 , n66454 , n66455 );
xor ( n66457 , n66452 , n66456 );
and ( n66458 , n65276 , n65281 );
and ( n66459 , n65281 , n65287 );
and ( n66460 , n65276 , n65287 );
or ( n66461 , n66458 , n66459 , n66460 );
and ( n66462 , n65305 , n65309 );
and ( n66463 , n65309 , n65315 );
and ( n66464 , n65305 , n65315 );
or ( n66465 , n66462 , n66463 , n66464 );
xor ( n66466 , n66461 , n66465 );
and ( n66467 , n65283 , n65284 );
and ( n66468 , n65284 , n65286 );
and ( n66469 , n65283 , n65286 );
or ( n66470 , n66467 , n66468 , n66469 );
and ( n66471 , n11015 , n20976 );
and ( n66472 , n11769 , n20156 );
xor ( n66473 , n66471 , n66472 );
and ( n66474 , n12320 , n19222 );
xor ( n66475 , n66473 , n66474 );
xor ( n66476 , n66470 , n66475 );
and ( n66477 , n8718 , n24137 );
and ( n66478 , n9400 , n23075 );
xor ( n66479 , n66477 , n66478 );
and ( n66480 , n10291 , n22065 );
xor ( n66481 , n66479 , n66480 );
xor ( n66482 , n66476 , n66481 );
xor ( n66483 , n66466 , n66482 );
xor ( n66484 , n66457 , n66483 );
xor ( n66485 , n66448 , n66484 );
xor ( n66486 , n66375 , n66485 );
and ( n66487 , n65297 , n65334 );
and ( n66488 , n65334 , n65342 );
and ( n66489 , n65297 , n65342 );
or ( n66490 , n66487 , n66488 , n66489 );
and ( n66491 , n65337 , n65340 );
and ( n66492 , n65336 , n65341 );
xor ( n66493 , n66491 , n66492 );
and ( n66494 , n65321 , n65326 );
and ( n66495 , n65326 , n65332 );
and ( n66496 , n65321 , n65332 );
or ( n66497 , n66494 , n66495 , n66496 );
and ( n66498 , n65311 , n65312 );
and ( n66499 , n65312 , n65314 );
and ( n66500 , n65311 , n65314 );
or ( n66501 , n66498 , n66499 , n66500 );
and ( n66502 , n65322 , n65323 );
and ( n66503 , n65323 , n65325 );
and ( n66504 , n65322 , n65325 );
or ( n66505 , n66502 , n66503 , n66504 );
xor ( n66506 , n66501 , n66505 );
and ( n66507 , n7385 , n27296 );
and ( n66508 , n7808 , n26216 );
xor ( n66509 , n66507 , n66508 );
and ( n66510 , n8079 , n25163 );
xor ( n66511 , n66509 , n66510 );
xor ( n66512 , n66506 , n66511 );
xor ( n66513 , n66497 , n66512 );
and ( n66514 , n65328 , n65329 );
and ( n66515 , n65329 , n65331 );
and ( n66516 , n65328 , n65331 );
or ( n66517 , n66514 , n66515 , n66516 );
and ( n66518 , n6187 , n30629 );
and ( n66519 , n6569 , n29508 );
xor ( n66520 , n66518 , n66519 );
and ( n66521 , n6816 , n28406 );
xor ( n66522 , n66520 , n66521 );
xor ( n66523 , n66517 , n66522 );
not ( n66524 , n4959 );
and ( n66525 , n34193 , n4959 );
nor ( n66526 , n66524 , n66525 );
and ( n66527 , n5459 , n32999 );
xor ( n66528 , n66526 , n66527 );
and ( n66529 , n5819 , n31761 );
xor ( n66530 , n66528 , n66529 );
xor ( n66531 , n66523 , n66530 );
xor ( n66532 , n66513 , n66531 );
xor ( n66533 , n66493 , n66532 );
xor ( n66534 , n66490 , n66533 );
xor ( n66535 , n66486 , n66534 );
xor ( n66536 , n66369 , n66535 );
xor ( n66537 , n66290 , n66536 );
xor ( n66538 , n66281 , n66537 );
and ( n66539 , n65083 , n65086 );
and ( n66540 , n65086 , n65347 );
and ( n66541 , n65083 , n65347 );
or ( n66542 , n66539 , n66540 , n66541 );
xor ( n66543 , n66538 , n66542 );
and ( n66544 , n65348 , n65352 );
and ( n66545 , n65353 , n65356 );
or ( n66546 , n66544 , n66545 );
xor ( n66547 , n66543 , n66546 );
buf ( n66548 , n66547 );
buf ( n66549 , n66548 );
not ( n66550 , n66549 );
nor ( n66551 , n66550 , n8739 );
xor ( n66552 , n66273 , n66551 );
and ( n66553 , n65079 , n65361 );
and ( n66554 , n65362 , n65365 );
or ( n66555 , n66553 , n66554 );
xor ( n66556 , n66552 , n66555 );
buf ( n66557 , n66556 );
buf ( n66558 , n66557 );
not ( n66559 , n66558 );
buf ( n66560 , n589 );
not ( n66561 , n66560 );
nor ( n66562 , n66559 , n66561 );
xor ( n66563 , n65899 , n66562 );
xor ( n66564 , n65377 , n65896 );
nor ( n66565 , n65369 , n66561 );
and ( n66566 , n66564 , n66565 );
xor ( n66567 , n66564 , n66565 );
xor ( n66568 , n65381 , n65894 );
nor ( n66569 , n64181 , n66561 );
and ( n66570 , n66568 , n66569 );
xor ( n66571 , n66568 , n66569 );
xor ( n66572 , n65385 , n65892 );
nor ( n66573 , n62991 , n66561 );
and ( n66574 , n66572 , n66573 );
xor ( n66575 , n66572 , n66573 );
xor ( n66576 , n65389 , n65890 );
nor ( n66577 , n61800 , n66561 );
and ( n66578 , n66576 , n66577 );
xor ( n66579 , n66576 , n66577 );
xor ( n66580 , n65393 , n65888 );
nor ( n66581 , n60609 , n66561 );
and ( n66582 , n66580 , n66581 );
xor ( n66583 , n66580 , n66581 );
xor ( n66584 , n65397 , n65886 );
nor ( n66585 , n59421 , n66561 );
and ( n66586 , n66584 , n66585 );
xor ( n66587 , n66584 , n66585 );
xor ( n66588 , n65401 , n65884 );
nor ( n66589 , n58226 , n66561 );
and ( n66590 , n66588 , n66589 );
xor ( n66591 , n66588 , n66589 );
xor ( n66592 , n65405 , n65882 );
nor ( n66593 , n57031 , n66561 );
and ( n66594 , n66592 , n66593 );
xor ( n66595 , n66592 , n66593 );
xor ( n66596 , n65409 , n65880 );
nor ( n66597 , n55835 , n66561 );
and ( n66598 , n66596 , n66597 );
xor ( n66599 , n66596 , n66597 );
xor ( n66600 , n65413 , n65878 );
nor ( n66601 , n54638 , n66561 );
and ( n66602 , n66600 , n66601 );
xor ( n66603 , n66600 , n66601 );
xor ( n66604 , n65417 , n65876 );
nor ( n66605 , n53441 , n66561 );
and ( n66606 , n66604 , n66605 );
xor ( n66607 , n66604 , n66605 );
xor ( n66608 , n65421 , n65874 );
nor ( n66609 , n52247 , n66561 );
and ( n66610 , n66608 , n66609 );
xor ( n66611 , n66608 , n66609 );
xor ( n66612 , n65425 , n65872 );
nor ( n66613 , n51049 , n66561 );
and ( n66614 , n66612 , n66613 );
xor ( n66615 , n66612 , n66613 );
xor ( n66616 , n65429 , n65870 );
nor ( n66617 , n49850 , n66561 );
and ( n66618 , n66616 , n66617 );
xor ( n66619 , n66616 , n66617 );
xor ( n66620 , n65433 , n65868 );
nor ( n66621 , n48650 , n66561 );
and ( n66622 , n66620 , n66621 );
xor ( n66623 , n66620 , n66621 );
xor ( n66624 , n65437 , n65866 );
nor ( n66625 , n47449 , n66561 );
and ( n66626 , n66624 , n66625 );
xor ( n66627 , n66624 , n66625 );
xor ( n66628 , n65441 , n65864 );
nor ( n66629 , n46248 , n66561 );
and ( n66630 , n66628 , n66629 );
xor ( n66631 , n66628 , n66629 );
xor ( n66632 , n65445 , n65862 );
nor ( n66633 , n45047 , n66561 );
and ( n66634 , n66632 , n66633 );
xor ( n66635 , n66632 , n66633 );
xor ( n66636 , n65449 , n65860 );
nor ( n66637 , n43843 , n66561 );
and ( n66638 , n66636 , n66637 );
xor ( n66639 , n66636 , n66637 );
xor ( n66640 , n65453 , n65858 );
nor ( n66641 , n42641 , n66561 );
and ( n66642 , n66640 , n66641 );
xor ( n66643 , n66640 , n66641 );
xor ( n66644 , n65457 , n65856 );
nor ( n66645 , n41437 , n66561 );
and ( n66646 , n66644 , n66645 );
xor ( n66647 , n66644 , n66645 );
xor ( n66648 , n65461 , n65854 );
nor ( n66649 , n40232 , n66561 );
and ( n66650 , n66648 , n66649 );
xor ( n66651 , n66648 , n66649 );
xor ( n66652 , n65465 , n65852 );
nor ( n66653 , n39027 , n66561 );
and ( n66654 , n66652 , n66653 );
xor ( n66655 , n66652 , n66653 );
xor ( n66656 , n65469 , n65850 );
nor ( n66657 , n37825 , n66561 );
and ( n66658 , n66656 , n66657 );
xor ( n66659 , n66656 , n66657 );
xor ( n66660 , n65473 , n65848 );
nor ( n66661 , n36620 , n66561 );
and ( n66662 , n66660 , n66661 );
xor ( n66663 , n66660 , n66661 );
xor ( n66664 , n65477 , n65846 );
nor ( n66665 , n35419 , n66561 );
and ( n66666 , n66664 , n66665 );
xor ( n66667 , n66664 , n66665 );
xor ( n66668 , n65481 , n65844 );
nor ( n66669 , n34224 , n66561 );
and ( n66670 , n66668 , n66669 );
xor ( n66671 , n66668 , n66669 );
xor ( n66672 , n65485 , n65842 );
nor ( n66673 , n33033 , n66561 );
and ( n66674 , n66672 , n66673 );
xor ( n66675 , n66672 , n66673 );
xor ( n66676 , n65489 , n65840 );
nor ( n66677 , n31867 , n66561 );
and ( n66678 , n66676 , n66677 );
xor ( n66679 , n66676 , n66677 );
xor ( n66680 , n65493 , n65838 );
nor ( n66681 , n30725 , n66561 );
and ( n66682 , n66680 , n66681 );
xor ( n66683 , n66680 , n66681 );
xor ( n66684 , n65497 , n65836 );
nor ( n66685 , n29596 , n66561 );
and ( n66686 , n66684 , n66685 );
xor ( n66687 , n66684 , n66685 );
xor ( n66688 , n65501 , n65834 );
nor ( n66689 , n28487 , n66561 );
and ( n66690 , n66688 , n66689 );
xor ( n66691 , n66688 , n66689 );
xor ( n66692 , n65505 , n65832 );
nor ( n66693 , n27397 , n66561 );
and ( n66694 , n66692 , n66693 );
xor ( n66695 , n66692 , n66693 );
xor ( n66696 , n65509 , n65830 );
nor ( n66697 , n26326 , n66561 );
and ( n66698 , n66696 , n66697 );
xor ( n66699 , n66696 , n66697 );
xor ( n66700 , n65513 , n65828 );
nor ( n66701 , n25272 , n66561 );
and ( n66702 , n66700 , n66701 );
xor ( n66703 , n66700 , n66701 );
xor ( n66704 , n65517 , n65826 );
nor ( n66705 , n24242 , n66561 );
and ( n66706 , n66704 , n66705 );
xor ( n66707 , n66704 , n66705 );
xor ( n66708 , n65521 , n65824 );
nor ( n66709 , n23225 , n66561 );
and ( n66710 , n66708 , n66709 );
xor ( n66711 , n66708 , n66709 );
xor ( n66712 , n65525 , n65822 );
nor ( n66713 , n22231 , n66561 );
and ( n66714 , n66712 , n66713 );
xor ( n66715 , n66712 , n66713 );
xor ( n66716 , n65529 , n65820 );
nor ( n66717 , n21258 , n66561 );
and ( n66718 , n66716 , n66717 );
xor ( n66719 , n66716 , n66717 );
xor ( n66720 , n65533 , n65818 );
nor ( n66721 , n20303 , n66561 );
and ( n66722 , n66720 , n66721 );
xor ( n66723 , n66720 , n66721 );
xor ( n66724 , n65537 , n65816 );
nor ( n66725 , n19365 , n66561 );
and ( n66726 , n66724 , n66725 );
xor ( n66727 , n66724 , n66725 );
xor ( n66728 , n65541 , n65814 );
nor ( n66729 , n18448 , n66561 );
and ( n66730 , n66728 , n66729 );
xor ( n66731 , n66728 , n66729 );
xor ( n66732 , n65545 , n65812 );
nor ( n66733 , n17548 , n66561 );
and ( n66734 , n66732 , n66733 );
xor ( n66735 , n66732 , n66733 );
xor ( n66736 , n65549 , n65810 );
nor ( n66737 , n16669 , n66561 );
and ( n66738 , n66736 , n66737 );
xor ( n66739 , n66736 , n66737 );
xor ( n66740 , n65553 , n65808 );
nor ( n66741 , n15809 , n66561 );
and ( n66742 , n66740 , n66741 );
xor ( n66743 , n66740 , n66741 );
xor ( n66744 , n65557 , n65806 );
nor ( n66745 , n14968 , n66561 );
and ( n66746 , n66744 , n66745 );
xor ( n66747 , n66744 , n66745 );
xor ( n66748 , n65561 , n65804 );
nor ( n66749 , n14147 , n66561 );
and ( n66750 , n66748 , n66749 );
xor ( n66751 , n66748 , n66749 );
xor ( n66752 , n65565 , n65802 );
nor ( n66753 , n13349 , n66561 );
and ( n66754 , n66752 , n66753 );
xor ( n66755 , n66752 , n66753 );
xor ( n66756 , n65569 , n65800 );
nor ( n66757 , n12564 , n66561 );
and ( n66758 , n66756 , n66757 );
xor ( n66759 , n66756 , n66757 );
xor ( n66760 , n65573 , n65798 );
nor ( n66761 , n11799 , n66561 );
and ( n66762 , n66760 , n66761 );
xor ( n66763 , n66760 , n66761 );
xor ( n66764 , n65577 , n65796 );
nor ( n66765 , n11050 , n66561 );
and ( n66766 , n66764 , n66765 );
xor ( n66767 , n66764 , n66765 );
xor ( n66768 , n65581 , n65794 );
nor ( n66769 , n10321 , n66561 );
and ( n66770 , n66768 , n66769 );
xor ( n66771 , n66768 , n66769 );
xor ( n66772 , n65585 , n65792 );
nor ( n66773 , n9429 , n66561 );
and ( n66774 , n66772 , n66773 );
xor ( n66775 , n66772 , n66773 );
xor ( n66776 , n65589 , n65790 );
nor ( n66777 , n8949 , n66561 );
and ( n66778 , n66776 , n66777 );
xor ( n66779 , n66776 , n66777 );
xor ( n66780 , n65593 , n65788 );
nor ( n66781 , n9437 , n66561 );
and ( n66782 , n66780 , n66781 );
xor ( n66783 , n66780 , n66781 );
xor ( n66784 , n65597 , n65786 );
nor ( n66785 , n9446 , n66561 );
and ( n66786 , n66784 , n66785 );
xor ( n66787 , n66784 , n66785 );
xor ( n66788 , n65601 , n65784 );
nor ( n66789 , n9455 , n66561 );
and ( n66790 , n66788 , n66789 );
xor ( n66791 , n66788 , n66789 );
xor ( n66792 , n65605 , n65782 );
nor ( n66793 , n9464 , n66561 );
and ( n66794 , n66792 , n66793 );
xor ( n66795 , n66792 , n66793 );
xor ( n66796 , n65609 , n65780 );
nor ( n66797 , n9473 , n66561 );
and ( n66798 , n66796 , n66797 );
xor ( n66799 , n66796 , n66797 );
xor ( n66800 , n65613 , n65778 );
nor ( n66801 , n9482 , n66561 );
and ( n66802 , n66800 , n66801 );
xor ( n66803 , n66800 , n66801 );
xor ( n66804 , n65617 , n65776 );
nor ( n66805 , n9491 , n66561 );
and ( n66806 , n66804 , n66805 );
xor ( n66807 , n66804 , n66805 );
xor ( n66808 , n65621 , n65774 );
nor ( n66809 , n9500 , n66561 );
and ( n66810 , n66808 , n66809 );
xor ( n66811 , n66808 , n66809 );
xor ( n66812 , n65625 , n65772 );
nor ( n66813 , n9509 , n66561 );
and ( n66814 , n66812 , n66813 );
xor ( n66815 , n66812 , n66813 );
xor ( n66816 , n65629 , n65770 );
nor ( n66817 , n9518 , n66561 );
and ( n66818 , n66816 , n66817 );
xor ( n66819 , n66816 , n66817 );
xor ( n66820 , n65633 , n65768 );
nor ( n66821 , n9527 , n66561 );
and ( n66822 , n66820 , n66821 );
xor ( n66823 , n66820 , n66821 );
xor ( n66824 , n65637 , n65766 );
nor ( n66825 , n9536 , n66561 );
and ( n66826 , n66824 , n66825 );
xor ( n66827 , n66824 , n66825 );
xor ( n66828 , n65641 , n65764 );
nor ( n66829 , n9545 , n66561 );
and ( n66830 , n66828 , n66829 );
xor ( n66831 , n66828 , n66829 );
xor ( n66832 , n65645 , n65762 );
nor ( n66833 , n9554 , n66561 );
and ( n66834 , n66832 , n66833 );
xor ( n66835 , n66832 , n66833 );
xor ( n66836 , n65649 , n65760 );
nor ( n66837 , n9563 , n66561 );
and ( n66838 , n66836 , n66837 );
xor ( n66839 , n66836 , n66837 );
xor ( n66840 , n65653 , n65758 );
nor ( n66841 , n9572 , n66561 );
and ( n66842 , n66840 , n66841 );
xor ( n66843 , n66840 , n66841 );
xor ( n66844 , n65657 , n65756 );
nor ( n66845 , n9581 , n66561 );
and ( n66846 , n66844 , n66845 );
xor ( n66847 , n66844 , n66845 );
xor ( n66848 , n65661 , n65754 );
nor ( n66849 , n9590 , n66561 );
and ( n66850 , n66848 , n66849 );
xor ( n66851 , n66848 , n66849 );
xor ( n66852 , n65665 , n65752 );
nor ( n66853 , n9599 , n66561 );
and ( n66854 , n66852 , n66853 );
xor ( n66855 , n66852 , n66853 );
xor ( n66856 , n65669 , n65750 );
nor ( n66857 , n9608 , n66561 );
and ( n66858 , n66856 , n66857 );
xor ( n66859 , n66856 , n66857 );
xor ( n66860 , n65673 , n65748 );
nor ( n66861 , n9617 , n66561 );
and ( n66862 , n66860 , n66861 );
xor ( n66863 , n66860 , n66861 );
xor ( n66864 , n65677 , n65746 );
nor ( n66865 , n9626 , n66561 );
and ( n66866 , n66864 , n66865 );
xor ( n66867 , n66864 , n66865 );
xor ( n66868 , n65681 , n65744 );
nor ( n66869 , n9635 , n66561 );
and ( n66870 , n66868 , n66869 );
xor ( n66871 , n66868 , n66869 );
xor ( n66872 , n65685 , n65742 );
nor ( n66873 , n9644 , n66561 );
and ( n66874 , n66872 , n66873 );
xor ( n66875 , n66872 , n66873 );
xor ( n66876 , n65689 , n65740 );
nor ( n66877 , n9653 , n66561 );
and ( n66878 , n66876 , n66877 );
xor ( n66879 , n66876 , n66877 );
xor ( n66880 , n65693 , n65738 );
nor ( n66881 , n9662 , n66561 );
and ( n66882 , n66880 , n66881 );
xor ( n66883 , n66880 , n66881 );
xor ( n66884 , n65697 , n65736 );
nor ( n66885 , n9671 , n66561 );
and ( n66886 , n66884 , n66885 );
xor ( n66887 , n66884 , n66885 );
xor ( n66888 , n65701 , n65734 );
nor ( n66889 , n9680 , n66561 );
and ( n66890 , n66888 , n66889 );
xor ( n66891 , n66888 , n66889 );
xor ( n66892 , n65705 , n65732 );
nor ( n66893 , n9689 , n66561 );
and ( n66894 , n66892 , n66893 );
xor ( n66895 , n66892 , n66893 );
xor ( n66896 , n65709 , n65730 );
nor ( n66897 , n9698 , n66561 );
and ( n66898 , n66896 , n66897 );
xor ( n66899 , n66896 , n66897 );
xor ( n66900 , n65713 , n65728 );
nor ( n66901 , n9707 , n66561 );
and ( n66902 , n66900 , n66901 );
xor ( n66903 , n66900 , n66901 );
xor ( n66904 , n65717 , n65726 );
nor ( n66905 , n9716 , n66561 );
and ( n66906 , n66904 , n66905 );
xor ( n66907 , n66904 , n66905 );
xor ( n66908 , n65721 , n65724 );
nor ( n66909 , n9725 , n66561 );
and ( n66910 , n66908 , n66909 );
xor ( n66911 , n66908 , n66909 );
xor ( n66912 , n65722 , n65723 );
nor ( n66913 , n9734 , n66561 );
and ( n66914 , n66912 , n66913 );
xor ( n66915 , n66912 , n66913 );
nor ( n66916 , n9752 , n65371 );
nor ( n66917 , n9743 , n66561 );
and ( n66918 , n66916 , n66917 );
and ( n66919 , n66915 , n66918 );
or ( n66920 , n66914 , n66919 );
and ( n66921 , n66911 , n66920 );
or ( n66922 , n66910 , n66921 );
and ( n66923 , n66907 , n66922 );
or ( n66924 , n66906 , n66923 );
and ( n66925 , n66903 , n66924 );
or ( n66926 , n66902 , n66925 );
and ( n66927 , n66899 , n66926 );
or ( n66928 , n66898 , n66927 );
and ( n66929 , n66895 , n66928 );
or ( n66930 , n66894 , n66929 );
and ( n66931 , n66891 , n66930 );
or ( n66932 , n66890 , n66931 );
and ( n66933 , n66887 , n66932 );
or ( n66934 , n66886 , n66933 );
and ( n66935 , n66883 , n66934 );
or ( n66936 , n66882 , n66935 );
and ( n66937 , n66879 , n66936 );
or ( n66938 , n66878 , n66937 );
and ( n66939 , n66875 , n66938 );
or ( n66940 , n66874 , n66939 );
and ( n66941 , n66871 , n66940 );
or ( n66942 , n66870 , n66941 );
and ( n66943 , n66867 , n66942 );
or ( n66944 , n66866 , n66943 );
and ( n66945 , n66863 , n66944 );
or ( n66946 , n66862 , n66945 );
and ( n66947 , n66859 , n66946 );
or ( n66948 , n66858 , n66947 );
and ( n66949 , n66855 , n66948 );
or ( n66950 , n66854 , n66949 );
and ( n66951 , n66851 , n66950 );
or ( n66952 , n66850 , n66951 );
and ( n66953 , n66847 , n66952 );
or ( n66954 , n66846 , n66953 );
and ( n66955 , n66843 , n66954 );
or ( n66956 , n66842 , n66955 );
and ( n66957 , n66839 , n66956 );
or ( n66958 , n66838 , n66957 );
and ( n66959 , n66835 , n66958 );
or ( n66960 , n66834 , n66959 );
and ( n66961 , n66831 , n66960 );
or ( n66962 , n66830 , n66961 );
and ( n66963 , n66827 , n66962 );
or ( n66964 , n66826 , n66963 );
and ( n66965 , n66823 , n66964 );
or ( n66966 , n66822 , n66965 );
and ( n66967 , n66819 , n66966 );
or ( n66968 , n66818 , n66967 );
and ( n66969 , n66815 , n66968 );
or ( n66970 , n66814 , n66969 );
and ( n66971 , n66811 , n66970 );
or ( n66972 , n66810 , n66971 );
and ( n66973 , n66807 , n66972 );
or ( n66974 , n66806 , n66973 );
and ( n66975 , n66803 , n66974 );
or ( n66976 , n66802 , n66975 );
and ( n66977 , n66799 , n66976 );
or ( n66978 , n66798 , n66977 );
and ( n66979 , n66795 , n66978 );
or ( n66980 , n66794 , n66979 );
and ( n66981 , n66791 , n66980 );
or ( n66982 , n66790 , n66981 );
and ( n66983 , n66787 , n66982 );
or ( n66984 , n66786 , n66983 );
and ( n66985 , n66783 , n66984 );
or ( n66986 , n66782 , n66985 );
and ( n66987 , n66779 , n66986 );
or ( n66988 , n66778 , n66987 );
and ( n66989 , n66775 , n66988 );
or ( n66990 , n66774 , n66989 );
and ( n66991 , n66771 , n66990 );
or ( n66992 , n66770 , n66991 );
and ( n66993 , n66767 , n66992 );
or ( n66994 , n66766 , n66993 );
and ( n66995 , n66763 , n66994 );
or ( n66996 , n66762 , n66995 );
and ( n66997 , n66759 , n66996 );
or ( n66998 , n66758 , n66997 );
and ( n66999 , n66755 , n66998 );
or ( n67000 , n66754 , n66999 );
and ( n67001 , n66751 , n67000 );
or ( n67002 , n66750 , n67001 );
and ( n67003 , n66747 , n67002 );
or ( n67004 , n66746 , n67003 );
and ( n67005 , n66743 , n67004 );
or ( n67006 , n66742 , n67005 );
and ( n67007 , n66739 , n67006 );
or ( n67008 , n66738 , n67007 );
and ( n67009 , n66735 , n67008 );
or ( n67010 , n66734 , n67009 );
and ( n67011 , n66731 , n67010 );
or ( n67012 , n66730 , n67011 );
and ( n67013 , n66727 , n67012 );
or ( n67014 , n66726 , n67013 );
and ( n67015 , n66723 , n67014 );
or ( n67016 , n66722 , n67015 );
and ( n67017 , n66719 , n67016 );
or ( n67018 , n66718 , n67017 );
and ( n67019 , n66715 , n67018 );
or ( n67020 , n66714 , n67019 );
and ( n67021 , n66711 , n67020 );
or ( n67022 , n66710 , n67021 );
and ( n67023 , n66707 , n67022 );
or ( n67024 , n66706 , n67023 );
and ( n67025 , n66703 , n67024 );
or ( n67026 , n66702 , n67025 );
and ( n67027 , n66699 , n67026 );
or ( n67028 , n66698 , n67027 );
and ( n67029 , n66695 , n67028 );
or ( n67030 , n66694 , n67029 );
and ( n67031 , n66691 , n67030 );
or ( n67032 , n66690 , n67031 );
and ( n67033 , n66687 , n67032 );
or ( n67034 , n66686 , n67033 );
and ( n67035 , n66683 , n67034 );
or ( n67036 , n66682 , n67035 );
and ( n67037 , n66679 , n67036 );
or ( n67038 , n66678 , n67037 );
and ( n67039 , n66675 , n67038 );
or ( n67040 , n66674 , n67039 );
and ( n67041 , n66671 , n67040 );
or ( n67042 , n66670 , n67041 );
and ( n67043 , n66667 , n67042 );
or ( n67044 , n66666 , n67043 );
and ( n67045 , n66663 , n67044 );
or ( n67046 , n66662 , n67045 );
and ( n67047 , n66659 , n67046 );
or ( n67048 , n66658 , n67047 );
and ( n67049 , n66655 , n67048 );
or ( n67050 , n66654 , n67049 );
and ( n67051 , n66651 , n67050 );
or ( n67052 , n66650 , n67051 );
and ( n67053 , n66647 , n67052 );
or ( n67054 , n66646 , n67053 );
and ( n67055 , n66643 , n67054 );
or ( n67056 , n66642 , n67055 );
and ( n67057 , n66639 , n67056 );
or ( n67058 , n66638 , n67057 );
and ( n67059 , n66635 , n67058 );
or ( n67060 , n66634 , n67059 );
and ( n67061 , n66631 , n67060 );
or ( n67062 , n66630 , n67061 );
and ( n67063 , n66627 , n67062 );
or ( n67064 , n66626 , n67063 );
and ( n67065 , n66623 , n67064 );
or ( n67066 , n66622 , n67065 );
and ( n67067 , n66619 , n67066 );
or ( n67068 , n66618 , n67067 );
and ( n67069 , n66615 , n67068 );
or ( n67070 , n66614 , n67069 );
and ( n67071 , n66611 , n67070 );
or ( n67072 , n66610 , n67071 );
and ( n67073 , n66607 , n67072 );
or ( n67074 , n66606 , n67073 );
and ( n67075 , n66603 , n67074 );
or ( n67076 , n66602 , n67075 );
and ( n67077 , n66599 , n67076 );
or ( n67078 , n66598 , n67077 );
and ( n67079 , n66595 , n67078 );
or ( n67080 , n66594 , n67079 );
and ( n67081 , n66591 , n67080 );
or ( n67082 , n66590 , n67081 );
and ( n67083 , n66587 , n67082 );
or ( n67084 , n66586 , n67083 );
and ( n67085 , n66583 , n67084 );
or ( n67086 , n66582 , n67085 );
and ( n67087 , n66579 , n67086 );
or ( n67088 , n66578 , n67087 );
and ( n67089 , n66575 , n67088 );
or ( n67090 , n66574 , n67089 );
and ( n67091 , n66571 , n67090 );
or ( n67092 , n66570 , n67091 );
and ( n67093 , n66567 , n67092 );
or ( n67094 , n66566 , n67093 );
xor ( n67095 , n66563 , n67094 );
and ( n67096 , n33403 , n5476 );
nor ( n67097 , n5477 , n67096 );
nor ( n67098 , n5838 , n32231 );
xor ( n67099 , n67097 , n67098 );
and ( n67100 , n65901 , n65902 );
and ( n67101 , n65903 , n65906 );
or ( n67102 , n67100 , n67101 );
xor ( n67103 , n67099 , n67102 );
nor ( n67104 , n6212 , n31083 );
xor ( n67105 , n67103 , n67104 );
and ( n67106 , n65907 , n65908 );
and ( n67107 , n65909 , n65912 );
or ( n67108 , n67106 , n67107 );
xor ( n67109 , n67105 , n67108 );
nor ( n67110 , n6596 , n29948 );
xor ( n67111 , n67109 , n67110 );
and ( n67112 , n65913 , n65914 );
and ( n67113 , n65915 , n65918 );
or ( n67114 , n67112 , n67113 );
xor ( n67115 , n67111 , n67114 );
nor ( n67116 , n6997 , n28833 );
xor ( n67117 , n67115 , n67116 );
and ( n67118 , n65919 , n65920 );
and ( n67119 , n65921 , n65924 );
or ( n67120 , n67118 , n67119 );
xor ( n67121 , n67117 , n67120 );
nor ( n67122 , n7413 , n27737 );
xor ( n67123 , n67121 , n67122 );
and ( n67124 , n65925 , n65926 );
and ( n67125 , n65927 , n65930 );
or ( n67126 , n67124 , n67125 );
xor ( n67127 , n67123 , n67126 );
nor ( n67128 , n7841 , n26660 );
xor ( n67129 , n67127 , n67128 );
and ( n67130 , n65931 , n65932 );
and ( n67131 , n65933 , n65936 );
or ( n67132 , n67130 , n67131 );
xor ( n67133 , n67129 , n67132 );
nor ( n67134 , n8281 , n25600 );
xor ( n67135 , n67133 , n67134 );
and ( n67136 , n65937 , n65938 );
and ( n67137 , n65939 , n65942 );
or ( n67138 , n67136 , n67137 );
xor ( n67139 , n67135 , n67138 );
nor ( n67140 , n8737 , n24564 );
xor ( n67141 , n67139 , n67140 );
and ( n67142 , n65943 , n65944 );
and ( n67143 , n65945 , n65948 );
or ( n67144 , n67142 , n67143 );
xor ( n67145 , n67141 , n67144 );
nor ( n67146 , n9420 , n23541 );
xor ( n67147 , n67145 , n67146 );
and ( n67148 , n65949 , n65950 );
and ( n67149 , n65951 , n65954 );
or ( n67150 , n67148 , n67149 );
xor ( n67151 , n67147 , n67150 );
nor ( n67152 , n10312 , n22541 );
xor ( n67153 , n67151 , n67152 );
and ( n67154 , n65955 , n65956 );
and ( n67155 , n65957 , n65960 );
or ( n67156 , n67154 , n67155 );
xor ( n67157 , n67153 , n67156 );
nor ( n67158 , n11041 , n21562 );
xor ( n67159 , n67157 , n67158 );
and ( n67160 , n65961 , n65962 );
and ( n67161 , n65963 , n65966 );
or ( n67162 , n67160 , n67161 );
xor ( n67163 , n67159 , n67162 );
nor ( n67164 , n11790 , n20601 );
xor ( n67165 , n67163 , n67164 );
and ( n67166 , n65967 , n65968 );
and ( n67167 , n65969 , n65972 );
or ( n67168 , n67166 , n67167 );
xor ( n67169 , n67165 , n67168 );
nor ( n67170 , n12555 , n19657 );
xor ( n67171 , n67169 , n67170 );
and ( n67172 , n65973 , n65974 );
and ( n67173 , n65975 , n65978 );
or ( n67174 , n67172 , n67173 );
xor ( n67175 , n67171 , n67174 );
nor ( n67176 , n13340 , n18734 );
xor ( n67177 , n67175 , n67176 );
and ( n67178 , n65979 , n65980 );
and ( n67179 , n65981 , n65984 );
or ( n67180 , n67178 , n67179 );
xor ( n67181 , n67177 , n67180 );
nor ( n67182 , n14138 , n17828 );
xor ( n67183 , n67181 , n67182 );
and ( n67184 , n65985 , n65986 );
and ( n67185 , n65987 , n65990 );
or ( n67186 , n67184 , n67185 );
xor ( n67187 , n67183 , n67186 );
nor ( n67188 , n14959 , n16943 );
xor ( n67189 , n67187 , n67188 );
and ( n67190 , n65991 , n65992 );
and ( n67191 , n65993 , n65996 );
or ( n67192 , n67190 , n67191 );
xor ( n67193 , n67189 , n67192 );
nor ( n67194 , n15800 , n16077 );
xor ( n67195 , n67193 , n67194 );
and ( n67196 , n65997 , n65998 );
and ( n67197 , n65999 , n66002 );
or ( n67198 , n67196 , n67197 );
xor ( n67199 , n67195 , n67198 );
nor ( n67200 , n16660 , n15230 );
xor ( n67201 , n67199 , n67200 );
and ( n67202 , n66003 , n66004 );
and ( n67203 , n66005 , n66008 );
or ( n67204 , n67202 , n67203 );
xor ( n67205 , n67201 , n67204 );
nor ( n67206 , n17539 , n14403 );
xor ( n67207 , n67205 , n67206 );
and ( n67208 , n66009 , n66010 );
and ( n67209 , n66011 , n66014 );
or ( n67210 , n67208 , n67209 );
xor ( n67211 , n67207 , n67210 );
nor ( n67212 , n18439 , n13599 );
xor ( n67213 , n67211 , n67212 );
and ( n67214 , n66015 , n66016 );
and ( n67215 , n66017 , n66020 );
or ( n67216 , n67214 , n67215 );
xor ( n67217 , n67213 , n67216 );
nor ( n67218 , n19356 , n12808 );
xor ( n67219 , n67217 , n67218 );
and ( n67220 , n66021 , n66022 );
and ( n67221 , n66023 , n66026 );
or ( n67222 , n67220 , n67221 );
xor ( n67223 , n67219 , n67222 );
nor ( n67224 , n20294 , n12037 );
xor ( n67225 , n67223 , n67224 );
and ( n67226 , n66027 , n66028 );
and ( n67227 , n66029 , n66032 );
or ( n67228 , n67226 , n67227 );
xor ( n67229 , n67225 , n67228 );
nor ( n67230 , n21249 , n11282 );
xor ( n67231 , n67229 , n67230 );
and ( n67232 , n66033 , n66034 );
and ( n67233 , n66035 , n66038 );
or ( n67234 , n67232 , n67233 );
xor ( n67235 , n67231 , n67234 );
nor ( n67236 , n22222 , n10547 );
xor ( n67237 , n67235 , n67236 );
and ( n67238 , n66039 , n66040 );
and ( n67239 , n66041 , n66044 );
or ( n67240 , n67238 , n67239 );
xor ( n67241 , n67237 , n67240 );
nor ( n67242 , n23216 , n9829 );
xor ( n67243 , n67241 , n67242 );
and ( n67244 , n66045 , n66046 );
and ( n67245 , n66047 , n66050 );
or ( n67246 , n67244 , n67245 );
xor ( n67247 , n67243 , n67246 );
nor ( n67248 , n24233 , n8955 );
xor ( n67249 , n67247 , n67248 );
and ( n67250 , n66051 , n66052 );
and ( n67251 , n66053 , n66056 );
or ( n67252 , n67250 , n67251 );
xor ( n67253 , n67249 , n67252 );
nor ( n67254 , n25263 , n603 );
xor ( n67255 , n67253 , n67254 );
and ( n67256 , n66057 , n66058 );
and ( n67257 , n66059 , n66062 );
or ( n67258 , n67256 , n67257 );
xor ( n67259 , n67255 , n67258 );
nor ( n67260 , n26317 , n652 );
xor ( n67261 , n67259 , n67260 );
and ( n67262 , n66063 , n66064 );
and ( n67263 , n66065 , n66068 );
or ( n67264 , n67262 , n67263 );
xor ( n67265 , n67261 , n67264 );
nor ( n67266 , n27388 , n624 );
xor ( n67267 , n67265 , n67266 );
and ( n67268 , n66069 , n66070 );
and ( n67269 , n66071 , n66074 );
or ( n67270 , n67268 , n67269 );
xor ( n67271 , n67267 , n67270 );
nor ( n67272 , n28478 , n648 );
xor ( n67273 , n67271 , n67272 );
and ( n67274 , n66075 , n66076 );
and ( n67275 , n66077 , n66080 );
or ( n67276 , n67274 , n67275 );
xor ( n67277 , n67273 , n67276 );
nor ( n67278 , n29587 , n686 );
xor ( n67279 , n67277 , n67278 );
and ( n67280 , n66081 , n66082 );
and ( n67281 , n66083 , n66086 );
or ( n67282 , n67280 , n67281 );
xor ( n67283 , n67279 , n67282 );
nor ( n67284 , n30716 , n735 );
xor ( n67285 , n67283 , n67284 );
and ( n67286 , n66087 , n66088 );
and ( n67287 , n66089 , n66092 );
or ( n67288 , n67286 , n67287 );
xor ( n67289 , n67285 , n67288 );
nor ( n67290 , n31858 , n798 );
xor ( n67291 , n67289 , n67290 );
and ( n67292 , n66093 , n66094 );
and ( n67293 , n66095 , n66098 );
or ( n67294 , n67292 , n67293 );
xor ( n67295 , n67291 , n67294 );
nor ( n67296 , n33024 , n870 );
xor ( n67297 , n67295 , n67296 );
and ( n67298 , n66099 , n66100 );
and ( n67299 , n66101 , n66104 );
or ( n67300 , n67298 , n67299 );
xor ( n67301 , n67297 , n67300 );
nor ( n67302 , n34215 , n960 );
xor ( n67303 , n67301 , n67302 );
and ( n67304 , n66105 , n66106 );
and ( n67305 , n66107 , n66110 );
or ( n67306 , n67304 , n67305 );
xor ( n67307 , n67303 , n67306 );
nor ( n67308 , n35410 , n1064 );
xor ( n67309 , n67307 , n67308 );
and ( n67310 , n66111 , n66112 );
and ( n67311 , n66113 , n66116 );
or ( n67312 , n67310 , n67311 );
xor ( n67313 , n67309 , n67312 );
nor ( n67314 , n36611 , n1178 );
xor ( n67315 , n67313 , n67314 );
and ( n67316 , n66117 , n66118 );
and ( n67317 , n66119 , n66122 );
or ( n67318 , n67316 , n67317 );
xor ( n67319 , n67315 , n67318 );
nor ( n67320 , n37816 , n1305 );
xor ( n67321 , n67319 , n67320 );
and ( n67322 , n66123 , n66124 );
and ( n67323 , n66125 , n66128 );
or ( n67324 , n67322 , n67323 );
xor ( n67325 , n67321 , n67324 );
nor ( n67326 , n39018 , n1447 );
xor ( n67327 , n67325 , n67326 );
and ( n67328 , n66129 , n66130 );
and ( n67329 , n66131 , n66134 );
or ( n67330 , n67328 , n67329 );
xor ( n67331 , n67327 , n67330 );
nor ( n67332 , n40223 , n1600 );
xor ( n67333 , n67331 , n67332 );
and ( n67334 , n66135 , n66136 );
and ( n67335 , n66137 , n66140 );
or ( n67336 , n67334 , n67335 );
xor ( n67337 , n67333 , n67336 );
nor ( n67338 , n41428 , n1768 );
xor ( n67339 , n67337 , n67338 );
and ( n67340 , n66141 , n66142 );
and ( n67341 , n66143 , n66146 );
or ( n67342 , n67340 , n67341 );
xor ( n67343 , n67339 , n67342 );
nor ( n67344 , n42632 , n1947 );
xor ( n67345 , n67343 , n67344 );
and ( n67346 , n66147 , n66148 );
and ( n67347 , n66149 , n66152 );
or ( n67348 , n67346 , n67347 );
xor ( n67349 , n67345 , n67348 );
nor ( n67350 , n43834 , n2139 );
xor ( n67351 , n67349 , n67350 );
and ( n67352 , n66153 , n66154 );
and ( n67353 , n66155 , n66158 );
or ( n67354 , n67352 , n67353 );
xor ( n67355 , n67351 , n67354 );
nor ( n67356 , n45038 , n2345 );
xor ( n67357 , n67355 , n67356 );
and ( n67358 , n66159 , n66160 );
and ( n67359 , n66161 , n66164 );
or ( n67360 , n67358 , n67359 );
xor ( n67361 , n67357 , n67360 );
nor ( n67362 , n46239 , n2568 );
xor ( n67363 , n67361 , n67362 );
and ( n67364 , n66165 , n66166 );
and ( n67365 , n66167 , n66170 );
or ( n67366 , n67364 , n67365 );
xor ( n67367 , n67363 , n67366 );
nor ( n67368 , n47440 , n2799 );
xor ( n67369 , n67367 , n67368 );
and ( n67370 , n66171 , n66172 );
and ( n67371 , n66173 , n66176 );
or ( n67372 , n67370 , n67371 );
xor ( n67373 , n67369 , n67372 );
nor ( n67374 , n48641 , n3045 );
xor ( n67375 , n67373 , n67374 );
and ( n67376 , n66177 , n66178 );
and ( n67377 , n66179 , n66182 );
or ( n67378 , n67376 , n67377 );
xor ( n67379 , n67375 , n67378 );
nor ( n67380 , n49841 , n3302 );
xor ( n67381 , n67379 , n67380 );
and ( n67382 , n66183 , n66184 );
and ( n67383 , n66185 , n66188 );
or ( n67384 , n67382 , n67383 );
xor ( n67385 , n67381 , n67384 );
nor ( n67386 , n51040 , n3572 );
xor ( n67387 , n67385 , n67386 );
and ( n67388 , n66189 , n66190 );
and ( n67389 , n66191 , n66194 );
or ( n67390 , n67388 , n67389 );
xor ( n67391 , n67387 , n67390 );
nor ( n67392 , n52238 , n3855 );
xor ( n67393 , n67391 , n67392 );
and ( n67394 , n66195 , n66196 );
and ( n67395 , n66197 , n66200 );
or ( n67396 , n67394 , n67395 );
xor ( n67397 , n67393 , n67396 );
nor ( n67398 , n53432 , n4153 );
xor ( n67399 , n67397 , n67398 );
and ( n67400 , n66201 , n66202 );
and ( n67401 , n66203 , n66206 );
or ( n67402 , n67400 , n67401 );
xor ( n67403 , n67399 , n67402 );
nor ( n67404 , n54629 , n4460 );
xor ( n67405 , n67403 , n67404 );
and ( n67406 , n66207 , n66208 );
and ( n67407 , n66209 , n66212 );
or ( n67408 , n67406 , n67407 );
xor ( n67409 , n67405 , n67408 );
nor ( n67410 , n55826 , n4788 );
xor ( n67411 , n67409 , n67410 );
and ( n67412 , n66213 , n66214 );
and ( n67413 , n66215 , n66218 );
or ( n67414 , n67412 , n67413 );
xor ( n67415 , n67411 , n67414 );
nor ( n67416 , n57022 , n5128 );
xor ( n67417 , n67415 , n67416 );
and ( n67418 , n66219 , n66220 );
and ( n67419 , n66221 , n66224 );
or ( n67420 , n67418 , n67419 );
xor ( n67421 , n67417 , n67420 );
nor ( n67422 , n58217 , n5479 );
xor ( n67423 , n67421 , n67422 );
and ( n67424 , n66225 , n66226 );
and ( n67425 , n66227 , n66230 );
or ( n67426 , n67424 , n67425 );
xor ( n67427 , n67423 , n67426 );
nor ( n67428 , n59412 , n5840 );
xor ( n67429 , n67427 , n67428 );
and ( n67430 , n66231 , n66232 );
and ( n67431 , n66233 , n66236 );
or ( n67432 , n67430 , n67431 );
xor ( n67433 , n67429 , n67432 );
nor ( n67434 , n60600 , n6214 );
xor ( n67435 , n67433 , n67434 );
and ( n67436 , n66237 , n66238 );
and ( n67437 , n66239 , n66242 );
or ( n67438 , n67436 , n67437 );
xor ( n67439 , n67435 , n67438 );
nor ( n67440 , n61791 , n6598 );
xor ( n67441 , n67439 , n67440 );
and ( n67442 , n66243 , n66244 );
and ( n67443 , n66245 , n66248 );
or ( n67444 , n67442 , n67443 );
xor ( n67445 , n67441 , n67444 );
nor ( n67446 , n62982 , n6999 );
xor ( n67447 , n67445 , n67446 );
and ( n67448 , n66249 , n66250 );
and ( n67449 , n66251 , n66254 );
or ( n67450 , n67448 , n67449 );
xor ( n67451 , n67447 , n67450 );
nor ( n67452 , n64172 , n7415 );
xor ( n67453 , n67451 , n67452 );
and ( n67454 , n66255 , n66256 );
and ( n67455 , n66257 , n66260 );
or ( n67456 , n67454 , n67455 );
xor ( n67457 , n67453 , n67456 );
nor ( n67458 , n65360 , n7843 );
xor ( n67459 , n67457 , n67458 );
and ( n67460 , n66261 , n66262 );
and ( n67461 , n66263 , n66266 );
or ( n67462 , n67460 , n67461 );
xor ( n67463 , n67459 , n67462 );
nor ( n67464 , n66550 , n8283 );
xor ( n67465 , n67463 , n67464 );
and ( n67466 , n66267 , n66268 );
and ( n67467 , n66269 , n66272 );
or ( n67468 , n67466 , n67467 );
xor ( n67469 , n67465 , n67468 );
and ( n67470 , n66285 , n66289 );
and ( n67471 , n66289 , n66536 );
and ( n67472 , n66285 , n66536 );
or ( n67473 , n67470 , n67471 , n67472 );
and ( n67474 , n33774 , n5408 );
not ( n67475 , n5408 );
nor ( n67476 , n67474 , n67475 );
xor ( n67477 , n67473 , n67476 );
and ( n67478 , n66295 , n66299 );
and ( n67479 , n66299 , n66367 );
and ( n67480 , n66295 , n66367 );
or ( n67481 , n67478 , n67479 , n67480 );
and ( n67482 , n66291 , n66368 );
and ( n67483 , n66368 , n66535 );
and ( n67484 , n66291 , n66535 );
or ( n67485 , n67482 , n67483 , n67484 );
xor ( n67486 , n67481 , n67485 );
and ( n67487 , n66486 , n66534 );
and ( n67488 , n66373 , n66374 );
and ( n67489 , n66374 , n66485 );
and ( n67490 , n66373 , n66485 );
or ( n67491 , n67488 , n67489 , n67490 );
and ( n67492 , n66304 , n66308 );
and ( n67493 , n66308 , n66366 );
and ( n67494 , n66304 , n66366 );
or ( n67495 , n67492 , n67493 , n67494 );
xor ( n67496 , n67491 , n67495 );
and ( n67497 , n66335 , n66339 );
and ( n67498 , n66339 , n66345 );
and ( n67499 , n66335 , n66345 );
or ( n67500 , n67497 , n67498 , n67499 );
and ( n67501 , n66313 , n66317 );
and ( n67502 , n66317 , n66365 );
and ( n67503 , n66313 , n66365 );
or ( n67504 , n67501 , n67502 , n67503 );
xor ( n67505 , n67500 , n67504 );
and ( n67506 , n66322 , n66326 );
and ( n67507 , n66326 , n66364 );
and ( n67508 , n66322 , n66364 );
or ( n67509 , n67506 , n67507 , n67508 );
and ( n67510 , n66383 , n66408 );
and ( n67511 , n66408 , n66446 );
and ( n67512 , n66383 , n66446 );
or ( n67513 , n67510 , n67511 , n67512 );
xor ( n67514 , n67509 , n67513 );
and ( n67515 , n66331 , n66346 );
and ( n67516 , n66346 , n66363 );
and ( n67517 , n66331 , n66363 );
or ( n67518 , n67515 , n67516 , n67517 );
and ( n67519 , n66387 , n66391 );
and ( n67520 , n66391 , n66407 );
and ( n67521 , n66387 , n66407 );
or ( n67522 , n67519 , n67520 , n67521 );
xor ( n67523 , n67518 , n67522 );
and ( n67524 , n66351 , n66356 );
and ( n67525 , n66356 , n66362 );
and ( n67526 , n66351 , n66362 );
or ( n67527 , n67524 , n67525 , n67526 );
and ( n67528 , n66341 , n66342 );
and ( n67529 , n66342 , n66344 );
and ( n67530 , n66341 , n66344 );
or ( n67531 , n67528 , n67529 , n67530 );
and ( n67532 , n66352 , n66353 );
and ( n67533 , n66353 , n66355 );
and ( n67534 , n66352 , n66355 );
or ( n67535 , n67532 , n67533 , n67534 );
xor ( n67536 , n67531 , n67535 );
and ( n67537 , n30695 , n6504 );
and ( n67538 , n31836 , n6132 );
xor ( n67539 , n67537 , n67538 );
and ( n67540 , n32649 , n5765 );
xor ( n67541 , n67539 , n67540 );
xor ( n67542 , n67536 , n67541 );
xor ( n67543 , n67527 , n67542 );
and ( n67544 , n66358 , n66359 );
and ( n67545 , n66359 , n66361 );
and ( n67546 , n66358 , n66361 );
or ( n67547 , n67544 , n67545 , n67546 );
and ( n67548 , n27361 , n7662 );
and ( n67549 , n28456 , n7310 );
xor ( n67550 , n67548 , n67549 );
and ( n67551 , n29559 , n6971 );
xor ( n67552 , n67550 , n67551 );
xor ( n67553 , n67547 , n67552 );
and ( n67554 , n24214 , n9348 );
and ( n67555 , n25243 , n8669 );
xor ( n67556 , n67554 , n67555 );
and ( n67557 , n26296 , n8243 );
xor ( n67558 , n67556 , n67557 );
xor ( n67559 , n67553 , n67558 );
xor ( n67560 , n67543 , n67559 );
xor ( n67561 , n67523 , n67560 );
xor ( n67562 , n67514 , n67561 );
xor ( n67563 , n67505 , n67562 );
xor ( n67564 , n67496 , n67563 );
xor ( n67565 , n67487 , n67564 );
and ( n67566 , n66379 , n66447 );
and ( n67567 , n66447 , n66484 );
and ( n67568 , n66379 , n66484 );
or ( n67569 , n67566 , n67567 , n67568 );
and ( n67570 , n66490 , n66533 );
xor ( n67571 , n67569 , n67570 );
and ( n67572 , n66452 , n66456 );
and ( n67573 , n66456 , n66483 );
and ( n67574 , n66452 , n66483 );
or ( n67575 , n67572 , n67573 , n67574 );
and ( n67576 , n66413 , n66429 );
and ( n67577 , n66429 , n66445 );
and ( n67578 , n66413 , n66445 );
or ( n67579 , n67576 , n67577 , n67578 );
and ( n67580 , n66396 , n66400 );
and ( n67581 , n66400 , n66406 );
and ( n67582 , n66396 , n66406 );
or ( n67583 , n67580 , n67581 , n67582 );
and ( n67584 , n66417 , n66422 );
and ( n67585 , n66422 , n66428 );
and ( n67586 , n66417 , n66428 );
or ( n67587 , n67584 , n67585 , n67586 );
xor ( n67588 , n67583 , n67587 );
and ( n67589 , n66402 , n66403 );
and ( n67590 , n66403 , n66405 );
and ( n67591 , n66402 , n66405 );
or ( n67592 , n67589 , n67590 , n67591 );
and ( n67593 , n66418 , n66419 );
and ( n67594 , n66419 , n66421 );
and ( n67595 , n66418 , n66421 );
or ( n67596 , n67593 , n67594 , n67595 );
xor ( n67597 , n67592 , n67596 );
and ( n67598 , n21216 , n11718 );
and ( n67599 , n22186 , n10977 );
xor ( n67600 , n67598 , n67599 );
and ( n67601 , n22892 , n10239 );
xor ( n67602 , n67600 , n67601 );
xor ( n67603 , n67597 , n67602 );
xor ( n67604 , n67588 , n67603 );
xor ( n67605 , n67579 , n67604 );
and ( n67606 , n66434 , n66438 );
and ( n67607 , n66438 , n66444 );
and ( n67608 , n66434 , n66444 );
or ( n67609 , n67606 , n67607 , n67608 );
and ( n67610 , n66424 , n66425 );
and ( n67611 , n66425 , n66427 );
and ( n67612 , n66424 , n66427 );
or ( n67613 , n67610 , n67611 , n67612 );
and ( n67614 , n18144 , n14044 );
and ( n67615 , n19324 , n13256 );
xor ( n67616 , n67614 , n67615 );
and ( n67617 , n20233 , n12531 );
xor ( n67618 , n67616 , n67617 );
xor ( n67619 , n67613 , n67618 );
and ( n67620 , n17512 , n14838 );
buf ( n67621 , n67620 );
xor ( n67622 , n67619 , n67621 );
xor ( n67623 , n67609 , n67622 );
and ( n67624 , n66440 , n66441 );
and ( n67625 , n66441 , n66443 );
and ( n67626 , n66440 , n66443 );
or ( n67627 , n67624 , n67625 , n67626 );
and ( n67628 , n66471 , n66472 );
and ( n67629 , n66472 , n66474 );
and ( n67630 , n66471 , n66474 );
or ( n67631 , n67628 , n67629 , n67630 );
xor ( n67632 , n67627 , n67631 );
and ( n67633 , n13322 , n19222 );
and ( n67634 , n14118 , n18407 );
xor ( n67635 , n67633 , n67634 );
and ( n67636 , n14938 , n17422 );
xor ( n67637 , n67635 , n67636 );
xor ( n67638 , n67632 , n67637 );
xor ( n67639 , n67623 , n67638 );
xor ( n67640 , n67605 , n67639 );
xor ( n67641 , n67575 , n67640 );
and ( n67642 , n66461 , n66465 );
and ( n67643 , n66465 , n66482 );
and ( n67644 , n66461 , n66482 );
or ( n67645 , n67642 , n67643 , n67644 );
and ( n67646 , n66497 , n66512 );
and ( n67647 , n66512 , n66531 );
and ( n67648 , n66497 , n66531 );
or ( n67649 , n67646 , n67647 , n67648 );
xor ( n67650 , n67645 , n67649 );
and ( n67651 , n66470 , n66475 );
and ( n67652 , n66475 , n66481 );
and ( n67653 , n66470 , n66481 );
or ( n67654 , n67651 , n67652 , n67653 );
and ( n67655 , n66501 , n66505 );
and ( n67656 , n66505 , n66511 );
and ( n67657 , n66501 , n66511 );
or ( n67658 , n67655 , n67656 , n67657 );
xor ( n67659 , n67654 , n67658 );
and ( n67660 , n66477 , n66478 );
and ( n67661 , n66478 , n66480 );
and ( n67662 , n66477 , n66480 );
or ( n67663 , n67660 , n67661 , n67662 );
and ( n67664 , n11015 , n22065 );
and ( n67665 , n11769 , n20976 );
xor ( n67666 , n67664 , n67665 );
and ( n67667 , n12320 , n20156 );
xor ( n67668 , n67666 , n67667 );
xor ( n67669 , n67663 , n67668 );
and ( n67670 , n8718 , n25163 );
and ( n67671 , n9400 , n24137 );
xor ( n67672 , n67670 , n67671 );
and ( n67673 , n10291 , n23075 );
xor ( n67674 , n67672 , n67673 );
xor ( n67675 , n67669 , n67674 );
xor ( n67676 , n67659 , n67675 );
xor ( n67677 , n67650 , n67676 );
xor ( n67678 , n67641 , n67677 );
xor ( n67679 , n67571 , n67678 );
and ( n67680 , n66492 , n66532 );
and ( n67681 , n66491 , n66532 );
or ( n67682 , 1'b0 , n67680 , n67681 );
and ( n67683 , n66517 , n66522 );
and ( n67684 , n66522 , n66530 );
and ( n67685 , n66517 , n66530 );
or ( n67686 , n67683 , n67684 , n67685 );
and ( n67687 , n66507 , n66508 );
and ( n67688 , n66508 , n66510 );
and ( n67689 , n66507 , n66510 );
or ( n67690 , n67687 , n67688 , n67689 );
and ( n67691 , n66518 , n66519 );
and ( n67692 , n66519 , n66521 );
and ( n67693 , n66518 , n66521 );
or ( n67694 , n67691 , n67692 , n67693 );
xor ( n67695 , n67690 , n67694 );
and ( n67696 , n7385 , n28406 );
and ( n67697 , n7808 , n27296 );
xor ( n67698 , n67696 , n67697 );
and ( n67699 , n8079 , n26216 );
xor ( n67700 , n67698 , n67699 );
xor ( n67701 , n67695 , n67700 );
xor ( n67702 , n67686 , n67701 );
and ( n67703 , n66526 , n66527 );
and ( n67704 , n66527 , n66529 );
and ( n67705 , n66526 , n66529 );
or ( n67706 , n67703 , n67704 , n67705 );
and ( n67707 , n6187 , n31761 );
and ( n67708 , n6569 , n30629 );
xor ( n67709 , n67707 , n67708 );
and ( n67710 , n6816 , n29508 );
xor ( n67711 , n67709 , n67710 );
xor ( n67712 , n67706 , n67711 );
not ( n67713 , n5459 );
and ( n67714 , n34193 , n5459 );
nor ( n67715 , n67713 , n67714 );
and ( n67716 , n5819 , n32999 );
xor ( n67717 , n67715 , n67716 );
xor ( n67718 , n67712 , n67717 );
xor ( n67719 , n67702 , n67718 );
xor ( n67720 , n67682 , n67719 );
xor ( n67721 , n67679 , n67720 );
xor ( n67722 , n67565 , n67721 );
xor ( n67723 , n67486 , n67722 );
xor ( n67724 , n67477 , n67723 );
and ( n67725 , n66277 , n66280 );
and ( n67726 , n66280 , n66537 );
and ( n67727 , n66277 , n66537 );
or ( n67728 , n67725 , n67726 , n67727 );
xor ( n67729 , n67724 , n67728 );
and ( n67730 , n66538 , n66542 );
and ( n67731 , n66543 , n66546 );
or ( n67732 , n67730 , n67731 );
xor ( n67733 , n67729 , n67732 );
buf ( n67734 , n67733 );
buf ( n67735 , n67734 );
not ( n67736 , n67735 );
nor ( n67737 , n67736 , n8739 );
xor ( n67738 , n67469 , n67737 );
and ( n67739 , n66273 , n66551 );
and ( n67740 , n66552 , n66555 );
or ( n67741 , n67739 , n67740 );
xor ( n67742 , n67738 , n67741 );
buf ( n67743 , n67742 );
buf ( n67744 , n67743 );
not ( n67745 , n67744 );
buf ( n67746 , n590 );
not ( n67747 , n67746 );
nor ( n67748 , n67745 , n67747 );
xor ( n67749 , n67095 , n67748 );
xor ( n67750 , n66567 , n67092 );
nor ( n67751 , n66559 , n67747 );
and ( n67752 , n67750 , n67751 );
xor ( n67753 , n67750 , n67751 );
xor ( n67754 , n66571 , n67090 );
nor ( n67755 , n65369 , n67747 );
and ( n67756 , n67754 , n67755 );
xor ( n67757 , n67754 , n67755 );
xor ( n67758 , n66575 , n67088 );
nor ( n67759 , n64181 , n67747 );
and ( n67760 , n67758 , n67759 );
xor ( n67761 , n67758 , n67759 );
xor ( n67762 , n66579 , n67086 );
nor ( n67763 , n62991 , n67747 );
and ( n67764 , n67762 , n67763 );
xor ( n67765 , n67762 , n67763 );
xor ( n67766 , n66583 , n67084 );
nor ( n67767 , n61800 , n67747 );
and ( n67768 , n67766 , n67767 );
xor ( n67769 , n67766 , n67767 );
xor ( n67770 , n66587 , n67082 );
nor ( n67771 , n60609 , n67747 );
and ( n67772 , n67770 , n67771 );
xor ( n67773 , n67770 , n67771 );
xor ( n67774 , n66591 , n67080 );
nor ( n67775 , n59421 , n67747 );
and ( n67776 , n67774 , n67775 );
xor ( n67777 , n67774 , n67775 );
xor ( n67778 , n66595 , n67078 );
nor ( n67779 , n58226 , n67747 );
and ( n67780 , n67778 , n67779 );
xor ( n67781 , n67778 , n67779 );
xor ( n67782 , n66599 , n67076 );
nor ( n67783 , n57031 , n67747 );
and ( n67784 , n67782 , n67783 );
xor ( n67785 , n67782 , n67783 );
xor ( n67786 , n66603 , n67074 );
nor ( n67787 , n55835 , n67747 );
and ( n67788 , n67786 , n67787 );
xor ( n67789 , n67786 , n67787 );
xor ( n67790 , n66607 , n67072 );
nor ( n67791 , n54638 , n67747 );
and ( n67792 , n67790 , n67791 );
xor ( n67793 , n67790 , n67791 );
xor ( n67794 , n66611 , n67070 );
nor ( n67795 , n53441 , n67747 );
and ( n67796 , n67794 , n67795 );
xor ( n67797 , n67794 , n67795 );
xor ( n67798 , n66615 , n67068 );
nor ( n67799 , n52247 , n67747 );
and ( n67800 , n67798 , n67799 );
xor ( n67801 , n67798 , n67799 );
xor ( n67802 , n66619 , n67066 );
nor ( n67803 , n51049 , n67747 );
and ( n67804 , n67802 , n67803 );
xor ( n67805 , n67802 , n67803 );
xor ( n67806 , n66623 , n67064 );
nor ( n67807 , n49850 , n67747 );
and ( n67808 , n67806 , n67807 );
xor ( n67809 , n67806 , n67807 );
xor ( n67810 , n66627 , n67062 );
nor ( n67811 , n48650 , n67747 );
and ( n67812 , n67810 , n67811 );
xor ( n67813 , n67810 , n67811 );
xor ( n67814 , n66631 , n67060 );
nor ( n67815 , n47449 , n67747 );
and ( n67816 , n67814 , n67815 );
xor ( n67817 , n67814 , n67815 );
xor ( n67818 , n66635 , n67058 );
nor ( n67819 , n46248 , n67747 );
and ( n67820 , n67818 , n67819 );
xor ( n67821 , n67818 , n67819 );
xor ( n67822 , n66639 , n67056 );
nor ( n67823 , n45047 , n67747 );
and ( n67824 , n67822 , n67823 );
xor ( n67825 , n67822 , n67823 );
xor ( n67826 , n66643 , n67054 );
nor ( n67827 , n43843 , n67747 );
and ( n67828 , n67826 , n67827 );
xor ( n67829 , n67826 , n67827 );
xor ( n67830 , n66647 , n67052 );
nor ( n67831 , n42641 , n67747 );
and ( n67832 , n67830 , n67831 );
xor ( n67833 , n67830 , n67831 );
xor ( n67834 , n66651 , n67050 );
nor ( n67835 , n41437 , n67747 );
and ( n67836 , n67834 , n67835 );
xor ( n67837 , n67834 , n67835 );
xor ( n67838 , n66655 , n67048 );
nor ( n67839 , n40232 , n67747 );
and ( n67840 , n67838 , n67839 );
xor ( n67841 , n67838 , n67839 );
xor ( n67842 , n66659 , n67046 );
nor ( n67843 , n39027 , n67747 );
and ( n67844 , n67842 , n67843 );
xor ( n67845 , n67842 , n67843 );
xor ( n67846 , n66663 , n67044 );
nor ( n67847 , n37825 , n67747 );
and ( n67848 , n67846 , n67847 );
xor ( n67849 , n67846 , n67847 );
xor ( n67850 , n66667 , n67042 );
nor ( n67851 , n36620 , n67747 );
and ( n67852 , n67850 , n67851 );
xor ( n67853 , n67850 , n67851 );
xor ( n67854 , n66671 , n67040 );
nor ( n67855 , n35419 , n67747 );
and ( n67856 , n67854 , n67855 );
xor ( n67857 , n67854 , n67855 );
xor ( n67858 , n66675 , n67038 );
nor ( n67859 , n34224 , n67747 );
and ( n67860 , n67858 , n67859 );
xor ( n67861 , n67858 , n67859 );
xor ( n67862 , n66679 , n67036 );
nor ( n67863 , n33033 , n67747 );
and ( n67864 , n67862 , n67863 );
xor ( n67865 , n67862 , n67863 );
xor ( n67866 , n66683 , n67034 );
nor ( n67867 , n31867 , n67747 );
and ( n67868 , n67866 , n67867 );
xor ( n67869 , n67866 , n67867 );
xor ( n67870 , n66687 , n67032 );
nor ( n67871 , n30725 , n67747 );
and ( n67872 , n67870 , n67871 );
xor ( n67873 , n67870 , n67871 );
xor ( n67874 , n66691 , n67030 );
nor ( n67875 , n29596 , n67747 );
and ( n67876 , n67874 , n67875 );
xor ( n67877 , n67874 , n67875 );
xor ( n67878 , n66695 , n67028 );
nor ( n67879 , n28487 , n67747 );
and ( n67880 , n67878 , n67879 );
xor ( n67881 , n67878 , n67879 );
xor ( n67882 , n66699 , n67026 );
nor ( n67883 , n27397 , n67747 );
and ( n67884 , n67882 , n67883 );
xor ( n67885 , n67882 , n67883 );
xor ( n67886 , n66703 , n67024 );
nor ( n67887 , n26326 , n67747 );
and ( n67888 , n67886 , n67887 );
xor ( n67889 , n67886 , n67887 );
xor ( n67890 , n66707 , n67022 );
nor ( n67891 , n25272 , n67747 );
and ( n67892 , n67890 , n67891 );
xor ( n67893 , n67890 , n67891 );
xor ( n67894 , n66711 , n67020 );
nor ( n67895 , n24242 , n67747 );
and ( n67896 , n67894 , n67895 );
xor ( n67897 , n67894 , n67895 );
xor ( n67898 , n66715 , n67018 );
nor ( n67899 , n23225 , n67747 );
and ( n67900 , n67898 , n67899 );
xor ( n67901 , n67898 , n67899 );
xor ( n67902 , n66719 , n67016 );
nor ( n67903 , n22231 , n67747 );
and ( n67904 , n67902 , n67903 );
xor ( n67905 , n67902 , n67903 );
xor ( n67906 , n66723 , n67014 );
nor ( n67907 , n21258 , n67747 );
and ( n67908 , n67906 , n67907 );
xor ( n67909 , n67906 , n67907 );
xor ( n67910 , n66727 , n67012 );
nor ( n67911 , n20303 , n67747 );
and ( n67912 , n67910 , n67911 );
xor ( n67913 , n67910 , n67911 );
xor ( n67914 , n66731 , n67010 );
nor ( n67915 , n19365 , n67747 );
and ( n67916 , n67914 , n67915 );
xor ( n67917 , n67914 , n67915 );
xor ( n67918 , n66735 , n67008 );
nor ( n67919 , n18448 , n67747 );
and ( n67920 , n67918 , n67919 );
xor ( n67921 , n67918 , n67919 );
xor ( n67922 , n66739 , n67006 );
nor ( n67923 , n17548 , n67747 );
and ( n67924 , n67922 , n67923 );
xor ( n67925 , n67922 , n67923 );
xor ( n67926 , n66743 , n67004 );
nor ( n67927 , n16669 , n67747 );
and ( n67928 , n67926 , n67927 );
xor ( n67929 , n67926 , n67927 );
xor ( n67930 , n66747 , n67002 );
nor ( n67931 , n15809 , n67747 );
and ( n67932 , n67930 , n67931 );
xor ( n67933 , n67930 , n67931 );
xor ( n67934 , n66751 , n67000 );
nor ( n67935 , n14968 , n67747 );
and ( n67936 , n67934 , n67935 );
xor ( n67937 , n67934 , n67935 );
xor ( n67938 , n66755 , n66998 );
nor ( n67939 , n14147 , n67747 );
and ( n67940 , n67938 , n67939 );
xor ( n67941 , n67938 , n67939 );
xor ( n67942 , n66759 , n66996 );
nor ( n67943 , n13349 , n67747 );
and ( n67944 , n67942 , n67943 );
xor ( n67945 , n67942 , n67943 );
xor ( n67946 , n66763 , n66994 );
nor ( n67947 , n12564 , n67747 );
and ( n67948 , n67946 , n67947 );
xor ( n67949 , n67946 , n67947 );
xor ( n67950 , n66767 , n66992 );
nor ( n67951 , n11799 , n67747 );
and ( n67952 , n67950 , n67951 );
xor ( n67953 , n67950 , n67951 );
xor ( n67954 , n66771 , n66990 );
nor ( n67955 , n11050 , n67747 );
and ( n67956 , n67954 , n67955 );
xor ( n67957 , n67954 , n67955 );
xor ( n67958 , n66775 , n66988 );
nor ( n67959 , n10321 , n67747 );
and ( n67960 , n67958 , n67959 );
xor ( n67961 , n67958 , n67959 );
xor ( n67962 , n66779 , n66986 );
nor ( n67963 , n9429 , n67747 );
and ( n67964 , n67962 , n67963 );
xor ( n67965 , n67962 , n67963 );
xor ( n67966 , n66783 , n66984 );
nor ( n67967 , n8949 , n67747 );
and ( n67968 , n67966 , n67967 );
xor ( n67969 , n67966 , n67967 );
xor ( n67970 , n66787 , n66982 );
nor ( n67971 , n9437 , n67747 );
and ( n67972 , n67970 , n67971 );
xor ( n67973 , n67970 , n67971 );
xor ( n67974 , n66791 , n66980 );
nor ( n67975 , n9446 , n67747 );
and ( n67976 , n67974 , n67975 );
xor ( n67977 , n67974 , n67975 );
xor ( n67978 , n66795 , n66978 );
nor ( n67979 , n9455 , n67747 );
and ( n67980 , n67978 , n67979 );
xor ( n67981 , n67978 , n67979 );
xor ( n67982 , n66799 , n66976 );
nor ( n67983 , n9464 , n67747 );
and ( n67984 , n67982 , n67983 );
xor ( n67985 , n67982 , n67983 );
xor ( n67986 , n66803 , n66974 );
nor ( n67987 , n9473 , n67747 );
and ( n67988 , n67986 , n67987 );
xor ( n67989 , n67986 , n67987 );
xor ( n67990 , n66807 , n66972 );
nor ( n67991 , n9482 , n67747 );
and ( n67992 , n67990 , n67991 );
xor ( n67993 , n67990 , n67991 );
xor ( n67994 , n66811 , n66970 );
nor ( n67995 , n9491 , n67747 );
and ( n67996 , n67994 , n67995 );
xor ( n67997 , n67994 , n67995 );
xor ( n67998 , n66815 , n66968 );
nor ( n67999 , n9500 , n67747 );
and ( n68000 , n67998 , n67999 );
xor ( n68001 , n67998 , n67999 );
xor ( n68002 , n66819 , n66966 );
nor ( n68003 , n9509 , n67747 );
and ( n68004 , n68002 , n68003 );
xor ( n68005 , n68002 , n68003 );
xor ( n68006 , n66823 , n66964 );
nor ( n68007 , n9518 , n67747 );
and ( n68008 , n68006 , n68007 );
xor ( n68009 , n68006 , n68007 );
xor ( n68010 , n66827 , n66962 );
nor ( n68011 , n9527 , n67747 );
and ( n68012 , n68010 , n68011 );
xor ( n68013 , n68010 , n68011 );
xor ( n68014 , n66831 , n66960 );
nor ( n68015 , n9536 , n67747 );
and ( n68016 , n68014 , n68015 );
xor ( n68017 , n68014 , n68015 );
xor ( n68018 , n66835 , n66958 );
nor ( n68019 , n9545 , n67747 );
and ( n68020 , n68018 , n68019 );
xor ( n68021 , n68018 , n68019 );
xor ( n68022 , n66839 , n66956 );
nor ( n68023 , n9554 , n67747 );
and ( n68024 , n68022 , n68023 );
xor ( n68025 , n68022 , n68023 );
xor ( n68026 , n66843 , n66954 );
nor ( n68027 , n9563 , n67747 );
and ( n68028 , n68026 , n68027 );
xor ( n68029 , n68026 , n68027 );
xor ( n68030 , n66847 , n66952 );
nor ( n68031 , n9572 , n67747 );
and ( n68032 , n68030 , n68031 );
xor ( n68033 , n68030 , n68031 );
xor ( n68034 , n66851 , n66950 );
nor ( n68035 , n9581 , n67747 );
and ( n68036 , n68034 , n68035 );
xor ( n68037 , n68034 , n68035 );
xor ( n68038 , n66855 , n66948 );
nor ( n68039 , n9590 , n67747 );
and ( n68040 , n68038 , n68039 );
xor ( n68041 , n68038 , n68039 );
xor ( n68042 , n66859 , n66946 );
nor ( n68043 , n9599 , n67747 );
and ( n68044 , n68042 , n68043 );
xor ( n68045 , n68042 , n68043 );
xor ( n68046 , n66863 , n66944 );
nor ( n68047 , n9608 , n67747 );
and ( n68048 , n68046 , n68047 );
xor ( n68049 , n68046 , n68047 );
xor ( n68050 , n66867 , n66942 );
nor ( n68051 , n9617 , n67747 );
and ( n68052 , n68050 , n68051 );
xor ( n68053 , n68050 , n68051 );
xor ( n68054 , n66871 , n66940 );
nor ( n68055 , n9626 , n67747 );
and ( n68056 , n68054 , n68055 );
xor ( n68057 , n68054 , n68055 );
xor ( n68058 , n66875 , n66938 );
nor ( n68059 , n9635 , n67747 );
and ( n68060 , n68058 , n68059 );
xor ( n68061 , n68058 , n68059 );
xor ( n68062 , n66879 , n66936 );
nor ( n68063 , n9644 , n67747 );
and ( n68064 , n68062 , n68063 );
xor ( n68065 , n68062 , n68063 );
xor ( n68066 , n66883 , n66934 );
nor ( n68067 , n9653 , n67747 );
and ( n68068 , n68066 , n68067 );
xor ( n68069 , n68066 , n68067 );
xor ( n68070 , n66887 , n66932 );
nor ( n68071 , n9662 , n67747 );
and ( n68072 , n68070 , n68071 );
xor ( n68073 , n68070 , n68071 );
xor ( n68074 , n66891 , n66930 );
nor ( n68075 , n9671 , n67747 );
and ( n68076 , n68074 , n68075 );
xor ( n68077 , n68074 , n68075 );
xor ( n68078 , n66895 , n66928 );
nor ( n68079 , n9680 , n67747 );
and ( n68080 , n68078 , n68079 );
xor ( n68081 , n68078 , n68079 );
xor ( n68082 , n66899 , n66926 );
nor ( n68083 , n9689 , n67747 );
and ( n68084 , n68082 , n68083 );
xor ( n68085 , n68082 , n68083 );
xor ( n68086 , n66903 , n66924 );
nor ( n68087 , n9698 , n67747 );
and ( n68088 , n68086 , n68087 );
xor ( n68089 , n68086 , n68087 );
xor ( n68090 , n66907 , n66922 );
nor ( n68091 , n9707 , n67747 );
and ( n68092 , n68090 , n68091 );
xor ( n68093 , n68090 , n68091 );
xor ( n68094 , n66911 , n66920 );
nor ( n68095 , n9716 , n67747 );
and ( n68096 , n68094 , n68095 );
xor ( n68097 , n68094 , n68095 );
xor ( n68098 , n66915 , n66918 );
nor ( n68099 , n9725 , n67747 );
and ( n68100 , n68098 , n68099 );
xor ( n68101 , n68098 , n68099 );
xor ( n68102 , n66916 , n66917 );
nor ( n68103 , n9734 , n67747 );
and ( n68104 , n68102 , n68103 );
xor ( n68105 , n68102 , n68103 );
nor ( n68106 , n9752 , n66561 );
nor ( n68107 , n9743 , n67747 );
and ( n68108 , n68106 , n68107 );
and ( n68109 , n68105 , n68108 );
or ( n68110 , n68104 , n68109 );
and ( n68111 , n68101 , n68110 );
or ( n68112 , n68100 , n68111 );
and ( n68113 , n68097 , n68112 );
or ( n68114 , n68096 , n68113 );
and ( n68115 , n68093 , n68114 );
or ( n68116 , n68092 , n68115 );
and ( n68117 , n68089 , n68116 );
or ( n68118 , n68088 , n68117 );
and ( n68119 , n68085 , n68118 );
or ( n68120 , n68084 , n68119 );
and ( n68121 , n68081 , n68120 );
or ( n68122 , n68080 , n68121 );
and ( n68123 , n68077 , n68122 );
or ( n68124 , n68076 , n68123 );
and ( n68125 , n68073 , n68124 );
or ( n68126 , n68072 , n68125 );
and ( n68127 , n68069 , n68126 );
or ( n68128 , n68068 , n68127 );
and ( n68129 , n68065 , n68128 );
or ( n68130 , n68064 , n68129 );
and ( n68131 , n68061 , n68130 );
or ( n68132 , n68060 , n68131 );
and ( n68133 , n68057 , n68132 );
or ( n68134 , n68056 , n68133 );
and ( n68135 , n68053 , n68134 );
or ( n68136 , n68052 , n68135 );
and ( n68137 , n68049 , n68136 );
or ( n68138 , n68048 , n68137 );
and ( n68139 , n68045 , n68138 );
or ( n68140 , n68044 , n68139 );
and ( n68141 , n68041 , n68140 );
or ( n68142 , n68040 , n68141 );
and ( n68143 , n68037 , n68142 );
or ( n68144 , n68036 , n68143 );
and ( n68145 , n68033 , n68144 );
or ( n68146 , n68032 , n68145 );
and ( n68147 , n68029 , n68146 );
or ( n68148 , n68028 , n68147 );
and ( n68149 , n68025 , n68148 );
or ( n68150 , n68024 , n68149 );
and ( n68151 , n68021 , n68150 );
or ( n68152 , n68020 , n68151 );
and ( n68153 , n68017 , n68152 );
or ( n68154 , n68016 , n68153 );
and ( n68155 , n68013 , n68154 );
or ( n68156 , n68012 , n68155 );
and ( n68157 , n68009 , n68156 );
or ( n68158 , n68008 , n68157 );
and ( n68159 , n68005 , n68158 );
or ( n68160 , n68004 , n68159 );
and ( n68161 , n68001 , n68160 );
or ( n68162 , n68000 , n68161 );
and ( n68163 , n67997 , n68162 );
or ( n68164 , n67996 , n68163 );
and ( n68165 , n67993 , n68164 );
or ( n68166 , n67992 , n68165 );
and ( n68167 , n67989 , n68166 );
or ( n68168 , n67988 , n68167 );
and ( n68169 , n67985 , n68168 );
or ( n68170 , n67984 , n68169 );
and ( n68171 , n67981 , n68170 );
or ( n68172 , n67980 , n68171 );
and ( n68173 , n67977 , n68172 );
or ( n68174 , n67976 , n68173 );
and ( n68175 , n67973 , n68174 );
or ( n68176 , n67972 , n68175 );
and ( n68177 , n67969 , n68176 );
or ( n68178 , n67968 , n68177 );
and ( n68179 , n67965 , n68178 );
or ( n68180 , n67964 , n68179 );
and ( n68181 , n67961 , n68180 );
or ( n68182 , n67960 , n68181 );
and ( n68183 , n67957 , n68182 );
or ( n68184 , n67956 , n68183 );
and ( n68185 , n67953 , n68184 );
or ( n68186 , n67952 , n68185 );
and ( n68187 , n67949 , n68186 );
or ( n68188 , n67948 , n68187 );
and ( n68189 , n67945 , n68188 );
or ( n68190 , n67944 , n68189 );
and ( n68191 , n67941 , n68190 );
or ( n68192 , n67940 , n68191 );
and ( n68193 , n67937 , n68192 );
or ( n68194 , n67936 , n68193 );
and ( n68195 , n67933 , n68194 );
or ( n68196 , n67932 , n68195 );
and ( n68197 , n67929 , n68196 );
or ( n68198 , n67928 , n68197 );
and ( n68199 , n67925 , n68198 );
or ( n68200 , n67924 , n68199 );
and ( n68201 , n67921 , n68200 );
or ( n68202 , n67920 , n68201 );
and ( n68203 , n67917 , n68202 );
or ( n68204 , n67916 , n68203 );
and ( n68205 , n67913 , n68204 );
or ( n68206 , n67912 , n68205 );
and ( n68207 , n67909 , n68206 );
or ( n68208 , n67908 , n68207 );
and ( n68209 , n67905 , n68208 );
or ( n68210 , n67904 , n68209 );
and ( n68211 , n67901 , n68210 );
or ( n68212 , n67900 , n68211 );
and ( n68213 , n67897 , n68212 );
or ( n68214 , n67896 , n68213 );
and ( n68215 , n67893 , n68214 );
or ( n68216 , n67892 , n68215 );
and ( n68217 , n67889 , n68216 );
or ( n68218 , n67888 , n68217 );
and ( n68219 , n67885 , n68218 );
or ( n68220 , n67884 , n68219 );
and ( n68221 , n67881 , n68220 );
or ( n68222 , n67880 , n68221 );
and ( n68223 , n67877 , n68222 );
or ( n68224 , n67876 , n68223 );
and ( n68225 , n67873 , n68224 );
or ( n68226 , n67872 , n68225 );
and ( n68227 , n67869 , n68226 );
or ( n68228 , n67868 , n68227 );
and ( n68229 , n67865 , n68228 );
or ( n68230 , n67864 , n68229 );
and ( n68231 , n67861 , n68230 );
or ( n68232 , n67860 , n68231 );
and ( n68233 , n67857 , n68232 );
or ( n68234 , n67856 , n68233 );
and ( n68235 , n67853 , n68234 );
or ( n68236 , n67852 , n68235 );
and ( n68237 , n67849 , n68236 );
or ( n68238 , n67848 , n68237 );
and ( n68239 , n67845 , n68238 );
or ( n68240 , n67844 , n68239 );
and ( n68241 , n67841 , n68240 );
or ( n68242 , n67840 , n68241 );
and ( n68243 , n67837 , n68242 );
or ( n68244 , n67836 , n68243 );
and ( n68245 , n67833 , n68244 );
or ( n68246 , n67832 , n68245 );
and ( n68247 , n67829 , n68246 );
or ( n68248 , n67828 , n68247 );
and ( n68249 , n67825 , n68248 );
or ( n68250 , n67824 , n68249 );
and ( n68251 , n67821 , n68250 );
or ( n68252 , n67820 , n68251 );
and ( n68253 , n67817 , n68252 );
or ( n68254 , n67816 , n68253 );
and ( n68255 , n67813 , n68254 );
or ( n68256 , n67812 , n68255 );
and ( n68257 , n67809 , n68256 );
or ( n68258 , n67808 , n68257 );
and ( n68259 , n67805 , n68258 );
or ( n68260 , n67804 , n68259 );
and ( n68261 , n67801 , n68260 );
or ( n68262 , n67800 , n68261 );
and ( n68263 , n67797 , n68262 );
or ( n68264 , n67796 , n68263 );
and ( n68265 , n67793 , n68264 );
or ( n68266 , n67792 , n68265 );
and ( n68267 , n67789 , n68266 );
or ( n68268 , n67788 , n68267 );
and ( n68269 , n67785 , n68268 );
or ( n68270 , n67784 , n68269 );
and ( n68271 , n67781 , n68270 );
or ( n68272 , n67780 , n68271 );
and ( n68273 , n67777 , n68272 );
or ( n68274 , n67776 , n68273 );
and ( n68275 , n67773 , n68274 );
or ( n68276 , n67772 , n68275 );
and ( n68277 , n67769 , n68276 );
or ( n68278 , n67768 , n68277 );
and ( n68279 , n67765 , n68278 );
or ( n68280 , n67764 , n68279 );
and ( n68281 , n67761 , n68280 );
or ( n68282 , n67760 , n68281 );
and ( n68283 , n67757 , n68282 );
or ( n68284 , n67756 , n68283 );
and ( n68285 , n67753 , n68284 );
or ( n68286 , n67752 , n68285 );
xor ( n68287 , n67749 , n68286 );
and ( n68288 , n33403 , n5837 );
nor ( n68289 , n5838 , n68288 );
nor ( n68290 , n6212 , n32231 );
xor ( n68291 , n68289 , n68290 );
and ( n68292 , n67097 , n67098 );
and ( n68293 , n67099 , n67102 );
or ( n68294 , n68292 , n68293 );
xor ( n68295 , n68291 , n68294 );
nor ( n68296 , n6596 , n31083 );
xor ( n68297 , n68295 , n68296 );
and ( n68298 , n67103 , n67104 );
and ( n68299 , n67105 , n67108 );
or ( n68300 , n68298 , n68299 );
xor ( n68301 , n68297 , n68300 );
nor ( n68302 , n6997 , n29948 );
xor ( n68303 , n68301 , n68302 );
and ( n68304 , n67109 , n67110 );
and ( n68305 , n67111 , n67114 );
or ( n68306 , n68304 , n68305 );
xor ( n68307 , n68303 , n68306 );
nor ( n68308 , n7413 , n28833 );
xor ( n68309 , n68307 , n68308 );
and ( n68310 , n67115 , n67116 );
and ( n68311 , n67117 , n67120 );
or ( n68312 , n68310 , n68311 );
xor ( n68313 , n68309 , n68312 );
nor ( n68314 , n7841 , n27737 );
xor ( n68315 , n68313 , n68314 );
and ( n68316 , n67121 , n67122 );
and ( n68317 , n67123 , n67126 );
or ( n68318 , n68316 , n68317 );
xor ( n68319 , n68315 , n68318 );
nor ( n68320 , n8281 , n26660 );
xor ( n68321 , n68319 , n68320 );
and ( n68322 , n67127 , n67128 );
and ( n68323 , n67129 , n67132 );
or ( n68324 , n68322 , n68323 );
xor ( n68325 , n68321 , n68324 );
nor ( n68326 , n8737 , n25600 );
xor ( n68327 , n68325 , n68326 );
and ( n68328 , n67133 , n67134 );
and ( n68329 , n67135 , n67138 );
or ( n68330 , n68328 , n68329 );
xor ( n68331 , n68327 , n68330 );
nor ( n68332 , n9420 , n24564 );
xor ( n68333 , n68331 , n68332 );
and ( n68334 , n67139 , n67140 );
and ( n68335 , n67141 , n67144 );
or ( n68336 , n68334 , n68335 );
xor ( n68337 , n68333 , n68336 );
nor ( n68338 , n10312 , n23541 );
xor ( n68339 , n68337 , n68338 );
and ( n68340 , n67145 , n67146 );
and ( n68341 , n67147 , n67150 );
or ( n68342 , n68340 , n68341 );
xor ( n68343 , n68339 , n68342 );
nor ( n68344 , n11041 , n22541 );
xor ( n68345 , n68343 , n68344 );
and ( n68346 , n67151 , n67152 );
and ( n68347 , n67153 , n67156 );
or ( n68348 , n68346 , n68347 );
xor ( n68349 , n68345 , n68348 );
nor ( n68350 , n11790 , n21562 );
xor ( n68351 , n68349 , n68350 );
and ( n68352 , n67157 , n67158 );
and ( n68353 , n67159 , n67162 );
or ( n68354 , n68352 , n68353 );
xor ( n68355 , n68351 , n68354 );
nor ( n68356 , n12555 , n20601 );
xor ( n68357 , n68355 , n68356 );
and ( n68358 , n67163 , n67164 );
and ( n68359 , n67165 , n67168 );
or ( n68360 , n68358 , n68359 );
xor ( n68361 , n68357 , n68360 );
nor ( n68362 , n13340 , n19657 );
xor ( n68363 , n68361 , n68362 );
and ( n68364 , n67169 , n67170 );
and ( n68365 , n67171 , n67174 );
or ( n68366 , n68364 , n68365 );
xor ( n68367 , n68363 , n68366 );
nor ( n68368 , n14138 , n18734 );
xor ( n68369 , n68367 , n68368 );
and ( n68370 , n67175 , n67176 );
and ( n68371 , n67177 , n67180 );
or ( n68372 , n68370 , n68371 );
xor ( n68373 , n68369 , n68372 );
nor ( n68374 , n14959 , n17828 );
xor ( n68375 , n68373 , n68374 );
and ( n68376 , n67181 , n67182 );
and ( n68377 , n67183 , n67186 );
or ( n68378 , n68376 , n68377 );
xor ( n68379 , n68375 , n68378 );
nor ( n68380 , n15800 , n16943 );
xor ( n68381 , n68379 , n68380 );
and ( n68382 , n67187 , n67188 );
and ( n68383 , n67189 , n67192 );
or ( n68384 , n68382 , n68383 );
xor ( n68385 , n68381 , n68384 );
nor ( n68386 , n16660 , n16077 );
xor ( n68387 , n68385 , n68386 );
and ( n68388 , n67193 , n67194 );
and ( n68389 , n67195 , n67198 );
or ( n68390 , n68388 , n68389 );
xor ( n68391 , n68387 , n68390 );
nor ( n68392 , n17539 , n15230 );
xor ( n68393 , n68391 , n68392 );
and ( n68394 , n67199 , n67200 );
and ( n68395 , n67201 , n67204 );
or ( n68396 , n68394 , n68395 );
xor ( n68397 , n68393 , n68396 );
nor ( n68398 , n18439 , n14403 );
xor ( n68399 , n68397 , n68398 );
and ( n68400 , n67205 , n67206 );
and ( n68401 , n67207 , n67210 );
or ( n68402 , n68400 , n68401 );
xor ( n68403 , n68399 , n68402 );
nor ( n68404 , n19356 , n13599 );
xor ( n68405 , n68403 , n68404 );
and ( n68406 , n67211 , n67212 );
and ( n68407 , n67213 , n67216 );
or ( n68408 , n68406 , n68407 );
xor ( n68409 , n68405 , n68408 );
nor ( n68410 , n20294 , n12808 );
xor ( n68411 , n68409 , n68410 );
and ( n68412 , n67217 , n67218 );
and ( n68413 , n67219 , n67222 );
or ( n68414 , n68412 , n68413 );
xor ( n68415 , n68411 , n68414 );
nor ( n68416 , n21249 , n12037 );
xor ( n68417 , n68415 , n68416 );
and ( n68418 , n67223 , n67224 );
and ( n68419 , n67225 , n67228 );
or ( n68420 , n68418 , n68419 );
xor ( n68421 , n68417 , n68420 );
nor ( n68422 , n22222 , n11282 );
xor ( n68423 , n68421 , n68422 );
and ( n68424 , n67229 , n67230 );
and ( n68425 , n67231 , n67234 );
or ( n68426 , n68424 , n68425 );
xor ( n68427 , n68423 , n68426 );
nor ( n68428 , n23216 , n10547 );
xor ( n68429 , n68427 , n68428 );
and ( n68430 , n67235 , n67236 );
and ( n68431 , n67237 , n67240 );
or ( n68432 , n68430 , n68431 );
xor ( n68433 , n68429 , n68432 );
nor ( n68434 , n24233 , n9829 );
xor ( n68435 , n68433 , n68434 );
and ( n68436 , n67241 , n67242 );
and ( n68437 , n67243 , n67246 );
or ( n68438 , n68436 , n68437 );
xor ( n68439 , n68435 , n68438 );
nor ( n68440 , n25263 , n8955 );
xor ( n68441 , n68439 , n68440 );
and ( n68442 , n67247 , n67248 );
and ( n68443 , n67249 , n67252 );
or ( n68444 , n68442 , n68443 );
xor ( n68445 , n68441 , n68444 );
nor ( n68446 , n26317 , n603 );
xor ( n68447 , n68445 , n68446 );
and ( n68448 , n67253 , n67254 );
and ( n68449 , n67255 , n67258 );
or ( n68450 , n68448 , n68449 );
xor ( n68451 , n68447 , n68450 );
nor ( n68452 , n27388 , n652 );
xor ( n68453 , n68451 , n68452 );
and ( n68454 , n67259 , n67260 );
and ( n68455 , n67261 , n67264 );
or ( n68456 , n68454 , n68455 );
xor ( n68457 , n68453 , n68456 );
nor ( n68458 , n28478 , n624 );
xor ( n68459 , n68457 , n68458 );
and ( n68460 , n67265 , n67266 );
and ( n68461 , n67267 , n67270 );
or ( n68462 , n68460 , n68461 );
xor ( n68463 , n68459 , n68462 );
nor ( n68464 , n29587 , n648 );
xor ( n68465 , n68463 , n68464 );
and ( n68466 , n67271 , n67272 );
and ( n68467 , n67273 , n67276 );
or ( n68468 , n68466 , n68467 );
xor ( n68469 , n68465 , n68468 );
nor ( n68470 , n30716 , n686 );
xor ( n68471 , n68469 , n68470 );
and ( n68472 , n67277 , n67278 );
and ( n68473 , n67279 , n67282 );
or ( n68474 , n68472 , n68473 );
xor ( n68475 , n68471 , n68474 );
nor ( n68476 , n31858 , n735 );
xor ( n68477 , n68475 , n68476 );
and ( n68478 , n67283 , n67284 );
and ( n68479 , n67285 , n67288 );
or ( n68480 , n68478 , n68479 );
xor ( n68481 , n68477 , n68480 );
nor ( n68482 , n33024 , n798 );
xor ( n68483 , n68481 , n68482 );
and ( n68484 , n67289 , n67290 );
and ( n68485 , n67291 , n67294 );
or ( n68486 , n68484 , n68485 );
xor ( n68487 , n68483 , n68486 );
nor ( n68488 , n34215 , n870 );
xor ( n68489 , n68487 , n68488 );
and ( n68490 , n67295 , n67296 );
and ( n68491 , n67297 , n67300 );
or ( n68492 , n68490 , n68491 );
xor ( n68493 , n68489 , n68492 );
nor ( n68494 , n35410 , n960 );
xor ( n68495 , n68493 , n68494 );
and ( n68496 , n67301 , n67302 );
and ( n68497 , n67303 , n67306 );
or ( n68498 , n68496 , n68497 );
xor ( n68499 , n68495 , n68498 );
nor ( n68500 , n36611 , n1064 );
xor ( n68501 , n68499 , n68500 );
and ( n68502 , n67307 , n67308 );
and ( n68503 , n67309 , n67312 );
or ( n68504 , n68502 , n68503 );
xor ( n68505 , n68501 , n68504 );
nor ( n68506 , n37816 , n1178 );
xor ( n68507 , n68505 , n68506 );
and ( n68508 , n67313 , n67314 );
and ( n68509 , n67315 , n67318 );
or ( n68510 , n68508 , n68509 );
xor ( n68511 , n68507 , n68510 );
nor ( n68512 , n39018 , n1305 );
xor ( n68513 , n68511 , n68512 );
and ( n68514 , n67319 , n67320 );
and ( n68515 , n67321 , n67324 );
or ( n68516 , n68514 , n68515 );
xor ( n68517 , n68513 , n68516 );
nor ( n68518 , n40223 , n1447 );
xor ( n68519 , n68517 , n68518 );
and ( n68520 , n67325 , n67326 );
and ( n68521 , n67327 , n67330 );
or ( n68522 , n68520 , n68521 );
xor ( n68523 , n68519 , n68522 );
nor ( n68524 , n41428 , n1600 );
xor ( n68525 , n68523 , n68524 );
and ( n68526 , n67331 , n67332 );
and ( n68527 , n67333 , n67336 );
or ( n68528 , n68526 , n68527 );
xor ( n68529 , n68525 , n68528 );
nor ( n68530 , n42632 , n1768 );
xor ( n68531 , n68529 , n68530 );
and ( n68532 , n67337 , n67338 );
and ( n68533 , n67339 , n67342 );
or ( n68534 , n68532 , n68533 );
xor ( n68535 , n68531 , n68534 );
nor ( n68536 , n43834 , n1947 );
xor ( n68537 , n68535 , n68536 );
and ( n68538 , n67343 , n67344 );
and ( n68539 , n67345 , n67348 );
or ( n68540 , n68538 , n68539 );
xor ( n68541 , n68537 , n68540 );
nor ( n68542 , n45038 , n2139 );
xor ( n68543 , n68541 , n68542 );
and ( n68544 , n67349 , n67350 );
and ( n68545 , n67351 , n67354 );
or ( n68546 , n68544 , n68545 );
xor ( n68547 , n68543 , n68546 );
nor ( n68548 , n46239 , n2345 );
xor ( n68549 , n68547 , n68548 );
and ( n68550 , n67355 , n67356 );
and ( n68551 , n67357 , n67360 );
or ( n68552 , n68550 , n68551 );
xor ( n68553 , n68549 , n68552 );
nor ( n68554 , n47440 , n2568 );
xor ( n68555 , n68553 , n68554 );
and ( n68556 , n67361 , n67362 );
and ( n68557 , n67363 , n67366 );
or ( n68558 , n68556 , n68557 );
xor ( n68559 , n68555 , n68558 );
nor ( n68560 , n48641 , n2799 );
xor ( n68561 , n68559 , n68560 );
and ( n68562 , n67367 , n67368 );
and ( n68563 , n67369 , n67372 );
or ( n68564 , n68562 , n68563 );
xor ( n68565 , n68561 , n68564 );
nor ( n68566 , n49841 , n3045 );
xor ( n68567 , n68565 , n68566 );
and ( n68568 , n67373 , n67374 );
and ( n68569 , n67375 , n67378 );
or ( n68570 , n68568 , n68569 );
xor ( n68571 , n68567 , n68570 );
nor ( n68572 , n51040 , n3302 );
xor ( n68573 , n68571 , n68572 );
and ( n68574 , n67379 , n67380 );
and ( n68575 , n67381 , n67384 );
or ( n68576 , n68574 , n68575 );
xor ( n68577 , n68573 , n68576 );
nor ( n68578 , n52238 , n3572 );
xor ( n68579 , n68577 , n68578 );
and ( n68580 , n67385 , n67386 );
and ( n68581 , n67387 , n67390 );
or ( n68582 , n68580 , n68581 );
xor ( n68583 , n68579 , n68582 );
nor ( n68584 , n53432 , n3855 );
xor ( n68585 , n68583 , n68584 );
and ( n68586 , n67391 , n67392 );
and ( n68587 , n67393 , n67396 );
or ( n68588 , n68586 , n68587 );
xor ( n68589 , n68585 , n68588 );
nor ( n68590 , n54629 , n4153 );
xor ( n68591 , n68589 , n68590 );
and ( n68592 , n67397 , n67398 );
and ( n68593 , n67399 , n67402 );
or ( n68594 , n68592 , n68593 );
xor ( n68595 , n68591 , n68594 );
nor ( n68596 , n55826 , n4460 );
xor ( n68597 , n68595 , n68596 );
and ( n68598 , n67403 , n67404 );
and ( n68599 , n67405 , n67408 );
or ( n68600 , n68598 , n68599 );
xor ( n68601 , n68597 , n68600 );
nor ( n68602 , n57022 , n4788 );
xor ( n68603 , n68601 , n68602 );
and ( n68604 , n67409 , n67410 );
and ( n68605 , n67411 , n67414 );
or ( n68606 , n68604 , n68605 );
xor ( n68607 , n68603 , n68606 );
nor ( n68608 , n58217 , n5128 );
xor ( n68609 , n68607 , n68608 );
and ( n68610 , n67415 , n67416 );
and ( n68611 , n67417 , n67420 );
or ( n68612 , n68610 , n68611 );
xor ( n68613 , n68609 , n68612 );
nor ( n68614 , n59412 , n5479 );
xor ( n68615 , n68613 , n68614 );
and ( n68616 , n67421 , n67422 );
and ( n68617 , n67423 , n67426 );
or ( n68618 , n68616 , n68617 );
xor ( n68619 , n68615 , n68618 );
nor ( n68620 , n60600 , n5840 );
xor ( n68621 , n68619 , n68620 );
and ( n68622 , n67427 , n67428 );
and ( n68623 , n67429 , n67432 );
or ( n68624 , n68622 , n68623 );
xor ( n68625 , n68621 , n68624 );
nor ( n68626 , n61791 , n6214 );
xor ( n68627 , n68625 , n68626 );
and ( n68628 , n67433 , n67434 );
and ( n68629 , n67435 , n67438 );
or ( n68630 , n68628 , n68629 );
xor ( n68631 , n68627 , n68630 );
nor ( n68632 , n62982 , n6598 );
xor ( n68633 , n68631 , n68632 );
and ( n68634 , n67439 , n67440 );
and ( n68635 , n67441 , n67444 );
or ( n68636 , n68634 , n68635 );
xor ( n68637 , n68633 , n68636 );
nor ( n68638 , n64172 , n6999 );
xor ( n68639 , n68637 , n68638 );
and ( n68640 , n67445 , n67446 );
and ( n68641 , n67447 , n67450 );
or ( n68642 , n68640 , n68641 );
xor ( n68643 , n68639 , n68642 );
nor ( n68644 , n65360 , n7415 );
xor ( n68645 , n68643 , n68644 );
and ( n68646 , n67451 , n67452 );
and ( n68647 , n67453 , n67456 );
or ( n68648 , n68646 , n68647 );
xor ( n68649 , n68645 , n68648 );
nor ( n68650 , n66550 , n7843 );
xor ( n68651 , n68649 , n68650 );
and ( n68652 , n67457 , n67458 );
and ( n68653 , n67459 , n67462 );
or ( n68654 , n68652 , n68653 );
xor ( n68655 , n68651 , n68654 );
nor ( n68656 , n67736 , n8283 );
xor ( n68657 , n68655 , n68656 );
and ( n68658 , n67463 , n67464 );
and ( n68659 , n67465 , n67468 );
or ( n68660 , n68658 , n68659 );
xor ( n68661 , n68657 , n68660 );
and ( n68662 , n67481 , n67485 );
and ( n68663 , n67485 , n67722 );
and ( n68664 , n67481 , n67722 );
or ( n68665 , n68662 , n68663 , n68664 );
and ( n68666 , n33774 , n5765 );
not ( n68667 , n5765 );
nor ( n68668 , n68666 , n68667 );
xor ( n68669 , n68665 , n68668 );
and ( n68670 , n67491 , n67495 );
and ( n68671 , n67495 , n67563 );
and ( n68672 , n67491 , n67563 );
or ( n68673 , n68670 , n68671 , n68672 );
and ( n68674 , n67487 , n67564 );
and ( n68675 , n67564 , n67721 );
and ( n68676 , n67487 , n67721 );
or ( n68677 , n68674 , n68675 , n68676 );
xor ( n68678 , n68673 , n68677 );
and ( n68679 , n67679 , n67720 );
and ( n68680 , n67569 , n67570 );
and ( n68681 , n67570 , n67678 );
and ( n68682 , n67569 , n67678 );
or ( n68683 , n68680 , n68681 , n68682 );
and ( n68684 , n67500 , n67504 );
and ( n68685 , n67504 , n67562 );
and ( n68686 , n67500 , n67562 );
or ( n68687 , n68684 , n68685 , n68686 );
xor ( n68688 , n68683 , n68687 );
and ( n68689 , n67531 , n67535 );
and ( n68690 , n67535 , n67541 );
and ( n68691 , n67531 , n67541 );
or ( n68692 , n68689 , n68690 , n68691 );
and ( n68693 , n67509 , n67513 );
and ( n68694 , n67513 , n67561 );
and ( n68695 , n67509 , n67561 );
or ( n68696 , n68693 , n68694 , n68695 );
xor ( n68697 , n68692 , n68696 );
and ( n68698 , n67518 , n67522 );
and ( n68699 , n67522 , n67560 );
and ( n68700 , n67518 , n67560 );
or ( n68701 , n68698 , n68699 , n68700 );
and ( n68702 , n67579 , n67604 );
and ( n68703 , n67604 , n67639 );
and ( n68704 , n67579 , n67639 );
or ( n68705 , n68702 , n68703 , n68704 );
xor ( n68706 , n68701 , n68705 );
and ( n68707 , n67527 , n67542 );
and ( n68708 , n67542 , n67559 );
and ( n68709 , n67527 , n67559 );
or ( n68710 , n68707 , n68708 , n68709 );
and ( n68711 , n67583 , n67587 );
and ( n68712 , n67587 , n67603 );
and ( n68713 , n67583 , n67603 );
or ( n68714 , n68711 , n68712 , n68713 );
xor ( n68715 , n68710 , n68714 );
and ( n68716 , n67547 , n67552 );
and ( n68717 , n67552 , n67558 );
and ( n68718 , n67547 , n67558 );
or ( n68719 , n68716 , n68717 , n68718 );
and ( n68720 , n67537 , n67538 );
and ( n68721 , n67538 , n67540 );
and ( n68722 , n67537 , n67540 );
or ( n68723 , n68720 , n68721 , n68722 );
and ( n68724 , n67548 , n67549 );
and ( n68725 , n67549 , n67551 );
and ( n68726 , n67548 , n67551 );
or ( n68727 , n68724 , n68725 , n68726 );
xor ( n68728 , n68723 , n68727 );
and ( n68729 , n30695 , n6971 );
and ( n68730 , n31836 , n6504 );
xor ( n68731 , n68729 , n68730 );
and ( n68732 , n32649 , n6132 );
xor ( n68733 , n68731 , n68732 );
xor ( n68734 , n68728 , n68733 );
xor ( n68735 , n68719 , n68734 );
and ( n68736 , n67554 , n67555 );
and ( n68737 , n67555 , n67557 );
and ( n68738 , n67554 , n67557 );
or ( n68739 , n68736 , n68737 , n68738 );
and ( n68740 , n27361 , n8243 );
and ( n68741 , n28456 , n7662 );
xor ( n68742 , n68740 , n68741 );
and ( n68743 , n29559 , n7310 );
xor ( n68744 , n68742 , n68743 );
xor ( n68745 , n68739 , n68744 );
and ( n68746 , n24214 , n10239 );
and ( n68747 , n25243 , n9348 );
xor ( n68748 , n68746 , n68747 );
and ( n68749 , n26296 , n8669 );
xor ( n68750 , n68748 , n68749 );
xor ( n68751 , n68745 , n68750 );
xor ( n68752 , n68735 , n68751 );
xor ( n68753 , n68715 , n68752 );
xor ( n68754 , n68706 , n68753 );
xor ( n68755 , n68697 , n68754 );
xor ( n68756 , n68688 , n68755 );
xor ( n68757 , n68679 , n68756 );
and ( n68758 , n67706 , n67711 );
and ( n68759 , n67711 , n67717 );
and ( n68760 , n67706 , n67717 );
or ( n68761 , n68758 , n68759 , n68760 );
and ( n68762 , n67696 , n67697 );
and ( n68763 , n67697 , n67699 );
and ( n68764 , n67696 , n67699 );
or ( n68765 , n68762 , n68763 , n68764 );
and ( n68766 , n67707 , n67708 );
and ( n68767 , n67708 , n67710 );
and ( n68768 , n67707 , n67710 );
or ( n68769 , n68766 , n68767 , n68768 );
xor ( n68770 , n68765 , n68769 );
and ( n68771 , n7385 , n29508 );
and ( n68772 , n7808 , n28406 );
xor ( n68773 , n68771 , n68772 );
and ( n68774 , n8079 , n27296 );
xor ( n68775 , n68773 , n68774 );
xor ( n68776 , n68770 , n68775 );
xor ( n68777 , n68761 , n68776 );
and ( n68778 , n67715 , n67716 );
not ( n68779 , n5819 );
and ( n68780 , n34193 , n5819 );
nor ( n68781 , n68779 , n68780 );
xor ( n68782 , n68778 , n68781 );
and ( n68783 , n6187 , n32999 );
and ( n68784 , n6569 , n31761 );
xor ( n68785 , n68783 , n68784 );
and ( n68786 , n6816 , n30629 );
xor ( n68787 , n68785 , n68786 );
xor ( n68788 , n68782 , n68787 );
xor ( n68789 , n68777 , n68788 );
and ( n68790 , n67575 , n67640 );
and ( n68791 , n67640 , n67677 );
and ( n68792 , n67575 , n67677 );
or ( n68793 , n68790 , n68791 , n68792 );
and ( n68794 , n67682 , n67719 );
xor ( n68795 , n68793 , n68794 );
and ( n68796 , n67645 , n67649 );
and ( n68797 , n67649 , n67676 );
and ( n68798 , n67645 , n67676 );
or ( n68799 , n68796 , n68797 , n68798 );
and ( n68800 , n67609 , n67622 );
and ( n68801 , n67622 , n67638 );
and ( n68802 , n67609 , n67638 );
or ( n68803 , n68800 , n68801 , n68802 );
and ( n68804 , n67592 , n67596 );
and ( n68805 , n67596 , n67602 );
and ( n68806 , n67592 , n67602 );
or ( n68807 , n68804 , n68805 , n68806 );
and ( n68808 , n67613 , n67618 );
and ( n68809 , n67618 , n67621 );
and ( n68810 , n67613 , n67621 );
or ( n68811 , n68808 , n68809 , n68810 );
xor ( n68812 , n68807 , n68811 );
and ( n68813 , n67598 , n67599 );
and ( n68814 , n67599 , n67601 );
and ( n68815 , n67598 , n67601 );
or ( n68816 , n68813 , n68814 , n68815 );
and ( n68817 , n67614 , n67615 );
and ( n68818 , n67615 , n67617 );
and ( n68819 , n67614 , n67617 );
or ( n68820 , n68817 , n68818 , n68819 );
xor ( n68821 , n68816 , n68820 );
and ( n68822 , n21216 , n12531 );
and ( n68823 , n22186 , n11718 );
xor ( n68824 , n68822 , n68823 );
and ( n68825 , n22892 , n10977 );
xor ( n68826 , n68824 , n68825 );
xor ( n68827 , n68821 , n68826 );
xor ( n68828 , n68812 , n68827 );
xor ( n68829 , n68803 , n68828 );
and ( n68830 , n67627 , n67631 );
and ( n68831 , n67631 , n67637 );
and ( n68832 , n67627 , n67637 );
or ( n68833 , n68830 , n68831 , n68832 );
and ( n68834 , n15758 , n16550 );
and ( n68835 , n16637 , n15691 );
and ( n68836 , n68834 , n68835 );
and ( n68837 , n68835 , n67620 );
and ( n68838 , n68834 , n67620 );
or ( n68839 , n68836 , n68837 , n68838 );
and ( n68840 , n18144 , n14838 );
and ( n68841 , n19324 , n14044 );
xor ( n68842 , n68840 , n68841 );
and ( n68843 , n20233 , n13256 );
xor ( n68844 , n68842 , n68843 );
xor ( n68845 , n68839 , n68844 );
and ( n68846 , n15758 , n17422 );
buf ( n68847 , n16637 );
xor ( n68848 , n68846 , n68847 );
and ( n68849 , n17512 , n15691 );
xor ( n68850 , n68848 , n68849 );
xor ( n68851 , n68845 , n68850 );
xor ( n68852 , n68833 , n68851 );
and ( n68853 , n67633 , n67634 );
and ( n68854 , n67634 , n67636 );
and ( n68855 , n67633 , n67636 );
or ( n68856 , n68853 , n68854 , n68855 );
and ( n68857 , n67664 , n67665 );
and ( n68858 , n67665 , n67667 );
and ( n68859 , n67664 , n67667 );
or ( n68860 , n68857 , n68858 , n68859 );
xor ( n68861 , n68856 , n68860 );
and ( n68862 , n13322 , n20156 );
and ( n68863 , n14118 , n19222 );
xor ( n68864 , n68862 , n68863 );
and ( n68865 , n14938 , n18407 );
xor ( n68866 , n68864 , n68865 );
xor ( n68867 , n68861 , n68866 );
xor ( n68868 , n68852 , n68867 );
xor ( n68869 , n68829 , n68868 );
xor ( n68870 , n68799 , n68869 );
and ( n68871 , n67654 , n67658 );
and ( n68872 , n67658 , n67675 );
and ( n68873 , n67654 , n67675 );
or ( n68874 , n68871 , n68872 , n68873 );
and ( n68875 , n67686 , n67701 );
and ( n68876 , n67701 , n67718 );
and ( n68877 , n67686 , n67718 );
or ( n68878 , n68875 , n68876 , n68877 );
xor ( n68879 , n68874 , n68878 );
and ( n68880 , n67663 , n67668 );
and ( n68881 , n67668 , n67674 );
and ( n68882 , n67663 , n67674 );
or ( n68883 , n68880 , n68881 , n68882 );
and ( n68884 , n67690 , n67694 );
and ( n68885 , n67694 , n67700 );
and ( n68886 , n67690 , n67700 );
or ( n68887 , n68884 , n68885 , n68886 );
xor ( n68888 , n68883 , n68887 );
and ( n68889 , n67670 , n67671 );
and ( n68890 , n67671 , n67673 );
and ( n68891 , n67670 , n67673 );
or ( n68892 , n68889 , n68890 , n68891 );
and ( n68893 , n11015 , n23075 );
and ( n68894 , n11769 , n22065 );
xor ( n68895 , n68893 , n68894 );
and ( n68896 , n12320 , n20976 );
xor ( n68897 , n68895 , n68896 );
xor ( n68898 , n68892 , n68897 );
and ( n68899 , n8718 , n26216 );
and ( n68900 , n9400 , n25163 );
xor ( n68901 , n68899 , n68900 );
and ( n68902 , n10291 , n24137 );
xor ( n68903 , n68901 , n68902 );
xor ( n68904 , n68898 , n68903 );
xor ( n68905 , n68888 , n68904 );
xor ( n68906 , n68879 , n68905 );
xor ( n68907 , n68870 , n68906 );
xor ( n68908 , n68795 , n68907 );
xor ( n68909 , n68789 , n68908 );
xor ( n68910 , n68757 , n68909 );
xor ( n68911 , n68678 , n68910 );
xor ( n68912 , n68669 , n68911 );
and ( n68913 , n67473 , n67476 );
and ( n68914 , n67476 , n67723 );
and ( n68915 , n67473 , n67723 );
or ( n68916 , n68913 , n68914 , n68915 );
xor ( n68917 , n68912 , n68916 );
and ( n68918 , n67724 , n67728 );
and ( n68919 , n67729 , n67732 );
or ( n68920 , n68918 , n68919 );
xor ( n68921 , n68917 , n68920 );
buf ( n68922 , n68921 );
buf ( n68923 , n68922 );
not ( n68924 , n68923 );
nor ( n68925 , n68924 , n8739 );
xor ( n68926 , n68661 , n68925 );
and ( n68927 , n67469 , n67737 );
and ( n68928 , n67738 , n67741 );
or ( n68929 , n68927 , n68928 );
xor ( n68930 , n68926 , n68929 );
buf ( n68931 , n68930 );
buf ( n68932 , n68931 );
not ( n68933 , n68932 );
buf ( n68934 , n591 );
not ( n68935 , n68934 );
nor ( n68936 , n68933 , n68935 );
xor ( n68937 , n68287 , n68936 );
xor ( n68938 , n67753 , n68284 );
nor ( n68939 , n67745 , n68935 );
and ( n68940 , n68938 , n68939 );
xor ( n68941 , n68938 , n68939 );
xor ( n68942 , n67757 , n68282 );
nor ( n68943 , n66559 , n68935 );
and ( n68944 , n68942 , n68943 );
xor ( n68945 , n68942 , n68943 );
xor ( n68946 , n67761 , n68280 );
nor ( n68947 , n65369 , n68935 );
and ( n68948 , n68946 , n68947 );
xor ( n68949 , n68946 , n68947 );
xor ( n68950 , n67765 , n68278 );
nor ( n68951 , n64181 , n68935 );
and ( n68952 , n68950 , n68951 );
xor ( n68953 , n68950 , n68951 );
xor ( n68954 , n67769 , n68276 );
nor ( n68955 , n62991 , n68935 );
and ( n68956 , n68954 , n68955 );
xor ( n68957 , n68954 , n68955 );
xor ( n68958 , n67773 , n68274 );
nor ( n68959 , n61800 , n68935 );
and ( n68960 , n68958 , n68959 );
xor ( n68961 , n68958 , n68959 );
xor ( n68962 , n67777 , n68272 );
nor ( n68963 , n60609 , n68935 );
and ( n68964 , n68962 , n68963 );
xor ( n68965 , n68962 , n68963 );
xor ( n68966 , n67781 , n68270 );
nor ( n68967 , n59421 , n68935 );
and ( n68968 , n68966 , n68967 );
xor ( n68969 , n68966 , n68967 );
xor ( n68970 , n67785 , n68268 );
nor ( n68971 , n58226 , n68935 );
and ( n68972 , n68970 , n68971 );
xor ( n68973 , n68970 , n68971 );
xor ( n68974 , n67789 , n68266 );
nor ( n68975 , n57031 , n68935 );
and ( n68976 , n68974 , n68975 );
xor ( n68977 , n68974 , n68975 );
xor ( n68978 , n67793 , n68264 );
nor ( n68979 , n55835 , n68935 );
and ( n68980 , n68978 , n68979 );
xor ( n68981 , n68978 , n68979 );
xor ( n68982 , n67797 , n68262 );
nor ( n68983 , n54638 , n68935 );
and ( n68984 , n68982 , n68983 );
xor ( n68985 , n68982 , n68983 );
xor ( n68986 , n67801 , n68260 );
nor ( n68987 , n53441 , n68935 );
and ( n68988 , n68986 , n68987 );
xor ( n68989 , n68986 , n68987 );
xor ( n68990 , n67805 , n68258 );
nor ( n68991 , n52247 , n68935 );
and ( n68992 , n68990 , n68991 );
xor ( n68993 , n68990 , n68991 );
xor ( n68994 , n67809 , n68256 );
nor ( n68995 , n51049 , n68935 );
and ( n68996 , n68994 , n68995 );
xor ( n68997 , n68994 , n68995 );
xor ( n68998 , n67813 , n68254 );
nor ( n68999 , n49850 , n68935 );
and ( n69000 , n68998 , n68999 );
xor ( n69001 , n68998 , n68999 );
xor ( n69002 , n67817 , n68252 );
nor ( n69003 , n48650 , n68935 );
and ( n69004 , n69002 , n69003 );
xor ( n69005 , n69002 , n69003 );
xor ( n69006 , n67821 , n68250 );
nor ( n69007 , n47449 , n68935 );
and ( n69008 , n69006 , n69007 );
xor ( n69009 , n69006 , n69007 );
xor ( n69010 , n67825 , n68248 );
nor ( n69011 , n46248 , n68935 );
and ( n69012 , n69010 , n69011 );
xor ( n69013 , n69010 , n69011 );
xor ( n69014 , n67829 , n68246 );
nor ( n69015 , n45047 , n68935 );
and ( n69016 , n69014 , n69015 );
xor ( n69017 , n69014 , n69015 );
xor ( n69018 , n67833 , n68244 );
nor ( n69019 , n43843 , n68935 );
and ( n69020 , n69018 , n69019 );
xor ( n69021 , n69018 , n69019 );
xor ( n69022 , n67837 , n68242 );
nor ( n69023 , n42641 , n68935 );
and ( n69024 , n69022 , n69023 );
xor ( n69025 , n69022 , n69023 );
xor ( n69026 , n67841 , n68240 );
nor ( n69027 , n41437 , n68935 );
and ( n69028 , n69026 , n69027 );
xor ( n69029 , n69026 , n69027 );
xor ( n69030 , n67845 , n68238 );
nor ( n69031 , n40232 , n68935 );
and ( n69032 , n69030 , n69031 );
xor ( n69033 , n69030 , n69031 );
xor ( n69034 , n67849 , n68236 );
nor ( n69035 , n39027 , n68935 );
and ( n69036 , n69034 , n69035 );
xor ( n69037 , n69034 , n69035 );
xor ( n69038 , n67853 , n68234 );
nor ( n69039 , n37825 , n68935 );
and ( n69040 , n69038 , n69039 );
xor ( n69041 , n69038 , n69039 );
xor ( n69042 , n67857 , n68232 );
nor ( n69043 , n36620 , n68935 );
and ( n69044 , n69042 , n69043 );
xor ( n69045 , n69042 , n69043 );
xor ( n69046 , n67861 , n68230 );
nor ( n69047 , n35419 , n68935 );
and ( n69048 , n69046 , n69047 );
xor ( n69049 , n69046 , n69047 );
xor ( n69050 , n67865 , n68228 );
nor ( n69051 , n34224 , n68935 );
and ( n69052 , n69050 , n69051 );
xor ( n69053 , n69050 , n69051 );
xor ( n69054 , n67869 , n68226 );
nor ( n69055 , n33033 , n68935 );
and ( n69056 , n69054 , n69055 );
xor ( n69057 , n69054 , n69055 );
xor ( n69058 , n67873 , n68224 );
nor ( n69059 , n31867 , n68935 );
and ( n69060 , n69058 , n69059 );
xor ( n69061 , n69058 , n69059 );
xor ( n69062 , n67877 , n68222 );
nor ( n69063 , n30725 , n68935 );
and ( n69064 , n69062 , n69063 );
xor ( n69065 , n69062 , n69063 );
xor ( n69066 , n67881 , n68220 );
nor ( n69067 , n29596 , n68935 );
and ( n69068 , n69066 , n69067 );
xor ( n69069 , n69066 , n69067 );
xor ( n69070 , n67885 , n68218 );
nor ( n69071 , n28487 , n68935 );
and ( n69072 , n69070 , n69071 );
xor ( n69073 , n69070 , n69071 );
xor ( n69074 , n67889 , n68216 );
nor ( n69075 , n27397 , n68935 );
and ( n69076 , n69074 , n69075 );
xor ( n69077 , n69074 , n69075 );
xor ( n69078 , n67893 , n68214 );
nor ( n69079 , n26326 , n68935 );
and ( n69080 , n69078 , n69079 );
xor ( n69081 , n69078 , n69079 );
xor ( n69082 , n67897 , n68212 );
nor ( n69083 , n25272 , n68935 );
and ( n69084 , n69082 , n69083 );
xor ( n69085 , n69082 , n69083 );
xor ( n69086 , n67901 , n68210 );
nor ( n69087 , n24242 , n68935 );
and ( n69088 , n69086 , n69087 );
xor ( n69089 , n69086 , n69087 );
xor ( n69090 , n67905 , n68208 );
nor ( n69091 , n23225 , n68935 );
and ( n69092 , n69090 , n69091 );
xor ( n69093 , n69090 , n69091 );
xor ( n69094 , n67909 , n68206 );
nor ( n69095 , n22231 , n68935 );
and ( n69096 , n69094 , n69095 );
xor ( n69097 , n69094 , n69095 );
xor ( n69098 , n67913 , n68204 );
nor ( n69099 , n21258 , n68935 );
and ( n69100 , n69098 , n69099 );
xor ( n69101 , n69098 , n69099 );
xor ( n69102 , n67917 , n68202 );
nor ( n69103 , n20303 , n68935 );
and ( n69104 , n69102 , n69103 );
xor ( n69105 , n69102 , n69103 );
xor ( n69106 , n67921 , n68200 );
nor ( n69107 , n19365 , n68935 );
and ( n69108 , n69106 , n69107 );
xor ( n69109 , n69106 , n69107 );
xor ( n69110 , n67925 , n68198 );
nor ( n69111 , n18448 , n68935 );
and ( n69112 , n69110 , n69111 );
xor ( n69113 , n69110 , n69111 );
xor ( n69114 , n67929 , n68196 );
nor ( n69115 , n17548 , n68935 );
and ( n69116 , n69114 , n69115 );
xor ( n69117 , n69114 , n69115 );
xor ( n69118 , n67933 , n68194 );
nor ( n69119 , n16669 , n68935 );
and ( n69120 , n69118 , n69119 );
xor ( n69121 , n69118 , n69119 );
xor ( n69122 , n67937 , n68192 );
nor ( n69123 , n15809 , n68935 );
and ( n69124 , n69122 , n69123 );
xor ( n69125 , n69122 , n69123 );
xor ( n69126 , n67941 , n68190 );
nor ( n69127 , n14968 , n68935 );
and ( n69128 , n69126 , n69127 );
xor ( n69129 , n69126 , n69127 );
xor ( n69130 , n67945 , n68188 );
nor ( n69131 , n14147 , n68935 );
and ( n69132 , n69130 , n69131 );
xor ( n69133 , n69130 , n69131 );
xor ( n69134 , n67949 , n68186 );
nor ( n69135 , n13349 , n68935 );
and ( n69136 , n69134 , n69135 );
xor ( n69137 , n69134 , n69135 );
xor ( n69138 , n67953 , n68184 );
nor ( n69139 , n12564 , n68935 );
and ( n69140 , n69138 , n69139 );
xor ( n69141 , n69138 , n69139 );
xor ( n69142 , n67957 , n68182 );
nor ( n69143 , n11799 , n68935 );
and ( n69144 , n69142 , n69143 );
xor ( n69145 , n69142 , n69143 );
xor ( n69146 , n67961 , n68180 );
nor ( n69147 , n11050 , n68935 );
and ( n69148 , n69146 , n69147 );
xor ( n69149 , n69146 , n69147 );
xor ( n69150 , n67965 , n68178 );
nor ( n69151 , n10321 , n68935 );
and ( n69152 , n69150 , n69151 );
xor ( n69153 , n69150 , n69151 );
xor ( n69154 , n67969 , n68176 );
nor ( n69155 , n9429 , n68935 );
and ( n69156 , n69154 , n69155 );
xor ( n69157 , n69154 , n69155 );
xor ( n69158 , n67973 , n68174 );
nor ( n69159 , n8949 , n68935 );
and ( n69160 , n69158 , n69159 );
xor ( n69161 , n69158 , n69159 );
xor ( n69162 , n67977 , n68172 );
nor ( n69163 , n9437 , n68935 );
and ( n69164 , n69162 , n69163 );
xor ( n69165 , n69162 , n69163 );
xor ( n69166 , n67981 , n68170 );
nor ( n69167 , n9446 , n68935 );
and ( n69168 , n69166 , n69167 );
xor ( n69169 , n69166 , n69167 );
xor ( n69170 , n67985 , n68168 );
nor ( n69171 , n9455 , n68935 );
and ( n69172 , n69170 , n69171 );
xor ( n69173 , n69170 , n69171 );
xor ( n69174 , n67989 , n68166 );
nor ( n69175 , n9464 , n68935 );
and ( n69176 , n69174 , n69175 );
xor ( n69177 , n69174 , n69175 );
xor ( n69178 , n67993 , n68164 );
nor ( n69179 , n9473 , n68935 );
and ( n69180 , n69178 , n69179 );
xor ( n69181 , n69178 , n69179 );
xor ( n69182 , n67997 , n68162 );
nor ( n69183 , n9482 , n68935 );
and ( n69184 , n69182 , n69183 );
xor ( n69185 , n69182 , n69183 );
xor ( n69186 , n68001 , n68160 );
nor ( n69187 , n9491 , n68935 );
and ( n69188 , n69186 , n69187 );
xor ( n69189 , n69186 , n69187 );
xor ( n69190 , n68005 , n68158 );
nor ( n69191 , n9500 , n68935 );
and ( n69192 , n69190 , n69191 );
xor ( n69193 , n69190 , n69191 );
xor ( n69194 , n68009 , n68156 );
nor ( n69195 , n9509 , n68935 );
and ( n69196 , n69194 , n69195 );
xor ( n69197 , n69194 , n69195 );
xor ( n69198 , n68013 , n68154 );
nor ( n69199 , n9518 , n68935 );
and ( n69200 , n69198 , n69199 );
xor ( n69201 , n69198 , n69199 );
xor ( n69202 , n68017 , n68152 );
nor ( n69203 , n9527 , n68935 );
and ( n69204 , n69202 , n69203 );
xor ( n69205 , n69202 , n69203 );
xor ( n69206 , n68021 , n68150 );
nor ( n69207 , n9536 , n68935 );
and ( n69208 , n69206 , n69207 );
xor ( n69209 , n69206 , n69207 );
xor ( n69210 , n68025 , n68148 );
nor ( n69211 , n9545 , n68935 );
and ( n69212 , n69210 , n69211 );
xor ( n69213 , n69210 , n69211 );
xor ( n69214 , n68029 , n68146 );
nor ( n69215 , n9554 , n68935 );
and ( n69216 , n69214 , n69215 );
xor ( n69217 , n69214 , n69215 );
xor ( n69218 , n68033 , n68144 );
nor ( n69219 , n9563 , n68935 );
and ( n69220 , n69218 , n69219 );
xor ( n69221 , n69218 , n69219 );
xor ( n69222 , n68037 , n68142 );
nor ( n69223 , n9572 , n68935 );
and ( n69224 , n69222 , n69223 );
xor ( n69225 , n69222 , n69223 );
xor ( n69226 , n68041 , n68140 );
nor ( n69227 , n9581 , n68935 );
and ( n69228 , n69226 , n69227 );
xor ( n69229 , n69226 , n69227 );
xor ( n69230 , n68045 , n68138 );
nor ( n69231 , n9590 , n68935 );
and ( n69232 , n69230 , n69231 );
xor ( n69233 , n69230 , n69231 );
xor ( n69234 , n68049 , n68136 );
nor ( n69235 , n9599 , n68935 );
and ( n69236 , n69234 , n69235 );
xor ( n69237 , n69234 , n69235 );
xor ( n69238 , n68053 , n68134 );
nor ( n69239 , n9608 , n68935 );
and ( n69240 , n69238 , n69239 );
xor ( n69241 , n69238 , n69239 );
xor ( n69242 , n68057 , n68132 );
nor ( n69243 , n9617 , n68935 );
and ( n69244 , n69242 , n69243 );
xor ( n69245 , n69242 , n69243 );
xor ( n69246 , n68061 , n68130 );
nor ( n69247 , n9626 , n68935 );
and ( n69248 , n69246 , n69247 );
xor ( n69249 , n69246 , n69247 );
xor ( n69250 , n68065 , n68128 );
nor ( n69251 , n9635 , n68935 );
and ( n69252 , n69250 , n69251 );
xor ( n69253 , n69250 , n69251 );
xor ( n69254 , n68069 , n68126 );
nor ( n69255 , n9644 , n68935 );
and ( n69256 , n69254 , n69255 );
xor ( n69257 , n69254 , n69255 );
xor ( n69258 , n68073 , n68124 );
nor ( n69259 , n9653 , n68935 );
and ( n69260 , n69258 , n69259 );
xor ( n69261 , n69258 , n69259 );
xor ( n69262 , n68077 , n68122 );
nor ( n69263 , n9662 , n68935 );
and ( n69264 , n69262 , n69263 );
xor ( n69265 , n69262 , n69263 );
xor ( n69266 , n68081 , n68120 );
nor ( n69267 , n9671 , n68935 );
and ( n69268 , n69266 , n69267 );
xor ( n69269 , n69266 , n69267 );
xor ( n69270 , n68085 , n68118 );
nor ( n69271 , n9680 , n68935 );
and ( n69272 , n69270 , n69271 );
xor ( n69273 , n69270 , n69271 );
xor ( n69274 , n68089 , n68116 );
nor ( n69275 , n9689 , n68935 );
and ( n69276 , n69274 , n69275 );
xor ( n69277 , n69274 , n69275 );
xor ( n69278 , n68093 , n68114 );
nor ( n69279 , n9698 , n68935 );
and ( n69280 , n69278 , n69279 );
xor ( n69281 , n69278 , n69279 );
xor ( n69282 , n68097 , n68112 );
nor ( n69283 , n9707 , n68935 );
and ( n69284 , n69282 , n69283 );
xor ( n69285 , n69282 , n69283 );
xor ( n69286 , n68101 , n68110 );
nor ( n69287 , n9716 , n68935 );
and ( n69288 , n69286 , n69287 );
xor ( n69289 , n69286 , n69287 );
xor ( n69290 , n68105 , n68108 );
nor ( n69291 , n9725 , n68935 );
and ( n69292 , n69290 , n69291 );
xor ( n69293 , n69290 , n69291 );
xor ( n69294 , n68106 , n68107 );
nor ( n69295 , n9734 , n68935 );
and ( n69296 , n69294 , n69295 );
xor ( n69297 , n69294 , n69295 );
nor ( n69298 , n9752 , n67747 );
nor ( n69299 , n9743 , n68935 );
and ( n69300 , n69298 , n69299 );
and ( n69301 , n69297 , n69300 );
or ( n69302 , n69296 , n69301 );
and ( n69303 , n69293 , n69302 );
or ( n69304 , n69292 , n69303 );
and ( n69305 , n69289 , n69304 );
or ( n69306 , n69288 , n69305 );
and ( n69307 , n69285 , n69306 );
or ( n69308 , n69284 , n69307 );
and ( n69309 , n69281 , n69308 );
or ( n69310 , n69280 , n69309 );
and ( n69311 , n69277 , n69310 );
or ( n69312 , n69276 , n69311 );
and ( n69313 , n69273 , n69312 );
or ( n69314 , n69272 , n69313 );
and ( n69315 , n69269 , n69314 );
or ( n69316 , n69268 , n69315 );
and ( n69317 , n69265 , n69316 );
or ( n69318 , n69264 , n69317 );
and ( n69319 , n69261 , n69318 );
or ( n69320 , n69260 , n69319 );
and ( n69321 , n69257 , n69320 );
or ( n69322 , n69256 , n69321 );
and ( n69323 , n69253 , n69322 );
or ( n69324 , n69252 , n69323 );
and ( n69325 , n69249 , n69324 );
or ( n69326 , n69248 , n69325 );
and ( n69327 , n69245 , n69326 );
or ( n69328 , n69244 , n69327 );
and ( n69329 , n69241 , n69328 );
or ( n69330 , n69240 , n69329 );
and ( n69331 , n69237 , n69330 );
or ( n69332 , n69236 , n69331 );
and ( n69333 , n69233 , n69332 );
or ( n69334 , n69232 , n69333 );
and ( n69335 , n69229 , n69334 );
or ( n69336 , n69228 , n69335 );
and ( n69337 , n69225 , n69336 );
or ( n69338 , n69224 , n69337 );
and ( n69339 , n69221 , n69338 );
or ( n69340 , n69220 , n69339 );
and ( n69341 , n69217 , n69340 );
or ( n69342 , n69216 , n69341 );
and ( n69343 , n69213 , n69342 );
or ( n69344 , n69212 , n69343 );
and ( n69345 , n69209 , n69344 );
or ( n69346 , n69208 , n69345 );
and ( n69347 , n69205 , n69346 );
or ( n69348 , n69204 , n69347 );
and ( n69349 , n69201 , n69348 );
or ( n69350 , n69200 , n69349 );
and ( n69351 , n69197 , n69350 );
or ( n69352 , n69196 , n69351 );
and ( n69353 , n69193 , n69352 );
or ( n69354 , n69192 , n69353 );
and ( n69355 , n69189 , n69354 );
or ( n69356 , n69188 , n69355 );
and ( n69357 , n69185 , n69356 );
or ( n69358 , n69184 , n69357 );
and ( n69359 , n69181 , n69358 );
or ( n69360 , n69180 , n69359 );
and ( n69361 , n69177 , n69360 );
or ( n69362 , n69176 , n69361 );
and ( n69363 , n69173 , n69362 );
or ( n69364 , n69172 , n69363 );
and ( n69365 , n69169 , n69364 );
or ( n69366 , n69168 , n69365 );
and ( n69367 , n69165 , n69366 );
or ( n69368 , n69164 , n69367 );
and ( n69369 , n69161 , n69368 );
or ( n69370 , n69160 , n69369 );
and ( n69371 , n69157 , n69370 );
or ( n69372 , n69156 , n69371 );
and ( n69373 , n69153 , n69372 );
or ( n69374 , n69152 , n69373 );
and ( n69375 , n69149 , n69374 );
or ( n69376 , n69148 , n69375 );
and ( n69377 , n69145 , n69376 );
or ( n69378 , n69144 , n69377 );
and ( n69379 , n69141 , n69378 );
or ( n69380 , n69140 , n69379 );
and ( n69381 , n69137 , n69380 );
or ( n69382 , n69136 , n69381 );
and ( n69383 , n69133 , n69382 );
or ( n69384 , n69132 , n69383 );
and ( n69385 , n69129 , n69384 );
or ( n69386 , n69128 , n69385 );
and ( n69387 , n69125 , n69386 );
or ( n69388 , n69124 , n69387 );
and ( n69389 , n69121 , n69388 );
or ( n69390 , n69120 , n69389 );
and ( n69391 , n69117 , n69390 );
or ( n69392 , n69116 , n69391 );
and ( n69393 , n69113 , n69392 );
or ( n69394 , n69112 , n69393 );
and ( n69395 , n69109 , n69394 );
or ( n69396 , n69108 , n69395 );
and ( n69397 , n69105 , n69396 );
or ( n69398 , n69104 , n69397 );
and ( n69399 , n69101 , n69398 );
or ( n69400 , n69100 , n69399 );
and ( n69401 , n69097 , n69400 );
or ( n69402 , n69096 , n69401 );
and ( n69403 , n69093 , n69402 );
or ( n69404 , n69092 , n69403 );
and ( n69405 , n69089 , n69404 );
or ( n69406 , n69088 , n69405 );
and ( n69407 , n69085 , n69406 );
or ( n69408 , n69084 , n69407 );
and ( n69409 , n69081 , n69408 );
or ( n69410 , n69080 , n69409 );
and ( n69411 , n69077 , n69410 );
or ( n69412 , n69076 , n69411 );
and ( n69413 , n69073 , n69412 );
or ( n69414 , n69072 , n69413 );
and ( n69415 , n69069 , n69414 );
or ( n69416 , n69068 , n69415 );
and ( n69417 , n69065 , n69416 );
or ( n69418 , n69064 , n69417 );
and ( n69419 , n69061 , n69418 );
or ( n69420 , n69060 , n69419 );
and ( n69421 , n69057 , n69420 );
or ( n69422 , n69056 , n69421 );
and ( n69423 , n69053 , n69422 );
or ( n69424 , n69052 , n69423 );
and ( n69425 , n69049 , n69424 );
or ( n69426 , n69048 , n69425 );
and ( n69427 , n69045 , n69426 );
or ( n69428 , n69044 , n69427 );
and ( n69429 , n69041 , n69428 );
or ( n69430 , n69040 , n69429 );
and ( n69431 , n69037 , n69430 );
or ( n69432 , n69036 , n69431 );
and ( n69433 , n69033 , n69432 );
or ( n69434 , n69032 , n69433 );
and ( n69435 , n69029 , n69434 );
or ( n69436 , n69028 , n69435 );
and ( n69437 , n69025 , n69436 );
or ( n69438 , n69024 , n69437 );
and ( n69439 , n69021 , n69438 );
or ( n69440 , n69020 , n69439 );
and ( n69441 , n69017 , n69440 );
or ( n69442 , n69016 , n69441 );
and ( n69443 , n69013 , n69442 );
or ( n69444 , n69012 , n69443 );
and ( n69445 , n69009 , n69444 );
or ( n69446 , n69008 , n69445 );
and ( n69447 , n69005 , n69446 );
or ( n69448 , n69004 , n69447 );
and ( n69449 , n69001 , n69448 );
or ( n69450 , n69000 , n69449 );
and ( n69451 , n68997 , n69450 );
or ( n69452 , n68996 , n69451 );
and ( n69453 , n68993 , n69452 );
or ( n69454 , n68992 , n69453 );
and ( n69455 , n68989 , n69454 );
or ( n69456 , n68988 , n69455 );
and ( n69457 , n68985 , n69456 );
or ( n69458 , n68984 , n69457 );
and ( n69459 , n68981 , n69458 );
or ( n69460 , n68980 , n69459 );
and ( n69461 , n68977 , n69460 );
or ( n69462 , n68976 , n69461 );
and ( n69463 , n68973 , n69462 );
or ( n69464 , n68972 , n69463 );
and ( n69465 , n68969 , n69464 );
or ( n69466 , n68968 , n69465 );
and ( n69467 , n68965 , n69466 );
or ( n69468 , n68964 , n69467 );
and ( n69469 , n68961 , n69468 );
or ( n69470 , n68960 , n69469 );
and ( n69471 , n68957 , n69470 );
or ( n69472 , n68956 , n69471 );
and ( n69473 , n68953 , n69472 );
or ( n69474 , n68952 , n69473 );
and ( n69475 , n68949 , n69474 );
or ( n69476 , n68948 , n69475 );
and ( n69477 , n68945 , n69476 );
or ( n69478 , n68944 , n69477 );
and ( n69479 , n68941 , n69478 );
or ( n69480 , n68940 , n69479 );
xor ( n69481 , n68937 , n69480 );
and ( n69482 , n33403 , n6211 );
nor ( n69483 , n6212 , n69482 );
nor ( n69484 , n6596 , n32231 );
xor ( n69485 , n69483 , n69484 );
and ( n69486 , n68289 , n68290 );
and ( n69487 , n68291 , n68294 );
or ( n69488 , n69486 , n69487 );
xor ( n69489 , n69485 , n69488 );
nor ( n69490 , n6997 , n31083 );
xor ( n69491 , n69489 , n69490 );
and ( n69492 , n68295 , n68296 );
and ( n69493 , n68297 , n68300 );
or ( n69494 , n69492 , n69493 );
xor ( n69495 , n69491 , n69494 );
nor ( n69496 , n7413 , n29948 );
xor ( n69497 , n69495 , n69496 );
and ( n69498 , n68301 , n68302 );
and ( n69499 , n68303 , n68306 );
or ( n69500 , n69498 , n69499 );
xor ( n69501 , n69497 , n69500 );
nor ( n69502 , n7841 , n28833 );
xor ( n69503 , n69501 , n69502 );
and ( n69504 , n68307 , n68308 );
and ( n69505 , n68309 , n68312 );
or ( n69506 , n69504 , n69505 );
xor ( n69507 , n69503 , n69506 );
nor ( n69508 , n8281 , n27737 );
xor ( n69509 , n69507 , n69508 );
and ( n69510 , n68313 , n68314 );
and ( n69511 , n68315 , n68318 );
or ( n69512 , n69510 , n69511 );
xor ( n69513 , n69509 , n69512 );
nor ( n69514 , n8737 , n26660 );
xor ( n69515 , n69513 , n69514 );
and ( n69516 , n68319 , n68320 );
and ( n69517 , n68321 , n68324 );
or ( n69518 , n69516 , n69517 );
xor ( n69519 , n69515 , n69518 );
nor ( n69520 , n9420 , n25600 );
xor ( n69521 , n69519 , n69520 );
and ( n69522 , n68325 , n68326 );
and ( n69523 , n68327 , n68330 );
or ( n69524 , n69522 , n69523 );
xor ( n69525 , n69521 , n69524 );
nor ( n69526 , n10312 , n24564 );
xor ( n69527 , n69525 , n69526 );
and ( n69528 , n68331 , n68332 );
and ( n69529 , n68333 , n68336 );
or ( n69530 , n69528 , n69529 );
xor ( n69531 , n69527 , n69530 );
nor ( n69532 , n11041 , n23541 );
xor ( n69533 , n69531 , n69532 );
and ( n69534 , n68337 , n68338 );
and ( n69535 , n68339 , n68342 );
or ( n69536 , n69534 , n69535 );
xor ( n69537 , n69533 , n69536 );
nor ( n69538 , n11790 , n22541 );
xor ( n69539 , n69537 , n69538 );
and ( n69540 , n68343 , n68344 );
and ( n69541 , n68345 , n68348 );
or ( n69542 , n69540 , n69541 );
xor ( n69543 , n69539 , n69542 );
nor ( n69544 , n12555 , n21562 );
xor ( n69545 , n69543 , n69544 );
and ( n69546 , n68349 , n68350 );
and ( n69547 , n68351 , n68354 );
or ( n69548 , n69546 , n69547 );
xor ( n69549 , n69545 , n69548 );
nor ( n69550 , n13340 , n20601 );
xor ( n69551 , n69549 , n69550 );
and ( n69552 , n68355 , n68356 );
and ( n69553 , n68357 , n68360 );
or ( n69554 , n69552 , n69553 );
xor ( n69555 , n69551 , n69554 );
nor ( n69556 , n14138 , n19657 );
xor ( n69557 , n69555 , n69556 );
and ( n69558 , n68361 , n68362 );
and ( n69559 , n68363 , n68366 );
or ( n69560 , n69558 , n69559 );
xor ( n69561 , n69557 , n69560 );
nor ( n69562 , n14959 , n18734 );
xor ( n69563 , n69561 , n69562 );
and ( n69564 , n68367 , n68368 );
and ( n69565 , n68369 , n68372 );
or ( n69566 , n69564 , n69565 );
xor ( n69567 , n69563 , n69566 );
nor ( n69568 , n15800 , n17828 );
xor ( n69569 , n69567 , n69568 );
and ( n69570 , n68373 , n68374 );
and ( n69571 , n68375 , n68378 );
or ( n69572 , n69570 , n69571 );
xor ( n69573 , n69569 , n69572 );
nor ( n69574 , n16660 , n16943 );
xor ( n69575 , n69573 , n69574 );
and ( n69576 , n68379 , n68380 );
and ( n69577 , n68381 , n68384 );
or ( n69578 , n69576 , n69577 );
xor ( n69579 , n69575 , n69578 );
nor ( n69580 , n17539 , n16077 );
xor ( n69581 , n69579 , n69580 );
and ( n69582 , n68385 , n68386 );
and ( n69583 , n68387 , n68390 );
or ( n69584 , n69582 , n69583 );
xor ( n69585 , n69581 , n69584 );
nor ( n69586 , n18439 , n15230 );
xor ( n69587 , n69585 , n69586 );
and ( n69588 , n68391 , n68392 );
and ( n69589 , n68393 , n68396 );
or ( n69590 , n69588 , n69589 );
xor ( n69591 , n69587 , n69590 );
nor ( n69592 , n19356 , n14403 );
xor ( n69593 , n69591 , n69592 );
and ( n69594 , n68397 , n68398 );
and ( n69595 , n68399 , n68402 );
or ( n69596 , n69594 , n69595 );
xor ( n69597 , n69593 , n69596 );
nor ( n69598 , n20294 , n13599 );
xor ( n69599 , n69597 , n69598 );
and ( n69600 , n68403 , n68404 );
and ( n69601 , n68405 , n68408 );
or ( n69602 , n69600 , n69601 );
xor ( n69603 , n69599 , n69602 );
nor ( n69604 , n21249 , n12808 );
xor ( n69605 , n69603 , n69604 );
and ( n69606 , n68409 , n68410 );
and ( n69607 , n68411 , n68414 );
or ( n69608 , n69606 , n69607 );
xor ( n69609 , n69605 , n69608 );
nor ( n69610 , n22222 , n12037 );
xor ( n69611 , n69609 , n69610 );
and ( n69612 , n68415 , n68416 );
and ( n69613 , n68417 , n68420 );
or ( n69614 , n69612 , n69613 );
xor ( n69615 , n69611 , n69614 );
nor ( n69616 , n23216 , n11282 );
xor ( n69617 , n69615 , n69616 );
and ( n69618 , n68421 , n68422 );
and ( n69619 , n68423 , n68426 );
or ( n69620 , n69618 , n69619 );
xor ( n69621 , n69617 , n69620 );
nor ( n69622 , n24233 , n10547 );
xor ( n69623 , n69621 , n69622 );
and ( n69624 , n68427 , n68428 );
and ( n69625 , n68429 , n68432 );
or ( n69626 , n69624 , n69625 );
xor ( n69627 , n69623 , n69626 );
nor ( n69628 , n25263 , n9829 );
xor ( n69629 , n69627 , n69628 );
and ( n69630 , n68433 , n68434 );
and ( n69631 , n68435 , n68438 );
or ( n69632 , n69630 , n69631 );
xor ( n69633 , n69629 , n69632 );
nor ( n69634 , n26317 , n8955 );
xor ( n69635 , n69633 , n69634 );
and ( n69636 , n68439 , n68440 );
and ( n69637 , n68441 , n68444 );
or ( n69638 , n69636 , n69637 );
xor ( n69639 , n69635 , n69638 );
nor ( n69640 , n27388 , n603 );
xor ( n69641 , n69639 , n69640 );
and ( n69642 , n68445 , n68446 );
and ( n69643 , n68447 , n68450 );
or ( n69644 , n69642 , n69643 );
xor ( n69645 , n69641 , n69644 );
nor ( n69646 , n28478 , n652 );
xor ( n69647 , n69645 , n69646 );
and ( n69648 , n68451 , n68452 );
and ( n69649 , n68453 , n68456 );
or ( n69650 , n69648 , n69649 );
xor ( n69651 , n69647 , n69650 );
nor ( n69652 , n29587 , n624 );
xor ( n69653 , n69651 , n69652 );
and ( n69654 , n68457 , n68458 );
and ( n69655 , n68459 , n68462 );
or ( n69656 , n69654 , n69655 );
xor ( n69657 , n69653 , n69656 );
nor ( n69658 , n30716 , n648 );
xor ( n69659 , n69657 , n69658 );
and ( n69660 , n68463 , n68464 );
and ( n69661 , n68465 , n68468 );
or ( n69662 , n69660 , n69661 );
xor ( n69663 , n69659 , n69662 );
nor ( n69664 , n31858 , n686 );
xor ( n69665 , n69663 , n69664 );
and ( n69666 , n68469 , n68470 );
and ( n69667 , n68471 , n68474 );
or ( n69668 , n69666 , n69667 );
xor ( n69669 , n69665 , n69668 );
nor ( n69670 , n33024 , n735 );
xor ( n69671 , n69669 , n69670 );
and ( n69672 , n68475 , n68476 );
and ( n69673 , n68477 , n68480 );
or ( n69674 , n69672 , n69673 );
xor ( n69675 , n69671 , n69674 );
nor ( n69676 , n34215 , n798 );
xor ( n69677 , n69675 , n69676 );
and ( n69678 , n68481 , n68482 );
and ( n69679 , n68483 , n68486 );
or ( n69680 , n69678 , n69679 );
xor ( n69681 , n69677 , n69680 );
nor ( n69682 , n35410 , n870 );
xor ( n69683 , n69681 , n69682 );
and ( n69684 , n68487 , n68488 );
and ( n69685 , n68489 , n68492 );
or ( n69686 , n69684 , n69685 );
xor ( n69687 , n69683 , n69686 );
nor ( n69688 , n36611 , n960 );
xor ( n69689 , n69687 , n69688 );
and ( n69690 , n68493 , n68494 );
and ( n69691 , n68495 , n68498 );
or ( n69692 , n69690 , n69691 );
xor ( n69693 , n69689 , n69692 );
nor ( n69694 , n37816 , n1064 );
xor ( n69695 , n69693 , n69694 );
and ( n69696 , n68499 , n68500 );
and ( n69697 , n68501 , n68504 );
or ( n69698 , n69696 , n69697 );
xor ( n69699 , n69695 , n69698 );
nor ( n69700 , n39018 , n1178 );
xor ( n69701 , n69699 , n69700 );
and ( n69702 , n68505 , n68506 );
and ( n69703 , n68507 , n68510 );
or ( n69704 , n69702 , n69703 );
xor ( n69705 , n69701 , n69704 );
nor ( n69706 , n40223 , n1305 );
xor ( n69707 , n69705 , n69706 );
and ( n69708 , n68511 , n68512 );
and ( n69709 , n68513 , n68516 );
or ( n69710 , n69708 , n69709 );
xor ( n69711 , n69707 , n69710 );
nor ( n69712 , n41428 , n1447 );
xor ( n69713 , n69711 , n69712 );
and ( n69714 , n68517 , n68518 );
and ( n69715 , n68519 , n68522 );
or ( n69716 , n69714 , n69715 );
xor ( n69717 , n69713 , n69716 );
nor ( n69718 , n42632 , n1600 );
xor ( n69719 , n69717 , n69718 );
and ( n69720 , n68523 , n68524 );
and ( n69721 , n68525 , n68528 );
or ( n69722 , n69720 , n69721 );
xor ( n69723 , n69719 , n69722 );
nor ( n69724 , n43834 , n1768 );
xor ( n69725 , n69723 , n69724 );
and ( n69726 , n68529 , n68530 );
and ( n69727 , n68531 , n68534 );
or ( n69728 , n69726 , n69727 );
xor ( n69729 , n69725 , n69728 );
nor ( n69730 , n45038 , n1947 );
xor ( n69731 , n69729 , n69730 );
and ( n69732 , n68535 , n68536 );
and ( n69733 , n68537 , n68540 );
or ( n69734 , n69732 , n69733 );
xor ( n69735 , n69731 , n69734 );
nor ( n69736 , n46239 , n2139 );
xor ( n69737 , n69735 , n69736 );
and ( n69738 , n68541 , n68542 );
and ( n69739 , n68543 , n68546 );
or ( n69740 , n69738 , n69739 );
xor ( n69741 , n69737 , n69740 );
nor ( n69742 , n47440 , n2345 );
xor ( n69743 , n69741 , n69742 );
and ( n69744 , n68547 , n68548 );
and ( n69745 , n68549 , n68552 );
or ( n69746 , n69744 , n69745 );
xor ( n69747 , n69743 , n69746 );
nor ( n69748 , n48641 , n2568 );
xor ( n69749 , n69747 , n69748 );
and ( n69750 , n68553 , n68554 );
and ( n69751 , n68555 , n68558 );
or ( n69752 , n69750 , n69751 );
xor ( n69753 , n69749 , n69752 );
nor ( n69754 , n49841 , n2799 );
xor ( n69755 , n69753 , n69754 );
and ( n69756 , n68559 , n68560 );
and ( n69757 , n68561 , n68564 );
or ( n69758 , n69756 , n69757 );
xor ( n69759 , n69755 , n69758 );
nor ( n69760 , n51040 , n3045 );
xor ( n69761 , n69759 , n69760 );
and ( n69762 , n68565 , n68566 );
and ( n69763 , n68567 , n68570 );
or ( n69764 , n69762 , n69763 );
xor ( n69765 , n69761 , n69764 );
nor ( n69766 , n52238 , n3302 );
xor ( n69767 , n69765 , n69766 );
and ( n69768 , n68571 , n68572 );
and ( n69769 , n68573 , n68576 );
or ( n69770 , n69768 , n69769 );
xor ( n69771 , n69767 , n69770 );
nor ( n69772 , n53432 , n3572 );
xor ( n69773 , n69771 , n69772 );
and ( n69774 , n68577 , n68578 );
and ( n69775 , n68579 , n68582 );
or ( n69776 , n69774 , n69775 );
xor ( n69777 , n69773 , n69776 );
nor ( n69778 , n54629 , n3855 );
xor ( n69779 , n69777 , n69778 );
and ( n69780 , n68583 , n68584 );
and ( n69781 , n68585 , n68588 );
or ( n69782 , n69780 , n69781 );
xor ( n69783 , n69779 , n69782 );
nor ( n69784 , n55826 , n4153 );
xor ( n69785 , n69783 , n69784 );
and ( n69786 , n68589 , n68590 );
and ( n69787 , n68591 , n68594 );
or ( n69788 , n69786 , n69787 );
xor ( n69789 , n69785 , n69788 );
nor ( n69790 , n57022 , n4460 );
xor ( n69791 , n69789 , n69790 );
and ( n69792 , n68595 , n68596 );
and ( n69793 , n68597 , n68600 );
or ( n69794 , n69792 , n69793 );
xor ( n69795 , n69791 , n69794 );
nor ( n69796 , n58217 , n4788 );
xor ( n69797 , n69795 , n69796 );
and ( n69798 , n68601 , n68602 );
and ( n69799 , n68603 , n68606 );
or ( n69800 , n69798 , n69799 );
xor ( n69801 , n69797 , n69800 );
nor ( n69802 , n59412 , n5128 );
xor ( n69803 , n69801 , n69802 );
and ( n69804 , n68607 , n68608 );
and ( n69805 , n68609 , n68612 );
or ( n69806 , n69804 , n69805 );
xor ( n69807 , n69803 , n69806 );
nor ( n69808 , n60600 , n5479 );
xor ( n69809 , n69807 , n69808 );
and ( n69810 , n68613 , n68614 );
and ( n69811 , n68615 , n68618 );
or ( n69812 , n69810 , n69811 );
xor ( n69813 , n69809 , n69812 );
nor ( n69814 , n61791 , n5840 );
xor ( n69815 , n69813 , n69814 );
and ( n69816 , n68619 , n68620 );
and ( n69817 , n68621 , n68624 );
or ( n69818 , n69816 , n69817 );
xor ( n69819 , n69815 , n69818 );
nor ( n69820 , n62982 , n6214 );
xor ( n69821 , n69819 , n69820 );
and ( n69822 , n68625 , n68626 );
and ( n69823 , n68627 , n68630 );
or ( n69824 , n69822 , n69823 );
xor ( n69825 , n69821 , n69824 );
nor ( n69826 , n64172 , n6598 );
xor ( n69827 , n69825 , n69826 );
and ( n69828 , n68631 , n68632 );
and ( n69829 , n68633 , n68636 );
or ( n69830 , n69828 , n69829 );
xor ( n69831 , n69827 , n69830 );
nor ( n69832 , n65360 , n6999 );
xor ( n69833 , n69831 , n69832 );
and ( n69834 , n68637 , n68638 );
and ( n69835 , n68639 , n68642 );
or ( n69836 , n69834 , n69835 );
xor ( n69837 , n69833 , n69836 );
nor ( n69838 , n66550 , n7415 );
xor ( n69839 , n69837 , n69838 );
and ( n69840 , n68643 , n68644 );
and ( n69841 , n68645 , n68648 );
or ( n69842 , n69840 , n69841 );
xor ( n69843 , n69839 , n69842 );
nor ( n69844 , n67736 , n7843 );
xor ( n69845 , n69843 , n69844 );
and ( n69846 , n68649 , n68650 );
and ( n69847 , n68651 , n68654 );
or ( n69848 , n69846 , n69847 );
xor ( n69849 , n69845 , n69848 );
nor ( n69850 , n68924 , n8283 );
xor ( n69851 , n69849 , n69850 );
and ( n69852 , n68655 , n68656 );
and ( n69853 , n68657 , n68660 );
or ( n69854 , n69852 , n69853 );
xor ( n69855 , n69851 , n69854 );
and ( n69856 , n68673 , n68677 );
and ( n69857 , n68677 , n68910 );
and ( n69858 , n68673 , n68910 );
or ( n69859 , n69856 , n69857 , n69858 );
and ( n69860 , n33774 , n6132 );
not ( n69861 , n6132 );
nor ( n69862 , n69860 , n69861 );
xor ( n69863 , n69859 , n69862 );
and ( n69864 , n68683 , n68687 );
and ( n69865 , n68687 , n68755 );
and ( n69866 , n68683 , n68755 );
or ( n69867 , n69864 , n69865 , n69866 );
and ( n69868 , n68679 , n68756 );
and ( n69869 , n68756 , n68909 );
and ( n69870 , n68679 , n68909 );
or ( n69871 , n69868 , n69869 , n69870 );
xor ( n69872 , n69867 , n69871 );
and ( n69873 , n68789 , n68908 );
and ( n69874 , n68793 , n68794 );
and ( n69875 , n68794 , n68907 );
and ( n69876 , n68793 , n68907 );
or ( n69877 , n69874 , n69875 , n69876 );
and ( n69878 , n68692 , n68696 );
and ( n69879 , n68696 , n68754 );
and ( n69880 , n68692 , n68754 );
or ( n69881 , n69878 , n69879 , n69880 );
xor ( n69882 , n69877 , n69881 );
and ( n69883 , n68723 , n68727 );
and ( n69884 , n68727 , n68733 );
and ( n69885 , n68723 , n68733 );
or ( n69886 , n69883 , n69884 , n69885 );
and ( n69887 , n68701 , n68705 );
and ( n69888 , n68705 , n68753 );
and ( n69889 , n68701 , n68753 );
or ( n69890 , n69887 , n69888 , n69889 );
xor ( n69891 , n69886 , n69890 );
and ( n69892 , n68710 , n68714 );
and ( n69893 , n68714 , n68752 );
and ( n69894 , n68710 , n68752 );
or ( n69895 , n69892 , n69893 , n69894 );
and ( n69896 , n68803 , n68828 );
and ( n69897 , n68828 , n68868 );
and ( n69898 , n68803 , n68868 );
or ( n69899 , n69896 , n69897 , n69898 );
xor ( n69900 , n69895 , n69899 );
and ( n69901 , n68719 , n68734 );
and ( n69902 , n68734 , n68751 );
and ( n69903 , n68719 , n68751 );
or ( n69904 , n69901 , n69902 , n69903 );
and ( n69905 , n68807 , n68811 );
and ( n69906 , n68811 , n68827 );
and ( n69907 , n68807 , n68827 );
or ( n69908 , n69905 , n69906 , n69907 );
xor ( n69909 , n69904 , n69908 );
and ( n69910 , n68739 , n68744 );
and ( n69911 , n68744 , n68750 );
and ( n69912 , n68739 , n68750 );
or ( n69913 , n69910 , n69911 , n69912 );
and ( n69914 , n68729 , n68730 );
and ( n69915 , n68730 , n68732 );
and ( n69916 , n68729 , n68732 );
or ( n69917 , n69914 , n69915 , n69916 );
and ( n69918 , n68740 , n68741 );
and ( n69919 , n68741 , n68743 );
and ( n69920 , n68740 , n68743 );
or ( n69921 , n69918 , n69919 , n69920 );
xor ( n69922 , n69917 , n69921 );
and ( n69923 , n30695 , n7310 );
and ( n69924 , n31836 , n6971 );
xor ( n69925 , n69923 , n69924 );
and ( n69926 , n32649 , n6504 );
xor ( n69927 , n69925 , n69926 );
xor ( n69928 , n69922 , n69927 );
xor ( n69929 , n69913 , n69928 );
and ( n69930 , n68746 , n68747 );
and ( n69931 , n68747 , n68749 );
and ( n69932 , n68746 , n68749 );
or ( n69933 , n69930 , n69931 , n69932 );
and ( n69934 , n27361 , n8669 );
and ( n69935 , n28456 , n8243 );
xor ( n69936 , n69934 , n69935 );
and ( n69937 , n29559 , n7662 );
xor ( n69938 , n69936 , n69937 );
xor ( n69939 , n69933 , n69938 );
and ( n69940 , n24214 , n10977 );
and ( n69941 , n25243 , n10239 );
xor ( n69942 , n69940 , n69941 );
and ( n69943 , n26296 , n9348 );
xor ( n69944 , n69942 , n69943 );
xor ( n69945 , n69939 , n69944 );
xor ( n69946 , n69929 , n69945 );
xor ( n69947 , n69909 , n69946 );
xor ( n69948 , n69900 , n69947 );
xor ( n69949 , n69891 , n69948 );
xor ( n69950 , n69882 , n69949 );
xor ( n69951 , n69873 , n69950 );
and ( n69952 , n68778 , n68781 );
and ( n69953 , n68781 , n68787 );
and ( n69954 , n68778 , n68787 );
or ( n69955 , n69952 , n69953 , n69954 );
not ( n69956 , n6187 );
and ( n69957 , n34193 , n6187 );
nor ( n69958 , n69956 , n69957 );
and ( n69959 , n6569 , n32999 );
xor ( n69960 , n69958 , n69959 );
and ( n69961 , n6816 , n31761 );
xor ( n69962 , n69960 , n69961 );
xor ( n69963 , n69955 , n69962 );
and ( n69964 , n68771 , n68772 );
and ( n69965 , n68772 , n68774 );
and ( n69966 , n68771 , n68774 );
or ( n69967 , n69964 , n69965 , n69966 );
and ( n69968 , n68783 , n68784 );
and ( n69969 , n68784 , n68786 );
and ( n69970 , n68783 , n68786 );
or ( n69971 , n69968 , n69969 , n69970 );
xor ( n69972 , n69967 , n69971 );
and ( n69973 , n7385 , n30629 );
and ( n69974 , n7808 , n29508 );
xor ( n69975 , n69973 , n69974 );
and ( n69976 , n8079 , n28406 );
xor ( n69977 , n69975 , n69976 );
xor ( n69978 , n69972 , n69977 );
xor ( n69979 , n69963 , n69978 );
and ( n69980 , n68799 , n68869 );
and ( n69981 , n68869 , n68906 );
and ( n69982 , n68799 , n68906 );
or ( n69983 , n69980 , n69981 , n69982 );
and ( n69984 , n68874 , n68878 );
and ( n69985 , n68878 , n68905 );
and ( n69986 , n68874 , n68905 );
or ( n69987 , n69984 , n69985 , n69986 );
and ( n69988 , n68833 , n68851 );
and ( n69989 , n68851 , n68867 );
and ( n69990 , n68833 , n68867 );
or ( n69991 , n69988 , n69989 , n69990 );
and ( n69992 , n68816 , n68820 );
and ( n69993 , n68820 , n68826 );
and ( n69994 , n68816 , n68826 );
or ( n69995 , n69992 , n69993 , n69994 );
and ( n69996 , n68839 , n68844 );
and ( n69997 , n68844 , n68850 );
and ( n69998 , n68839 , n68850 );
or ( n69999 , n69996 , n69997 , n69998 );
xor ( n70000 , n69995 , n69999 );
and ( n70001 , n68822 , n68823 );
and ( n70002 , n68823 , n68825 );
and ( n70003 , n68822 , n68825 );
or ( n70004 , n70001 , n70002 , n70003 );
and ( n70005 , n68840 , n68841 );
and ( n70006 , n68841 , n68843 );
and ( n70007 , n68840 , n68843 );
or ( n70008 , n70005 , n70006 , n70007 );
xor ( n70009 , n70004 , n70008 );
and ( n70010 , n21216 , n13256 );
and ( n70011 , n22186 , n12531 );
xor ( n70012 , n70010 , n70011 );
and ( n70013 , n22892 , n11718 );
xor ( n70014 , n70012 , n70013 );
xor ( n70015 , n70009 , n70014 );
xor ( n70016 , n70000 , n70015 );
xor ( n70017 , n69991 , n70016 );
and ( n70018 , n68856 , n68860 );
and ( n70019 , n68860 , n68866 );
and ( n70020 , n68856 , n68866 );
or ( n70021 , n70018 , n70019 , n70020 );
and ( n70022 , n68846 , n68847 );
and ( n70023 , n68847 , n68849 );
and ( n70024 , n68846 , n68849 );
or ( n70025 , n70022 , n70023 , n70024 );
and ( n70026 , n18144 , n15691 );
and ( n70027 , n19324 , n14838 );
xor ( n70028 , n70026 , n70027 );
and ( n70029 , n20233 , n14044 );
xor ( n70030 , n70028 , n70029 );
xor ( n70031 , n70025 , n70030 );
and ( n70032 , n15758 , n18407 );
and ( n70033 , n16637 , n17422 );
xor ( n70034 , n70032 , n70033 );
and ( n70035 , n17512 , n16550 );
xor ( n70036 , n70034 , n70035 );
xor ( n70037 , n70031 , n70036 );
xor ( n70038 , n70021 , n70037 );
and ( n70039 , n68862 , n68863 );
and ( n70040 , n68863 , n68865 );
and ( n70041 , n68862 , n68865 );
or ( n70042 , n70039 , n70040 , n70041 );
and ( n70043 , n68893 , n68894 );
and ( n70044 , n68894 , n68896 );
and ( n70045 , n68893 , n68896 );
or ( n70046 , n70043 , n70044 , n70045 );
xor ( n70047 , n70042 , n70046 );
and ( n70048 , n13322 , n20976 );
and ( n70049 , n14118 , n20156 );
xor ( n70050 , n70048 , n70049 );
and ( n70051 , n14938 , n19222 );
xor ( n70052 , n70050 , n70051 );
xor ( n70053 , n70047 , n70052 );
xor ( n70054 , n70038 , n70053 );
xor ( n70055 , n70017 , n70054 );
xor ( n70056 , n69987 , n70055 );
and ( n70057 , n68761 , n68776 );
and ( n70058 , n68776 , n68788 );
and ( n70059 , n68761 , n68788 );
or ( n70060 , n70057 , n70058 , n70059 );
and ( n70061 , n68883 , n68887 );
and ( n70062 , n68887 , n68904 );
and ( n70063 , n68883 , n68904 );
or ( n70064 , n70061 , n70062 , n70063 );
xor ( n70065 , n70060 , n70064 );
and ( n70066 , n68892 , n68897 );
and ( n70067 , n68897 , n68903 );
and ( n70068 , n68892 , n68903 );
or ( n70069 , n70066 , n70067 , n70068 );
and ( n70070 , n68765 , n68769 );
and ( n70071 , n68769 , n68775 );
and ( n70072 , n68765 , n68775 );
or ( n70073 , n70070 , n70071 , n70072 );
xor ( n70074 , n70069 , n70073 );
and ( n70075 , n68899 , n68900 );
and ( n70076 , n68900 , n68902 );
and ( n70077 , n68899 , n68902 );
or ( n70078 , n70075 , n70076 , n70077 );
and ( n70079 , n11015 , n24137 );
and ( n70080 , n11769 , n23075 );
xor ( n70081 , n70079 , n70080 );
and ( n70082 , n12320 , n22065 );
xor ( n70083 , n70081 , n70082 );
xor ( n70084 , n70078 , n70083 );
and ( n70085 , n8718 , n27296 );
and ( n70086 , n9400 , n26216 );
xor ( n70087 , n70085 , n70086 );
and ( n70088 , n10291 , n25163 );
xor ( n70089 , n70087 , n70088 );
xor ( n70090 , n70084 , n70089 );
xor ( n70091 , n70074 , n70090 );
xor ( n70092 , n70065 , n70091 );
xor ( n70093 , n70056 , n70092 );
xor ( n70094 , n69983 , n70093 );
xor ( n70095 , n69979 , n70094 );
xor ( n70096 , n69951 , n70095 );
xor ( n70097 , n69872 , n70096 );
xor ( n70098 , n69863 , n70097 );
and ( n70099 , n68665 , n68668 );
and ( n70100 , n68668 , n68911 );
and ( n70101 , n68665 , n68911 );
or ( n70102 , n70099 , n70100 , n70101 );
xor ( n70103 , n70098 , n70102 );
and ( n70104 , n68912 , n68916 );
and ( n70105 , n68917 , n68920 );
or ( n70106 , n70104 , n70105 );
xor ( n70107 , n70103 , n70106 );
buf ( n70108 , n70107 );
buf ( n70109 , n70108 );
not ( n70110 , n70109 );
nor ( n70111 , n70110 , n8739 );
xor ( n70112 , n69855 , n70111 );
and ( n70113 , n68661 , n68925 );
and ( n70114 , n68926 , n68929 );
or ( n70115 , n70113 , n70114 );
xor ( n70116 , n70112 , n70115 );
buf ( n70117 , n70116 );
buf ( n70118 , n70117 );
not ( n70119 , n70118 );
buf ( n70120 , n592 );
not ( n70121 , n70120 );
nor ( n70122 , n70119 , n70121 );
xor ( n70123 , n69481 , n70122 );
xor ( n70124 , n68941 , n69478 );
nor ( n70125 , n68933 , n70121 );
and ( n70126 , n70124 , n70125 );
xor ( n70127 , n70124 , n70125 );
xor ( n70128 , n68945 , n69476 );
nor ( n70129 , n67745 , n70121 );
and ( n70130 , n70128 , n70129 );
xor ( n70131 , n70128 , n70129 );
xor ( n70132 , n68949 , n69474 );
nor ( n70133 , n66559 , n70121 );
and ( n70134 , n70132 , n70133 );
xor ( n70135 , n70132 , n70133 );
xor ( n70136 , n68953 , n69472 );
nor ( n70137 , n65369 , n70121 );
and ( n70138 , n70136 , n70137 );
xor ( n70139 , n70136 , n70137 );
xor ( n70140 , n68957 , n69470 );
nor ( n70141 , n64181 , n70121 );
and ( n70142 , n70140 , n70141 );
xor ( n70143 , n70140 , n70141 );
xor ( n70144 , n68961 , n69468 );
nor ( n70145 , n62991 , n70121 );
and ( n70146 , n70144 , n70145 );
xor ( n70147 , n70144 , n70145 );
xor ( n70148 , n68965 , n69466 );
nor ( n70149 , n61800 , n70121 );
and ( n70150 , n70148 , n70149 );
xor ( n70151 , n70148 , n70149 );
xor ( n70152 , n68969 , n69464 );
nor ( n70153 , n60609 , n70121 );
and ( n70154 , n70152 , n70153 );
xor ( n70155 , n70152 , n70153 );
xor ( n70156 , n68973 , n69462 );
nor ( n70157 , n59421 , n70121 );
and ( n70158 , n70156 , n70157 );
xor ( n70159 , n70156 , n70157 );
xor ( n70160 , n68977 , n69460 );
nor ( n70161 , n58226 , n70121 );
and ( n70162 , n70160 , n70161 );
xor ( n70163 , n70160 , n70161 );
xor ( n70164 , n68981 , n69458 );
nor ( n70165 , n57031 , n70121 );
and ( n70166 , n70164 , n70165 );
xor ( n70167 , n70164 , n70165 );
xor ( n70168 , n68985 , n69456 );
nor ( n70169 , n55835 , n70121 );
and ( n70170 , n70168 , n70169 );
xor ( n70171 , n70168 , n70169 );
xor ( n70172 , n68989 , n69454 );
nor ( n70173 , n54638 , n70121 );
and ( n70174 , n70172 , n70173 );
xor ( n70175 , n70172 , n70173 );
xor ( n70176 , n68993 , n69452 );
nor ( n70177 , n53441 , n70121 );
and ( n70178 , n70176 , n70177 );
xor ( n70179 , n70176 , n70177 );
xor ( n70180 , n68997 , n69450 );
nor ( n70181 , n52247 , n70121 );
and ( n70182 , n70180 , n70181 );
xor ( n70183 , n70180 , n70181 );
xor ( n70184 , n69001 , n69448 );
nor ( n70185 , n51049 , n70121 );
and ( n70186 , n70184 , n70185 );
xor ( n70187 , n70184 , n70185 );
xor ( n70188 , n69005 , n69446 );
nor ( n70189 , n49850 , n70121 );
and ( n70190 , n70188 , n70189 );
xor ( n70191 , n70188 , n70189 );
xor ( n70192 , n69009 , n69444 );
nor ( n70193 , n48650 , n70121 );
and ( n70194 , n70192 , n70193 );
xor ( n70195 , n70192 , n70193 );
xor ( n70196 , n69013 , n69442 );
nor ( n70197 , n47449 , n70121 );
and ( n70198 , n70196 , n70197 );
xor ( n70199 , n70196 , n70197 );
xor ( n70200 , n69017 , n69440 );
nor ( n70201 , n46248 , n70121 );
and ( n70202 , n70200 , n70201 );
xor ( n70203 , n70200 , n70201 );
xor ( n70204 , n69021 , n69438 );
nor ( n70205 , n45047 , n70121 );
and ( n70206 , n70204 , n70205 );
xor ( n70207 , n70204 , n70205 );
xor ( n70208 , n69025 , n69436 );
nor ( n70209 , n43843 , n70121 );
and ( n70210 , n70208 , n70209 );
xor ( n70211 , n70208 , n70209 );
xor ( n70212 , n69029 , n69434 );
nor ( n70213 , n42641 , n70121 );
and ( n70214 , n70212 , n70213 );
xor ( n70215 , n70212 , n70213 );
xor ( n70216 , n69033 , n69432 );
nor ( n70217 , n41437 , n70121 );
and ( n70218 , n70216 , n70217 );
xor ( n70219 , n70216 , n70217 );
xor ( n70220 , n69037 , n69430 );
nor ( n70221 , n40232 , n70121 );
and ( n70222 , n70220 , n70221 );
xor ( n70223 , n70220 , n70221 );
xor ( n70224 , n69041 , n69428 );
nor ( n70225 , n39027 , n70121 );
and ( n70226 , n70224 , n70225 );
xor ( n70227 , n70224 , n70225 );
xor ( n70228 , n69045 , n69426 );
nor ( n70229 , n37825 , n70121 );
and ( n70230 , n70228 , n70229 );
xor ( n70231 , n70228 , n70229 );
xor ( n70232 , n69049 , n69424 );
nor ( n70233 , n36620 , n70121 );
and ( n70234 , n70232 , n70233 );
xor ( n70235 , n70232 , n70233 );
xor ( n70236 , n69053 , n69422 );
nor ( n70237 , n35419 , n70121 );
and ( n70238 , n70236 , n70237 );
xor ( n70239 , n70236 , n70237 );
xor ( n70240 , n69057 , n69420 );
nor ( n70241 , n34224 , n70121 );
and ( n70242 , n70240 , n70241 );
xor ( n70243 , n70240 , n70241 );
xor ( n70244 , n69061 , n69418 );
nor ( n70245 , n33033 , n70121 );
and ( n70246 , n70244 , n70245 );
xor ( n70247 , n70244 , n70245 );
xor ( n70248 , n69065 , n69416 );
nor ( n70249 , n31867 , n70121 );
and ( n70250 , n70248 , n70249 );
xor ( n70251 , n70248 , n70249 );
xor ( n70252 , n69069 , n69414 );
nor ( n70253 , n30725 , n70121 );
and ( n70254 , n70252 , n70253 );
xor ( n70255 , n70252 , n70253 );
xor ( n70256 , n69073 , n69412 );
nor ( n70257 , n29596 , n70121 );
and ( n70258 , n70256 , n70257 );
xor ( n70259 , n70256 , n70257 );
xor ( n70260 , n69077 , n69410 );
nor ( n70261 , n28487 , n70121 );
and ( n70262 , n70260 , n70261 );
xor ( n70263 , n70260 , n70261 );
xor ( n70264 , n69081 , n69408 );
nor ( n70265 , n27397 , n70121 );
and ( n70266 , n70264 , n70265 );
xor ( n70267 , n70264 , n70265 );
xor ( n70268 , n69085 , n69406 );
nor ( n70269 , n26326 , n70121 );
and ( n70270 , n70268 , n70269 );
xor ( n70271 , n70268 , n70269 );
xor ( n70272 , n69089 , n69404 );
nor ( n70273 , n25272 , n70121 );
and ( n70274 , n70272 , n70273 );
xor ( n70275 , n70272 , n70273 );
xor ( n70276 , n69093 , n69402 );
nor ( n70277 , n24242 , n70121 );
and ( n70278 , n70276 , n70277 );
xor ( n70279 , n70276 , n70277 );
xor ( n70280 , n69097 , n69400 );
nor ( n70281 , n23225 , n70121 );
and ( n70282 , n70280 , n70281 );
xor ( n70283 , n70280 , n70281 );
xor ( n70284 , n69101 , n69398 );
nor ( n70285 , n22231 , n70121 );
and ( n70286 , n70284 , n70285 );
xor ( n70287 , n70284 , n70285 );
xor ( n70288 , n69105 , n69396 );
nor ( n70289 , n21258 , n70121 );
and ( n70290 , n70288 , n70289 );
xor ( n70291 , n70288 , n70289 );
xor ( n70292 , n69109 , n69394 );
nor ( n70293 , n20303 , n70121 );
and ( n70294 , n70292 , n70293 );
xor ( n70295 , n70292 , n70293 );
xor ( n70296 , n69113 , n69392 );
nor ( n70297 , n19365 , n70121 );
and ( n70298 , n70296 , n70297 );
xor ( n70299 , n70296 , n70297 );
xor ( n70300 , n69117 , n69390 );
nor ( n70301 , n18448 , n70121 );
and ( n70302 , n70300 , n70301 );
xor ( n70303 , n70300 , n70301 );
xor ( n70304 , n69121 , n69388 );
nor ( n70305 , n17548 , n70121 );
and ( n70306 , n70304 , n70305 );
xor ( n70307 , n70304 , n70305 );
xor ( n70308 , n69125 , n69386 );
nor ( n70309 , n16669 , n70121 );
and ( n70310 , n70308 , n70309 );
xor ( n70311 , n70308 , n70309 );
xor ( n70312 , n69129 , n69384 );
nor ( n70313 , n15809 , n70121 );
and ( n70314 , n70312 , n70313 );
xor ( n70315 , n70312 , n70313 );
xor ( n70316 , n69133 , n69382 );
nor ( n70317 , n14968 , n70121 );
and ( n70318 , n70316 , n70317 );
xor ( n70319 , n70316 , n70317 );
xor ( n70320 , n69137 , n69380 );
nor ( n70321 , n14147 , n70121 );
and ( n70322 , n70320 , n70321 );
xor ( n70323 , n70320 , n70321 );
xor ( n70324 , n69141 , n69378 );
nor ( n70325 , n13349 , n70121 );
and ( n70326 , n70324 , n70325 );
xor ( n70327 , n70324 , n70325 );
xor ( n70328 , n69145 , n69376 );
nor ( n70329 , n12564 , n70121 );
and ( n70330 , n70328 , n70329 );
xor ( n70331 , n70328 , n70329 );
xor ( n70332 , n69149 , n69374 );
nor ( n70333 , n11799 , n70121 );
and ( n70334 , n70332 , n70333 );
xor ( n70335 , n70332 , n70333 );
xor ( n70336 , n69153 , n69372 );
nor ( n70337 , n11050 , n70121 );
and ( n70338 , n70336 , n70337 );
xor ( n70339 , n70336 , n70337 );
xor ( n70340 , n69157 , n69370 );
nor ( n70341 , n10321 , n70121 );
and ( n70342 , n70340 , n70341 );
xor ( n70343 , n70340 , n70341 );
xor ( n70344 , n69161 , n69368 );
nor ( n70345 , n9429 , n70121 );
and ( n70346 , n70344 , n70345 );
xor ( n70347 , n70344 , n70345 );
xor ( n70348 , n69165 , n69366 );
nor ( n70349 , n8949 , n70121 );
and ( n70350 , n70348 , n70349 );
xor ( n70351 , n70348 , n70349 );
xor ( n70352 , n69169 , n69364 );
nor ( n70353 , n9437 , n70121 );
and ( n70354 , n70352 , n70353 );
xor ( n70355 , n70352 , n70353 );
xor ( n70356 , n69173 , n69362 );
nor ( n70357 , n9446 , n70121 );
and ( n70358 , n70356 , n70357 );
xor ( n70359 , n70356 , n70357 );
xor ( n70360 , n69177 , n69360 );
nor ( n70361 , n9455 , n70121 );
and ( n70362 , n70360 , n70361 );
xor ( n70363 , n70360 , n70361 );
xor ( n70364 , n69181 , n69358 );
nor ( n70365 , n9464 , n70121 );
and ( n70366 , n70364 , n70365 );
xor ( n70367 , n70364 , n70365 );
xor ( n70368 , n69185 , n69356 );
nor ( n70369 , n9473 , n70121 );
and ( n70370 , n70368 , n70369 );
xor ( n70371 , n70368 , n70369 );
xor ( n70372 , n69189 , n69354 );
nor ( n70373 , n9482 , n70121 );
and ( n70374 , n70372 , n70373 );
xor ( n70375 , n70372 , n70373 );
xor ( n70376 , n69193 , n69352 );
nor ( n70377 , n9491 , n70121 );
and ( n70378 , n70376 , n70377 );
xor ( n70379 , n70376 , n70377 );
xor ( n70380 , n69197 , n69350 );
nor ( n70381 , n9500 , n70121 );
and ( n70382 , n70380 , n70381 );
xor ( n70383 , n70380 , n70381 );
xor ( n70384 , n69201 , n69348 );
nor ( n70385 , n9509 , n70121 );
and ( n70386 , n70384 , n70385 );
xor ( n70387 , n70384 , n70385 );
xor ( n70388 , n69205 , n69346 );
nor ( n70389 , n9518 , n70121 );
and ( n70390 , n70388 , n70389 );
xor ( n70391 , n70388 , n70389 );
xor ( n70392 , n69209 , n69344 );
nor ( n70393 , n9527 , n70121 );
and ( n70394 , n70392 , n70393 );
xor ( n70395 , n70392 , n70393 );
xor ( n70396 , n69213 , n69342 );
nor ( n70397 , n9536 , n70121 );
and ( n70398 , n70396 , n70397 );
xor ( n70399 , n70396 , n70397 );
xor ( n70400 , n69217 , n69340 );
nor ( n70401 , n9545 , n70121 );
and ( n70402 , n70400 , n70401 );
xor ( n70403 , n70400 , n70401 );
xor ( n70404 , n69221 , n69338 );
nor ( n70405 , n9554 , n70121 );
and ( n70406 , n70404 , n70405 );
xor ( n70407 , n70404 , n70405 );
xor ( n70408 , n69225 , n69336 );
nor ( n70409 , n9563 , n70121 );
and ( n70410 , n70408 , n70409 );
xor ( n70411 , n70408 , n70409 );
xor ( n70412 , n69229 , n69334 );
nor ( n70413 , n9572 , n70121 );
and ( n70414 , n70412 , n70413 );
xor ( n70415 , n70412 , n70413 );
xor ( n70416 , n69233 , n69332 );
nor ( n70417 , n9581 , n70121 );
and ( n70418 , n70416 , n70417 );
xor ( n70419 , n70416 , n70417 );
xor ( n70420 , n69237 , n69330 );
nor ( n70421 , n9590 , n70121 );
and ( n70422 , n70420 , n70421 );
xor ( n70423 , n70420 , n70421 );
xor ( n70424 , n69241 , n69328 );
nor ( n70425 , n9599 , n70121 );
and ( n70426 , n70424 , n70425 );
xor ( n70427 , n70424 , n70425 );
xor ( n70428 , n69245 , n69326 );
nor ( n70429 , n9608 , n70121 );
and ( n70430 , n70428 , n70429 );
xor ( n70431 , n70428 , n70429 );
xor ( n70432 , n69249 , n69324 );
nor ( n70433 , n9617 , n70121 );
and ( n70434 , n70432 , n70433 );
xor ( n70435 , n70432 , n70433 );
xor ( n70436 , n69253 , n69322 );
nor ( n70437 , n9626 , n70121 );
and ( n70438 , n70436 , n70437 );
xor ( n70439 , n70436 , n70437 );
xor ( n70440 , n69257 , n69320 );
nor ( n70441 , n9635 , n70121 );
and ( n70442 , n70440 , n70441 );
xor ( n70443 , n70440 , n70441 );
xor ( n70444 , n69261 , n69318 );
nor ( n70445 , n9644 , n70121 );
and ( n70446 , n70444 , n70445 );
xor ( n70447 , n70444 , n70445 );
xor ( n70448 , n69265 , n69316 );
nor ( n70449 , n9653 , n70121 );
and ( n70450 , n70448 , n70449 );
xor ( n70451 , n70448 , n70449 );
xor ( n70452 , n69269 , n69314 );
nor ( n70453 , n9662 , n70121 );
and ( n70454 , n70452 , n70453 );
xor ( n70455 , n70452 , n70453 );
xor ( n70456 , n69273 , n69312 );
nor ( n70457 , n9671 , n70121 );
and ( n70458 , n70456 , n70457 );
xor ( n70459 , n70456 , n70457 );
xor ( n70460 , n69277 , n69310 );
nor ( n70461 , n9680 , n70121 );
and ( n70462 , n70460 , n70461 );
xor ( n70463 , n70460 , n70461 );
xor ( n70464 , n69281 , n69308 );
nor ( n70465 , n9689 , n70121 );
and ( n70466 , n70464 , n70465 );
xor ( n70467 , n70464 , n70465 );
xor ( n70468 , n69285 , n69306 );
nor ( n70469 , n9698 , n70121 );
and ( n70470 , n70468 , n70469 );
xor ( n70471 , n70468 , n70469 );
xor ( n70472 , n69289 , n69304 );
nor ( n70473 , n9707 , n70121 );
and ( n70474 , n70472 , n70473 );
xor ( n70475 , n70472 , n70473 );
xor ( n70476 , n69293 , n69302 );
nor ( n70477 , n9716 , n70121 );
and ( n70478 , n70476 , n70477 );
xor ( n70479 , n70476 , n70477 );
xor ( n70480 , n69297 , n69300 );
nor ( n70481 , n9725 , n70121 );
and ( n70482 , n70480 , n70481 );
xor ( n70483 , n70480 , n70481 );
xor ( n70484 , n69298 , n69299 );
nor ( n70485 , n9734 , n70121 );
and ( n70486 , n70484 , n70485 );
xor ( n70487 , n70484 , n70485 );
nor ( n70488 , n9752 , n68935 );
nor ( n70489 , n9743 , n70121 );
and ( n70490 , n70488 , n70489 );
and ( n70491 , n70487 , n70490 );
or ( n70492 , n70486 , n70491 );
and ( n70493 , n70483 , n70492 );
or ( n70494 , n70482 , n70493 );
and ( n70495 , n70479 , n70494 );
or ( n70496 , n70478 , n70495 );
and ( n70497 , n70475 , n70496 );
or ( n70498 , n70474 , n70497 );
and ( n70499 , n70471 , n70498 );
or ( n70500 , n70470 , n70499 );
and ( n70501 , n70467 , n70500 );
or ( n70502 , n70466 , n70501 );
and ( n70503 , n70463 , n70502 );
or ( n70504 , n70462 , n70503 );
and ( n70505 , n70459 , n70504 );
or ( n70506 , n70458 , n70505 );
and ( n70507 , n70455 , n70506 );
or ( n70508 , n70454 , n70507 );
and ( n70509 , n70451 , n70508 );
or ( n70510 , n70450 , n70509 );
and ( n70511 , n70447 , n70510 );
or ( n70512 , n70446 , n70511 );
and ( n70513 , n70443 , n70512 );
or ( n70514 , n70442 , n70513 );
and ( n70515 , n70439 , n70514 );
or ( n70516 , n70438 , n70515 );
and ( n70517 , n70435 , n70516 );
or ( n70518 , n70434 , n70517 );
and ( n70519 , n70431 , n70518 );
or ( n70520 , n70430 , n70519 );
and ( n70521 , n70427 , n70520 );
or ( n70522 , n70426 , n70521 );
and ( n70523 , n70423 , n70522 );
or ( n70524 , n70422 , n70523 );
and ( n70525 , n70419 , n70524 );
or ( n70526 , n70418 , n70525 );
and ( n70527 , n70415 , n70526 );
or ( n70528 , n70414 , n70527 );
and ( n70529 , n70411 , n70528 );
or ( n70530 , n70410 , n70529 );
and ( n70531 , n70407 , n70530 );
or ( n70532 , n70406 , n70531 );
and ( n70533 , n70403 , n70532 );
or ( n70534 , n70402 , n70533 );
and ( n70535 , n70399 , n70534 );
or ( n70536 , n70398 , n70535 );
and ( n70537 , n70395 , n70536 );
or ( n70538 , n70394 , n70537 );
and ( n70539 , n70391 , n70538 );
or ( n70540 , n70390 , n70539 );
and ( n70541 , n70387 , n70540 );
or ( n70542 , n70386 , n70541 );
and ( n70543 , n70383 , n70542 );
or ( n70544 , n70382 , n70543 );
and ( n70545 , n70379 , n70544 );
or ( n70546 , n70378 , n70545 );
and ( n70547 , n70375 , n70546 );
or ( n70548 , n70374 , n70547 );
and ( n70549 , n70371 , n70548 );
or ( n70550 , n70370 , n70549 );
and ( n70551 , n70367 , n70550 );
or ( n70552 , n70366 , n70551 );
and ( n70553 , n70363 , n70552 );
or ( n70554 , n70362 , n70553 );
and ( n70555 , n70359 , n70554 );
or ( n70556 , n70358 , n70555 );
and ( n70557 , n70355 , n70556 );
or ( n70558 , n70354 , n70557 );
and ( n70559 , n70351 , n70558 );
or ( n70560 , n70350 , n70559 );
and ( n70561 , n70347 , n70560 );
or ( n70562 , n70346 , n70561 );
and ( n70563 , n70343 , n70562 );
or ( n70564 , n70342 , n70563 );
and ( n70565 , n70339 , n70564 );
or ( n70566 , n70338 , n70565 );
and ( n70567 , n70335 , n70566 );
or ( n70568 , n70334 , n70567 );
and ( n70569 , n70331 , n70568 );
or ( n70570 , n70330 , n70569 );
and ( n70571 , n70327 , n70570 );
or ( n70572 , n70326 , n70571 );
and ( n70573 , n70323 , n70572 );
or ( n70574 , n70322 , n70573 );
and ( n70575 , n70319 , n70574 );
or ( n70576 , n70318 , n70575 );
and ( n70577 , n70315 , n70576 );
or ( n70578 , n70314 , n70577 );
and ( n70579 , n70311 , n70578 );
or ( n70580 , n70310 , n70579 );
and ( n70581 , n70307 , n70580 );
or ( n70582 , n70306 , n70581 );
and ( n70583 , n70303 , n70582 );
or ( n70584 , n70302 , n70583 );
and ( n70585 , n70299 , n70584 );
or ( n70586 , n70298 , n70585 );
and ( n70587 , n70295 , n70586 );
or ( n70588 , n70294 , n70587 );
and ( n70589 , n70291 , n70588 );
or ( n70590 , n70290 , n70589 );
and ( n70591 , n70287 , n70590 );
or ( n70592 , n70286 , n70591 );
and ( n70593 , n70283 , n70592 );
or ( n70594 , n70282 , n70593 );
and ( n70595 , n70279 , n70594 );
or ( n70596 , n70278 , n70595 );
and ( n70597 , n70275 , n70596 );
or ( n70598 , n70274 , n70597 );
and ( n70599 , n70271 , n70598 );
or ( n70600 , n70270 , n70599 );
and ( n70601 , n70267 , n70600 );
or ( n70602 , n70266 , n70601 );
and ( n70603 , n70263 , n70602 );
or ( n70604 , n70262 , n70603 );
and ( n70605 , n70259 , n70604 );
or ( n70606 , n70258 , n70605 );
and ( n70607 , n70255 , n70606 );
or ( n70608 , n70254 , n70607 );
and ( n70609 , n70251 , n70608 );
or ( n70610 , n70250 , n70609 );
and ( n70611 , n70247 , n70610 );
or ( n70612 , n70246 , n70611 );
and ( n70613 , n70243 , n70612 );
or ( n70614 , n70242 , n70613 );
and ( n70615 , n70239 , n70614 );
or ( n70616 , n70238 , n70615 );
and ( n70617 , n70235 , n70616 );
or ( n70618 , n70234 , n70617 );
and ( n70619 , n70231 , n70618 );
or ( n70620 , n70230 , n70619 );
and ( n70621 , n70227 , n70620 );
or ( n70622 , n70226 , n70621 );
and ( n70623 , n70223 , n70622 );
or ( n70624 , n70222 , n70623 );
and ( n70625 , n70219 , n70624 );
or ( n70626 , n70218 , n70625 );
and ( n70627 , n70215 , n70626 );
or ( n70628 , n70214 , n70627 );
and ( n70629 , n70211 , n70628 );
or ( n70630 , n70210 , n70629 );
and ( n70631 , n70207 , n70630 );
or ( n70632 , n70206 , n70631 );
and ( n70633 , n70203 , n70632 );
or ( n70634 , n70202 , n70633 );
and ( n70635 , n70199 , n70634 );
or ( n70636 , n70198 , n70635 );
and ( n70637 , n70195 , n70636 );
or ( n70638 , n70194 , n70637 );
and ( n70639 , n70191 , n70638 );
or ( n70640 , n70190 , n70639 );
and ( n70641 , n70187 , n70640 );
or ( n70642 , n70186 , n70641 );
and ( n70643 , n70183 , n70642 );
or ( n70644 , n70182 , n70643 );
and ( n70645 , n70179 , n70644 );
or ( n70646 , n70178 , n70645 );
and ( n70647 , n70175 , n70646 );
or ( n70648 , n70174 , n70647 );
and ( n70649 , n70171 , n70648 );
or ( n70650 , n70170 , n70649 );
and ( n70651 , n70167 , n70650 );
or ( n70652 , n70166 , n70651 );
and ( n70653 , n70163 , n70652 );
or ( n70654 , n70162 , n70653 );
and ( n70655 , n70159 , n70654 );
or ( n70656 , n70158 , n70655 );
and ( n70657 , n70155 , n70656 );
or ( n70658 , n70154 , n70657 );
and ( n70659 , n70151 , n70658 );
or ( n70660 , n70150 , n70659 );
and ( n70661 , n70147 , n70660 );
or ( n70662 , n70146 , n70661 );
and ( n70663 , n70143 , n70662 );
or ( n70664 , n70142 , n70663 );
and ( n70665 , n70139 , n70664 );
or ( n70666 , n70138 , n70665 );
and ( n70667 , n70135 , n70666 );
or ( n70668 , n70134 , n70667 );
and ( n70669 , n70131 , n70668 );
or ( n70670 , n70130 , n70669 );
and ( n70671 , n70127 , n70670 );
or ( n70672 , n70126 , n70671 );
xor ( n70673 , n70123 , n70672 );
and ( n70674 , n33403 , n6595 );
nor ( n70675 , n6596 , n70674 );
nor ( n70676 , n6997 , n32231 );
xor ( n70677 , n70675 , n70676 );
and ( n70678 , n69483 , n69484 );
and ( n70679 , n69485 , n69488 );
or ( n70680 , n70678 , n70679 );
xor ( n70681 , n70677 , n70680 );
nor ( n70682 , n7413 , n31083 );
xor ( n70683 , n70681 , n70682 );
and ( n70684 , n69489 , n69490 );
and ( n70685 , n69491 , n69494 );
or ( n70686 , n70684 , n70685 );
xor ( n70687 , n70683 , n70686 );
nor ( n70688 , n7841 , n29948 );
xor ( n70689 , n70687 , n70688 );
and ( n70690 , n69495 , n69496 );
and ( n70691 , n69497 , n69500 );
or ( n70692 , n70690 , n70691 );
xor ( n70693 , n70689 , n70692 );
nor ( n70694 , n8281 , n28833 );
xor ( n70695 , n70693 , n70694 );
and ( n70696 , n69501 , n69502 );
and ( n70697 , n69503 , n69506 );
or ( n70698 , n70696 , n70697 );
xor ( n70699 , n70695 , n70698 );
nor ( n70700 , n8737 , n27737 );
xor ( n70701 , n70699 , n70700 );
and ( n70702 , n69507 , n69508 );
and ( n70703 , n69509 , n69512 );
or ( n70704 , n70702 , n70703 );
xor ( n70705 , n70701 , n70704 );
nor ( n70706 , n9420 , n26660 );
xor ( n70707 , n70705 , n70706 );
and ( n70708 , n69513 , n69514 );
and ( n70709 , n69515 , n69518 );
or ( n70710 , n70708 , n70709 );
xor ( n70711 , n70707 , n70710 );
nor ( n70712 , n10312 , n25600 );
xor ( n70713 , n70711 , n70712 );
and ( n70714 , n69519 , n69520 );
and ( n70715 , n69521 , n69524 );
or ( n70716 , n70714 , n70715 );
xor ( n70717 , n70713 , n70716 );
nor ( n70718 , n11041 , n24564 );
xor ( n70719 , n70717 , n70718 );
and ( n70720 , n69525 , n69526 );
and ( n70721 , n69527 , n69530 );
or ( n70722 , n70720 , n70721 );
xor ( n70723 , n70719 , n70722 );
nor ( n70724 , n11790 , n23541 );
xor ( n70725 , n70723 , n70724 );
and ( n70726 , n69531 , n69532 );
and ( n70727 , n69533 , n69536 );
or ( n70728 , n70726 , n70727 );
xor ( n70729 , n70725 , n70728 );
nor ( n70730 , n12555 , n22541 );
xor ( n70731 , n70729 , n70730 );
and ( n70732 , n69537 , n69538 );
and ( n70733 , n69539 , n69542 );
or ( n70734 , n70732 , n70733 );
xor ( n70735 , n70731 , n70734 );
nor ( n70736 , n13340 , n21562 );
xor ( n70737 , n70735 , n70736 );
and ( n70738 , n69543 , n69544 );
and ( n70739 , n69545 , n69548 );
or ( n70740 , n70738 , n70739 );
xor ( n70741 , n70737 , n70740 );
nor ( n70742 , n14138 , n20601 );
xor ( n70743 , n70741 , n70742 );
and ( n70744 , n69549 , n69550 );
and ( n70745 , n69551 , n69554 );
or ( n70746 , n70744 , n70745 );
xor ( n70747 , n70743 , n70746 );
nor ( n70748 , n14959 , n19657 );
xor ( n70749 , n70747 , n70748 );
and ( n70750 , n69555 , n69556 );
and ( n70751 , n69557 , n69560 );
or ( n70752 , n70750 , n70751 );
xor ( n70753 , n70749 , n70752 );
nor ( n70754 , n15800 , n18734 );
xor ( n70755 , n70753 , n70754 );
and ( n70756 , n69561 , n69562 );
and ( n70757 , n69563 , n69566 );
or ( n70758 , n70756 , n70757 );
xor ( n70759 , n70755 , n70758 );
nor ( n70760 , n16660 , n17828 );
xor ( n70761 , n70759 , n70760 );
and ( n70762 , n69567 , n69568 );
and ( n70763 , n69569 , n69572 );
or ( n70764 , n70762 , n70763 );
xor ( n70765 , n70761 , n70764 );
nor ( n70766 , n17539 , n16943 );
xor ( n70767 , n70765 , n70766 );
and ( n70768 , n69573 , n69574 );
and ( n70769 , n69575 , n69578 );
or ( n70770 , n70768 , n70769 );
xor ( n70771 , n70767 , n70770 );
nor ( n70772 , n18439 , n16077 );
xor ( n70773 , n70771 , n70772 );
and ( n70774 , n69579 , n69580 );
and ( n70775 , n69581 , n69584 );
or ( n70776 , n70774 , n70775 );
xor ( n70777 , n70773 , n70776 );
nor ( n70778 , n19356 , n15230 );
xor ( n70779 , n70777 , n70778 );
and ( n70780 , n69585 , n69586 );
and ( n70781 , n69587 , n69590 );
or ( n70782 , n70780 , n70781 );
xor ( n70783 , n70779 , n70782 );
nor ( n70784 , n20294 , n14403 );
xor ( n70785 , n70783 , n70784 );
and ( n70786 , n69591 , n69592 );
and ( n70787 , n69593 , n69596 );
or ( n70788 , n70786 , n70787 );
xor ( n70789 , n70785 , n70788 );
nor ( n70790 , n21249 , n13599 );
xor ( n70791 , n70789 , n70790 );
and ( n70792 , n69597 , n69598 );
and ( n70793 , n69599 , n69602 );
or ( n70794 , n70792 , n70793 );
xor ( n70795 , n70791 , n70794 );
nor ( n70796 , n22222 , n12808 );
xor ( n70797 , n70795 , n70796 );
and ( n70798 , n69603 , n69604 );
and ( n70799 , n69605 , n69608 );
or ( n70800 , n70798 , n70799 );
xor ( n70801 , n70797 , n70800 );
nor ( n70802 , n23216 , n12037 );
xor ( n70803 , n70801 , n70802 );
and ( n70804 , n69609 , n69610 );
and ( n70805 , n69611 , n69614 );
or ( n70806 , n70804 , n70805 );
xor ( n70807 , n70803 , n70806 );
nor ( n70808 , n24233 , n11282 );
xor ( n70809 , n70807 , n70808 );
and ( n70810 , n69615 , n69616 );
and ( n70811 , n69617 , n69620 );
or ( n70812 , n70810 , n70811 );
xor ( n70813 , n70809 , n70812 );
nor ( n70814 , n25263 , n10547 );
xor ( n70815 , n70813 , n70814 );
and ( n70816 , n69621 , n69622 );
and ( n70817 , n69623 , n69626 );
or ( n70818 , n70816 , n70817 );
xor ( n70819 , n70815 , n70818 );
nor ( n70820 , n26317 , n9829 );
xor ( n70821 , n70819 , n70820 );
and ( n70822 , n69627 , n69628 );
and ( n70823 , n69629 , n69632 );
or ( n70824 , n70822 , n70823 );
xor ( n70825 , n70821 , n70824 );
nor ( n70826 , n27388 , n8955 );
xor ( n70827 , n70825 , n70826 );
and ( n70828 , n69633 , n69634 );
and ( n70829 , n69635 , n69638 );
or ( n70830 , n70828 , n70829 );
xor ( n70831 , n70827 , n70830 );
nor ( n70832 , n28478 , n603 );
xor ( n70833 , n70831 , n70832 );
and ( n70834 , n69639 , n69640 );
and ( n70835 , n69641 , n69644 );
or ( n70836 , n70834 , n70835 );
xor ( n70837 , n70833 , n70836 );
nor ( n70838 , n29587 , n652 );
xor ( n70839 , n70837 , n70838 );
and ( n70840 , n69645 , n69646 );
and ( n70841 , n69647 , n69650 );
or ( n70842 , n70840 , n70841 );
xor ( n70843 , n70839 , n70842 );
nor ( n70844 , n30716 , n624 );
xor ( n70845 , n70843 , n70844 );
and ( n70846 , n69651 , n69652 );
and ( n70847 , n69653 , n69656 );
or ( n70848 , n70846 , n70847 );
xor ( n70849 , n70845 , n70848 );
nor ( n70850 , n31858 , n648 );
xor ( n70851 , n70849 , n70850 );
and ( n70852 , n69657 , n69658 );
and ( n70853 , n69659 , n69662 );
or ( n70854 , n70852 , n70853 );
xor ( n70855 , n70851 , n70854 );
nor ( n70856 , n33024 , n686 );
xor ( n70857 , n70855 , n70856 );
and ( n70858 , n69663 , n69664 );
and ( n70859 , n69665 , n69668 );
or ( n70860 , n70858 , n70859 );
xor ( n70861 , n70857 , n70860 );
nor ( n70862 , n34215 , n735 );
xor ( n70863 , n70861 , n70862 );
and ( n70864 , n69669 , n69670 );
and ( n70865 , n69671 , n69674 );
or ( n70866 , n70864 , n70865 );
xor ( n70867 , n70863 , n70866 );
nor ( n70868 , n35410 , n798 );
xor ( n70869 , n70867 , n70868 );
and ( n70870 , n69675 , n69676 );
and ( n70871 , n69677 , n69680 );
or ( n70872 , n70870 , n70871 );
xor ( n70873 , n70869 , n70872 );
nor ( n70874 , n36611 , n870 );
xor ( n70875 , n70873 , n70874 );
and ( n70876 , n69681 , n69682 );
and ( n70877 , n69683 , n69686 );
or ( n70878 , n70876 , n70877 );
xor ( n70879 , n70875 , n70878 );
nor ( n70880 , n37816 , n960 );
xor ( n70881 , n70879 , n70880 );
and ( n70882 , n69687 , n69688 );
and ( n70883 , n69689 , n69692 );
or ( n70884 , n70882 , n70883 );
xor ( n70885 , n70881 , n70884 );
nor ( n70886 , n39018 , n1064 );
xor ( n70887 , n70885 , n70886 );
and ( n70888 , n69693 , n69694 );
and ( n70889 , n69695 , n69698 );
or ( n70890 , n70888 , n70889 );
xor ( n70891 , n70887 , n70890 );
nor ( n70892 , n40223 , n1178 );
xor ( n70893 , n70891 , n70892 );
and ( n70894 , n69699 , n69700 );
and ( n70895 , n69701 , n69704 );
or ( n70896 , n70894 , n70895 );
xor ( n70897 , n70893 , n70896 );
nor ( n70898 , n41428 , n1305 );
xor ( n70899 , n70897 , n70898 );
and ( n70900 , n69705 , n69706 );
and ( n70901 , n69707 , n69710 );
or ( n70902 , n70900 , n70901 );
xor ( n70903 , n70899 , n70902 );
nor ( n70904 , n42632 , n1447 );
xor ( n70905 , n70903 , n70904 );
and ( n70906 , n69711 , n69712 );
and ( n70907 , n69713 , n69716 );
or ( n70908 , n70906 , n70907 );
xor ( n70909 , n70905 , n70908 );
nor ( n70910 , n43834 , n1600 );
xor ( n70911 , n70909 , n70910 );
and ( n70912 , n69717 , n69718 );
and ( n70913 , n69719 , n69722 );
or ( n70914 , n70912 , n70913 );
xor ( n70915 , n70911 , n70914 );
nor ( n70916 , n45038 , n1768 );
xor ( n70917 , n70915 , n70916 );
and ( n70918 , n69723 , n69724 );
and ( n70919 , n69725 , n69728 );
or ( n70920 , n70918 , n70919 );
xor ( n70921 , n70917 , n70920 );
nor ( n70922 , n46239 , n1947 );
xor ( n70923 , n70921 , n70922 );
and ( n70924 , n69729 , n69730 );
and ( n70925 , n69731 , n69734 );
or ( n70926 , n70924 , n70925 );
xor ( n70927 , n70923 , n70926 );
nor ( n70928 , n47440 , n2139 );
xor ( n70929 , n70927 , n70928 );
and ( n70930 , n69735 , n69736 );
and ( n70931 , n69737 , n69740 );
or ( n70932 , n70930 , n70931 );
xor ( n70933 , n70929 , n70932 );
nor ( n70934 , n48641 , n2345 );
xor ( n70935 , n70933 , n70934 );
and ( n70936 , n69741 , n69742 );
and ( n70937 , n69743 , n69746 );
or ( n70938 , n70936 , n70937 );
xor ( n70939 , n70935 , n70938 );
nor ( n70940 , n49841 , n2568 );
xor ( n70941 , n70939 , n70940 );
and ( n70942 , n69747 , n69748 );
and ( n70943 , n69749 , n69752 );
or ( n70944 , n70942 , n70943 );
xor ( n70945 , n70941 , n70944 );
nor ( n70946 , n51040 , n2799 );
xor ( n70947 , n70945 , n70946 );
and ( n70948 , n69753 , n69754 );
and ( n70949 , n69755 , n69758 );
or ( n70950 , n70948 , n70949 );
xor ( n70951 , n70947 , n70950 );
nor ( n70952 , n52238 , n3045 );
xor ( n70953 , n70951 , n70952 );
and ( n70954 , n69759 , n69760 );
and ( n70955 , n69761 , n69764 );
or ( n70956 , n70954 , n70955 );
xor ( n70957 , n70953 , n70956 );
nor ( n70958 , n53432 , n3302 );
xor ( n70959 , n70957 , n70958 );
and ( n70960 , n69765 , n69766 );
and ( n70961 , n69767 , n69770 );
or ( n70962 , n70960 , n70961 );
xor ( n70963 , n70959 , n70962 );
nor ( n70964 , n54629 , n3572 );
xor ( n70965 , n70963 , n70964 );
and ( n70966 , n69771 , n69772 );
and ( n70967 , n69773 , n69776 );
or ( n70968 , n70966 , n70967 );
xor ( n70969 , n70965 , n70968 );
nor ( n70970 , n55826 , n3855 );
xor ( n70971 , n70969 , n70970 );
and ( n70972 , n69777 , n69778 );
and ( n70973 , n69779 , n69782 );
or ( n70974 , n70972 , n70973 );
xor ( n70975 , n70971 , n70974 );
nor ( n70976 , n57022 , n4153 );
xor ( n70977 , n70975 , n70976 );
and ( n70978 , n69783 , n69784 );
and ( n70979 , n69785 , n69788 );
or ( n70980 , n70978 , n70979 );
xor ( n70981 , n70977 , n70980 );
nor ( n70982 , n58217 , n4460 );
xor ( n70983 , n70981 , n70982 );
and ( n70984 , n69789 , n69790 );
and ( n70985 , n69791 , n69794 );
or ( n70986 , n70984 , n70985 );
xor ( n70987 , n70983 , n70986 );
nor ( n70988 , n59412 , n4788 );
xor ( n70989 , n70987 , n70988 );
and ( n70990 , n69795 , n69796 );
and ( n70991 , n69797 , n69800 );
or ( n70992 , n70990 , n70991 );
xor ( n70993 , n70989 , n70992 );
nor ( n70994 , n60600 , n5128 );
xor ( n70995 , n70993 , n70994 );
and ( n70996 , n69801 , n69802 );
and ( n70997 , n69803 , n69806 );
or ( n70998 , n70996 , n70997 );
xor ( n70999 , n70995 , n70998 );
nor ( n71000 , n61791 , n5479 );
xor ( n71001 , n70999 , n71000 );
and ( n71002 , n69807 , n69808 );
and ( n71003 , n69809 , n69812 );
or ( n71004 , n71002 , n71003 );
xor ( n71005 , n71001 , n71004 );
nor ( n71006 , n62982 , n5840 );
xor ( n71007 , n71005 , n71006 );
and ( n71008 , n69813 , n69814 );
and ( n71009 , n69815 , n69818 );
or ( n71010 , n71008 , n71009 );
xor ( n71011 , n71007 , n71010 );
nor ( n71012 , n64172 , n6214 );
xor ( n71013 , n71011 , n71012 );
and ( n71014 , n69819 , n69820 );
and ( n71015 , n69821 , n69824 );
or ( n71016 , n71014 , n71015 );
xor ( n71017 , n71013 , n71016 );
nor ( n71018 , n65360 , n6598 );
xor ( n71019 , n71017 , n71018 );
and ( n71020 , n69825 , n69826 );
and ( n71021 , n69827 , n69830 );
or ( n71022 , n71020 , n71021 );
xor ( n71023 , n71019 , n71022 );
nor ( n71024 , n66550 , n6999 );
xor ( n71025 , n71023 , n71024 );
and ( n71026 , n69831 , n69832 );
and ( n71027 , n69833 , n69836 );
or ( n71028 , n71026 , n71027 );
xor ( n71029 , n71025 , n71028 );
nor ( n71030 , n67736 , n7415 );
xor ( n71031 , n71029 , n71030 );
and ( n71032 , n69837 , n69838 );
and ( n71033 , n69839 , n69842 );
or ( n71034 , n71032 , n71033 );
xor ( n71035 , n71031 , n71034 );
nor ( n71036 , n68924 , n7843 );
xor ( n71037 , n71035 , n71036 );
and ( n71038 , n69843 , n69844 );
and ( n71039 , n69845 , n69848 );
or ( n71040 , n71038 , n71039 );
xor ( n71041 , n71037 , n71040 );
nor ( n71042 , n70110 , n8283 );
xor ( n71043 , n71041 , n71042 );
and ( n71044 , n69849 , n69850 );
and ( n71045 , n69851 , n69854 );
or ( n71046 , n71044 , n71045 );
xor ( n71047 , n71043 , n71046 );
and ( n71048 , n69867 , n69871 );
and ( n71049 , n69871 , n70096 );
and ( n71050 , n69867 , n70096 );
or ( n71051 , n71048 , n71049 , n71050 );
and ( n71052 , n33774 , n6504 );
not ( n71053 , n6504 );
nor ( n71054 , n71052 , n71053 );
xor ( n71055 , n71051 , n71054 );
and ( n71056 , n69877 , n69881 );
and ( n71057 , n69881 , n69949 );
and ( n71058 , n69877 , n69949 );
or ( n71059 , n71056 , n71057 , n71058 );
and ( n71060 , n69873 , n69950 );
and ( n71061 , n69950 , n70095 );
and ( n71062 , n69873 , n70095 );
or ( n71063 , n71060 , n71061 , n71062 );
xor ( n71064 , n71059 , n71063 );
and ( n71065 , n69979 , n70094 );
and ( n71066 , n69886 , n69890 );
and ( n71067 , n69890 , n69948 );
and ( n71068 , n69886 , n69948 );
or ( n71069 , n71066 , n71067 , n71068 );
and ( n71070 , n69983 , n70093 );
xor ( n71071 , n71069 , n71070 );
and ( n71072 , n69917 , n69921 );
and ( n71073 , n69921 , n69927 );
and ( n71074 , n69917 , n69927 );
or ( n71075 , n71072 , n71073 , n71074 );
and ( n71076 , n69895 , n69899 );
and ( n71077 , n69899 , n69947 );
and ( n71078 , n69895 , n69947 );
or ( n71079 , n71076 , n71077 , n71078 );
xor ( n71080 , n71075 , n71079 );
and ( n71081 , n69904 , n69908 );
and ( n71082 , n69908 , n69946 );
and ( n71083 , n69904 , n69946 );
or ( n71084 , n71081 , n71082 , n71083 );
and ( n71085 , n69991 , n70016 );
and ( n71086 , n70016 , n70054 );
and ( n71087 , n69991 , n70054 );
or ( n71088 , n71085 , n71086 , n71087 );
xor ( n71089 , n71084 , n71088 );
and ( n71090 , n69913 , n69928 );
and ( n71091 , n69928 , n69945 );
and ( n71092 , n69913 , n69945 );
or ( n71093 , n71090 , n71091 , n71092 );
and ( n71094 , n69995 , n69999 );
and ( n71095 , n69999 , n70015 );
and ( n71096 , n69995 , n70015 );
or ( n71097 , n71094 , n71095 , n71096 );
xor ( n71098 , n71093 , n71097 );
and ( n71099 , n69933 , n69938 );
and ( n71100 , n69938 , n69944 );
and ( n71101 , n69933 , n69944 );
or ( n71102 , n71099 , n71100 , n71101 );
and ( n71103 , n69923 , n69924 );
and ( n71104 , n69924 , n69926 );
and ( n71105 , n69923 , n69926 );
or ( n71106 , n71103 , n71104 , n71105 );
and ( n71107 , n69934 , n69935 );
and ( n71108 , n69935 , n69937 );
and ( n71109 , n69934 , n69937 );
or ( n71110 , n71107 , n71108 , n71109 );
xor ( n71111 , n71106 , n71110 );
and ( n71112 , n30695 , n7662 );
and ( n71113 , n31836 , n7310 );
xor ( n71114 , n71112 , n71113 );
and ( n71115 , n32649 , n6971 );
xor ( n71116 , n71114 , n71115 );
xor ( n71117 , n71111 , n71116 );
xor ( n71118 , n71102 , n71117 );
and ( n71119 , n69940 , n69941 );
and ( n71120 , n69941 , n69943 );
and ( n71121 , n69940 , n69943 );
or ( n71122 , n71119 , n71120 , n71121 );
and ( n71123 , n27361 , n9348 );
and ( n71124 , n28456 , n8669 );
xor ( n71125 , n71123 , n71124 );
and ( n71126 , n29559 , n8243 );
xor ( n71127 , n71125 , n71126 );
xor ( n71128 , n71122 , n71127 );
and ( n71129 , n24214 , n11718 );
and ( n71130 , n25243 , n10977 );
xor ( n71131 , n71129 , n71130 );
and ( n71132 , n26296 , n10239 );
xor ( n71133 , n71131 , n71132 );
xor ( n71134 , n71128 , n71133 );
xor ( n71135 , n71118 , n71134 );
xor ( n71136 , n71098 , n71135 );
xor ( n71137 , n71089 , n71136 );
xor ( n71138 , n71080 , n71137 );
xor ( n71139 , n71071 , n71138 );
xor ( n71140 , n71065 , n71139 );
and ( n71141 , n69958 , n69959 );
and ( n71142 , n69959 , n69961 );
and ( n71143 , n69958 , n69961 );
or ( n71144 , n71141 , n71142 , n71143 );
and ( n71145 , n69973 , n69974 );
and ( n71146 , n69974 , n69976 );
and ( n71147 , n69973 , n69976 );
or ( n71148 , n71145 , n71146 , n71147 );
xor ( n71149 , n71144 , n71148 );
and ( n71150 , n7385 , n31761 );
and ( n71151 , n7808 , n30629 );
xor ( n71152 , n71150 , n71151 );
and ( n71153 , n8079 , n29508 );
xor ( n71154 , n71152 , n71153 );
xor ( n71155 , n71149 , n71154 );
not ( n71156 , n6569 );
and ( n71157 , n34193 , n6569 );
nor ( n71158 , n71156 , n71157 );
and ( n71159 , n6816 , n32999 );
xor ( n71160 , n71158 , n71159 );
xor ( n71161 , n71155 , n71160 );
and ( n71162 , n69987 , n70055 );
and ( n71163 , n70055 , n70092 );
and ( n71164 , n69987 , n70092 );
or ( n71165 , n71162 , n71163 , n71164 );
and ( n71166 , n70060 , n70064 );
and ( n71167 , n70064 , n70091 );
and ( n71168 , n70060 , n70091 );
or ( n71169 , n71166 , n71167 , n71168 );
and ( n71170 , n70021 , n70037 );
and ( n71171 , n70037 , n70053 );
and ( n71172 , n70021 , n70053 );
or ( n71173 , n71170 , n71171 , n71172 );
and ( n71174 , n70004 , n70008 );
and ( n71175 , n70008 , n70014 );
and ( n71176 , n70004 , n70014 );
or ( n71177 , n71174 , n71175 , n71176 );
and ( n71178 , n70025 , n70030 );
and ( n71179 , n70030 , n70036 );
and ( n71180 , n70025 , n70036 );
or ( n71181 , n71178 , n71179 , n71180 );
xor ( n71182 , n71177 , n71181 );
and ( n71183 , n70010 , n70011 );
and ( n71184 , n70011 , n70013 );
and ( n71185 , n70010 , n70013 );
or ( n71186 , n71183 , n71184 , n71185 );
and ( n71187 , n70026 , n70027 );
and ( n71188 , n70027 , n70029 );
and ( n71189 , n70026 , n70029 );
or ( n71190 , n71187 , n71188 , n71189 );
xor ( n71191 , n71186 , n71190 );
and ( n71192 , n21216 , n14044 );
and ( n71193 , n22186 , n13256 );
xor ( n71194 , n71192 , n71193 );
and ( n71195 , n22892 , n12531 );
xor ( n71196 , n71194 , n71195 );
xor ( n71197 , n71191 , n71196 );
xor ( n71198 , n71182 , n71197 );
xor ( n71199 , n71173 , n71198 );
and ( n71200 , n70042 , n70046 );
and ( n71201 , n70046 , n70052 );
and ( n71202 , n70042 , n70052 );
or ( n71203 , n71200 , n71201 , n71202 );
and ( n71204 , n70032 , n70033 );
and ( n71205 , n70033 , n70035 );
and ( n71206 , n70032 , n70035 );
or ( n71207 , n71204 , n71205 , n71206 );
and ( n71208 , n18144 , n16550 );
and ( n71209 , n19324 , n15691 );
xor ( n71210 , n71208 , n71209 );
and ( n71211 , n20233 , n14838 );
xor ( n71212 , n71210 , n71211 );
xor ( n71213 , n71207 , n71212 );
and ( n71214 , n15758 , n19222 );
and ( n71215 , n16637 , n18407 );
xor ( n71216 , n71214 , n71215 );
buf ( n71217 , n17512 );
xor ( n71218 , n71216 , n71217 );
xor ( n71219 , n71213 , n71218 );
xor ( n71220 , n71203 , n71219 );
and ( n71221 , n70048 , n70049 );
and ( n71222 , n70049 , n70051 );
and ( n71223 , n70048 , n70051 );
or ( n71224 , n71221 , n71222 , n71223 );
and ( n71225 , n70079 , n70080 );
and ( n71226 , n70080 , n70082 );
and ( n71227 , n70079 , n70082 );
or ( n71228 , n71225 , n71226 , n71227 );
xor ( n71229 , n71224 , n71228 );
and ( n71230 , n13322 , n22065 );
and ( n71231 , n14118 , n20976 );
xor ( n71232 , n71230 , n71231 );
and ( n71233 , n14938 , n20156 );
xor ( n71234 , n71232 , n71233 );
xor ( n71235 , n71229 , n71234 );
xor ( n71236 , n71220 , n71235 );
xor ( n71237 , n71199 , n71236 );
xor ( n71238 , n71169 , n71237 );
and ( n71239 , n69955 , n69962 );
and ( n71240 , n69962 , n69978 );
and ( n71241 , n69955 , n69978 );
or ( n71242 , n71239 , n71240 , n71241 );
and ( n71243 , n70069 , n70073 );
and ( n71244 , n70073 , n70090 );
and ( n71245 , n70069 , n70090 );
or ( n71246 , n71243 , n71244 , n71245 );
xor ( n71247 , n71242 , n71246 );
and ( n71248 , n70078 , n70083 );
and ( n71249 , n70083 , n70089 );
and ( n71250 , n70078 , n70089 );
or ( n71251 , n71248 , n71249 , n71250 );
and ( n71252 , n69967 , n69971 );
and ( n71253 , n69971 , n69977 );
and ( n71254 , n69967 , n69977 );
or ( n71255 , n71252 , n71253 , n71254 );
xor ( n71256 , n71251 , n71255 );
and ( n71257 , n70085 , n70086 );
and ( n71258 , n70086 , n70088 );
and ( n71259 , n70085 , n70088 );
or ( n71260 , n71257 , n71258 , n71259 );
and ( n71261 , n11015 , n25163 );
and ( n71262 , n11769 , n24137 );
xor ( n71263 , n71261 , n71262 );
and ( n71264 , n12320 , n23075 );
xor ( n71265 , n71263 , n71264 );
xor ( n71266 , n71260 , n71265 );
and ( n71267 , n8718 , n28406 );
and ( n71268 , n9400 , n27296 );
xor ( n71269 , n71267 , n71268 );
and ( n71270 , n10291 , n26216 );
xor ( n71271 , n71269 , n71270 );
xor ( n71272 , n71266 , n71271 );
xor ( n71273 , n71256 , n71272 );
xor ( n71274 , n71247 , n71273 );
xor ( n71275 , n71238 , n71274 );
xor ( n71276 , n71165 , n71275 );
xor ( n71277 , n71161 , n71276 );
xor ( n71278 , n71140 , n71277 );
xor ( n71279 , n71064 , n71278 );
xor ( n71280 , n71055 , n71279 );
and ( n71281 , n69859 , n69862 );
and ( n71282 , n69862 , n70097 );
and ( n71283 , n69859 , n70097 );
or ( n71284 , n71281 , n71282 , n71283 );
xor ( n71285 , n71280 , n71284 );
and ( n71286 , n70098 , n70102 );
and ( n71287 , n70103 , n70106 );
or ( n71288 , n71286 , n71287 );
xor ( n71289 , n71285 , n71288 );
buf ( n71290 , n71289 );
buf ( n71291 , n71290 );
not ( n71292 , n71291 );
nor ( n71293 , n71292 , n8739 );
xor ( n71294 , n71047 , n71293 );
and ( n71295 , n69855 , n70111 );
and ( n71296 , n70112 , n70115 );
or ( n71297 , n71295 , n71296 );
xor ( n71298 , n71294 , n71297 );
buf ( n71299 , n71298 );
buf ( n71300 , n71299 );
not ( n71301 , n71300 );
buf ( n71302 , n593 );
not ( n71303 , n71302 );
nor ( n71304 , n71301 , n71303 );
xor ( n71305 , n70673 , n71304 );
xor ( n71306 , n70127 , n70670 );
nor ( n71307 , n70119 , n71303 );
and ( n71308 , n71306 , n71307 );
xor ( n71309 , n71306 , n71307 );
xor ( n71310 , n70131 , n70668 );
nor ( n71311 , n68933 , n71303 );
and ( n71312 , n71310 , n71311 );
xor ( n71313 , n71310 , n71311 );
xor ( n71314 , n70135 , n70666 );
nor ( n71315 , n67745 , n71303 );
and ( n71316 , n71314 , n71315 );
xor ( n71317 , n71314 , n71315 );
xor ( n71318 , n70139 , n70664 );
nor ( n71319 , n66559 , n71303 );
and ( n71320 , n71318 , n71319 );
xor ( n71321 , n71318 , n71319 );
xor ( n71322 , n70143 , n70662 );
nor ( n71323 , n65369 , n71303 );
and ( n71324 , n71322 , n71323 );
xor ( n71325 , n71322 , n71323 );
xor ( n71326 , n70147 , n70660 );
nor ( n71327 , n64181 , n71303 );
and ( n71328 , n71326 , n71327 );
xor ( n71329 , n71326 , n71327 );
xor ( n71330 , n70151 , n70658 );
nor ( n71331 , n62991 , n71303 );
and ( n71332 , n71330 , n71331 );
xor ( n71333 , n71330 , n71331 );
xor ( n71334 , n70155 , n70656 );
nor ( n71335 , n61800 , n71303 );
and ( n71336 , n71334 , n71335 );
xor ( n71337 , n71334 , n71335 );
xor ( n71338 , n70159 , n70654 );
nor ( n71339 , n60609 , n71303 );
and ( n71340 , n71338 , n71339 );
xor ( n71341 , n71338 , n71339 );
xor ( n71342 , n70163 , n70652 );
nor ( n71343 , n59421 , n71303 );
and ( n71344 , n71342 , n71343 );
xor ( n71345 , n71342 , n71343 );
xor ( n71346 , n70167 , n70650 );
nor ( n71347 , n58226 , n71303 );
and ( n71348 , n71346 , n71347 );
xor ( n71349 , n71346 , n71347 );
xor ( n71350 , n70171 , n70648 );
nor ( n71351 , n57031 , n71303 );
and ( n71352 , n71350 , n71351 );
xor ( n71353 , n71350 , n71351 );
xor ( n71354 , n70175 , n70646 );
nor ( n71355 , n55835 , n71303 );
and ( n71356 , n71354 , n71355 );
xor ( n71357 , n71354 , n71355 );
xor ( n71358 , n70179 , n70644 );
nor ( n71359 , n54638 , n71303 );
and ( n71360 , n71358 , n71359 );
xor ( n71361 , n71358 , n71359 );
xor ( n71362 , n70183 , n70642 );
nor ( n71363 , n53441 , n71303 );
and ( n71364 , n71362 , n71363 );
xor ( n71365 , n71362 , n71363 );
xor ( n71366 , n70187 , n70640 );
nor ( n71367 , n52247 , n71303 );
and ( n71368 , n71366 , n71367 );
xor ( n71369 , n71366 , n71367 );
xor ( n71370 , n70191 , n70638 );
nor ( n71371 , n51049 , n71303 );
and ( n71372 , n71370 , n71371 );
xor ( n71373 , n71370 , n71371 );
xor ( n71374 , n70195 , n70636 );
nor ( n71375 , n49850 , n71303 );
and ( n71376 , n71374 , n71375 );
xor ( n71377 , n71374 , n71375 );
xor ( n71378 , n70199 , n70634 );
nor ( n71379 , n48650 , n71303 );
and ( n71380 , n71378 , n71379 );
xor ( n71381 , n71378 , n71379 );
xor ( n71382 , n70203 , n70632 );
nor ( n71383 , n47449 , n71303 );
and ( n71384 , n71382 , n71383 );
xor ( n71385 , n71382 , n71383 );
xor ( n71386 , n70207 , n70630 );
nor ( n71387 , n46248 , n71303 );
and ( n71388 , n71386 , n71387 );
xor ( n71389 , n71386 , n71387 );
xor ( n71390 , n70211 , n70628 );
nor ( n71391 , n45047 , n71303 );
and ( n71392 , n71390 , n71391 );
xor ( n71393 , n71390 , n71391 );
xor ( n71394 , n70215 , n70626 );
nor ( n71395 , n43843 , n71303 );
and ( n71396 , n71394 , n71395 );
xor ( n71397 , n71394 , n71395 );
xor ( n71398 , n70219 , n70624 );
nor ( n71399 , n42641 , n71303 );
and ( n71400 , n71398 , n71399 );
xor ( n71401 , n71398 , n71399 );
xor ( n71402 , n70223 , n70622 );
nor ( n71403 , n41437 , n71303 );
and ( n71404 , n71402 , n71403 );
xor ( n71405 , n71402 , n71403 );
xor ( n71406 , n70227 , n70620 );
nor ( n71407 , n40232 , n71303 );
and ( n71408 , n71406 , n71407 );
xor ( n71409 , n71406 , n71407 );
xor ( n71410 , n70231 , n70618 );
nor ( n71411 , n39027 , n71303 );
and ( n71412 , n71410 , n71411 );
xor ( n71413 , n71410 , n71411 );
xor ( n71414 , n70235 , n70616 );
nor ( n71415 , n37825 , n71303 );
and ( n71416 , n71414 , n71415 );
xor ( n71417 , n71414 , n71415 );
xor ( n71418 , n70239 , n70614 );
nor ( n71419 , n36620 , n71303 );
and ( n71420 , n71418 , n71419 );
xor ( n71421 , n71418 , n71419 );
xor ( n71422 , n70243 , n70612 );
nor ( n71423 , n35419 , n71303 );
and ( n71424 , n71422 , n71423 );
xor ( n71425 , n71422 , n71423 );
xor ( n71426 , n70247 , n70610 );
nor ( n71427 , n34224 , n71303 );
and ( n71428 , n71426 , n71427 );
xor ( n71429 , n71426 , n71427 );
xor ( n71430 , n70251 , n70608 );
nor ( n71431 , n33033 , n71303 );
and ( n71432 , n71430 , n71431 );
xor ( n71433 , n71430 , n71431 );
xor ( n71434 , n70255 , n70606 );
nor ( n71435 , n31867 , n71303 );
and ( n71436 , n71434 , n71435 );
xor ( n71437 , n71434 , n71435 );
xor ( n71438 , n70259 , n70604 );
nor ( n71439 , n30725 , n71303 );
and ( n71440 , n71438 , n71439 );
xor ( n71441 , n71438 , n71439 );
xor ( n71442 , n70263 , n70602 );
nor ( n71443 , n29596 , n71303 );
and ( n71444 , n71442 , n71443 );
xor ( n71445 , n71442 , n71443 );
xor ( n71446 , n70267 , n70600 );
nor ( n71447 , n28487 , n71303 );
and ( n71448 , n71446 , n71447 );
xor ( n71449 , n71446 , n71447 );
xor ( n71450 , n70271 , n70598 );
nor ( n71451 , n27397 , n71303 );
and ( n71452 , n71450 , n71451 );
xor ( n71453 , n71450 , n71451 );
xor ( n71454 , n70275 , n70596 );
nor ( n71455 , n26326 , n71303 );
and ( n71456 , n71454 , n71455 );
xor ( n71457 , n71454 , n71455 );
xor ( n71458 , n70279 , n70594 );
nor ( n71459 , n25272 , n71303 );
and ( n71460 , n71458 , n71459 );
xor ( n71461 , n71458 , n71459 );
xor ( n71462 , n70283 , n70592 );
nor ( n71463 , n24242 , n71303 );
and ( n71464 , n71462 , n71463 );
xor ( n71465 , n71462 , n71463 );
xor ( n71466 , n70287 , n70590 );
nor ( n71467 , n23225 , n71303 );
and ( n71468 , n71466 , n71467 );
xor ( n71469 , n71466 , n71467 );
xor ( n71470 , n70291 , n70588 );
nor ( n71471 , n22231 , n71303 );
and ( n71472 , n71470 , n71471 );
xor ( n71473 , n71470 , n71471 );
xor ( n71474 , n70295 , n70586 );
nor ( n71475 , n21258 , n71303 );
and ( n71476 , n71474 , n71475 );
xor ( n71477 , n71474 , n71475 );
xor ( n71478 , n70299 , n70584 );
nor ( n71479 , n20303 , n71303 );
and ( n71480 , n71478 , n71479 );
xor ( n71481 , n71478 , n71479 );
xor ( n71482 , n70303 , n70582 );
nor ( n71483 , n19365 , n71303 );
and ( n71484 , n71482 , n71483 );
xor ( n71485 , n71482 , n71483 );
xor ( n71486 , n70307 , n70580 );
nor ( n71487 , n18448 , n71303 );
and ( n71488 , n71486 , n71487 );
xor ( n71489 , n71486 , n71487 );
xor ( n71490 , n70311 , n70578 );
nor ( n71491 , n17548 , n71303 );
and ( n71492 , n71490 , n71491 );
xor ( n71493 , n71490 , n71491 );
xor ( n71494 , n70315 , n70576 );
nor ( n71495 , n16669 , n71303 );
and ( n71496 , n71494 , n71495 );
xor ( n71497 , n71494 , n71495 );
xor ( n71498 , n70319 , n70574 );
nor ( n71499 , n15809 , n71303 );
and ( n71500 , n71498 , n71499 );
xor ( n71501 , n71498 , n71499 );
xor ( n71502 , n70323 , n70572 );
nor ( n71503 , n14968 , n71303 );
and ( n71504 , n71502 , n71503 );
xor ( n71505 , n71502 , n71503 );
xor ( n71506 , n70327 , n70570 );
nor ( n71507 , n14147 , n71303 );
and ( n71508 , n71506 , n71507 );
xor ( n71509 , n71506 , n71507 );
xor ( n71510 , n70331 , n70568 );
nor ( n71511 , n13349 , n71303 );
and ( n71512 , n71510 , n71511 );
xor ( n71513 , n71510 , n71511 );
xor ( n71514 , n70335 , n70566 );
nor ( n71515 , n12564 , n71303 );
and ( n71516 , n71514 , n71515 );
xor ( n71517 , n71514 , n71515 );
xor ( n71518 , n70339 , n70564 );
nor ( n71519 , n11799 , n71303 );
and ( n71520 , n71518 , n71519 );
xor ( n71521 , n71518 , n71519 );
xor ( n71522 , n70343 , n70562 );
nor ( n71523 , n11050 , n71303 );
and ( n71524 , n71522 , n71523 );
xor ( n71525 , n71522 , n71523 );
xor ( n71526 , n70347 , n70560 );
nor ( n71527 , n10321 , n71303 );
and ( n71528 , n71526 , n71527 );
xor ( n71529 , n71526 , n71527 );
xor ( n71530 , n70351 , n70558 );
nor ( n71531 , n9429 , n71303 );
and ( n71532 , n71530 , n71531 );
xor ( n71533 , n71530 , n71531 );
xor ( n71534 , n70355 , n70556 );
nor ( n71535 , n8949 , n71303 );
and ( n71536 , n71534 , n71535 );
xor ( n71537 , n71534 , n71535 );
xor ( n71538 , n70359 , n70554 );
nor ( n71539 , n9437 , n71303 );
and ( n71540 , n71538 , n71539 );
xor ( n71541 , n71538 , n71539 );
xor ( n71542 , n70363 , n70552 );
nor ( n71543 , n9446 , n71303 );
and ( n71544 , n71542 , n71543 );
xor ( n71545 , n71542 , n71543 );
xor ( n71546 , n70367 , n70550 );
nor ( n71547 , n9455 , n71303 );
and ( n71548 , n71546 , n71547 );
xor ( n71549 , n71546 , n71547 );
xor ( n71550 , n70371 , n70548 );
nor ( n71551 , n9464 , n71303 );
and ( n71552 , n71550 , n71551 );
xor ( n71553 , n71550 , n71551 );
xor ( n71554 , n70375 , n70546 );
nor ( n71555 , n9473 , n71303 );
and ( n71556 , n71554 , n71555 );
xor ( n71557 , n71554 , n71555 );
xor ( n71558 , n70379 , n70544 );
nor ( n71559 , n9482 , n71303 );
and ( n71560 , n71558 , n71559 );
xor ( n71561 , n71558 , n71559 );
xor ( n71562 , n70383 , n70542 );
nor ( n71563 , n9491 , n71303 );
and ( n71564 , n71562 , n71563 );
xor ( n71565 , n71562 , n71563 );
xor ( n71566 , n70387 , n70540 );
nor ( n71567 , n9500 , n71303 );
and ( n71568 , n71566 , n71567 );
xor ( n71569 , n71566 , n71567 );
xor ( n71570 , n70391 , n70538 );
nor ( n71571 , n9509 , n71303 );
and ( n71572 , n71570 , n71571 );
xor ( n71573 , n71570 , n71571 );
xor ( n71574 , n70395 , n70536 );
nor ( n71575 , n9518 , n71303 );
and ( n71576 , n71574 , n71575 );
xor ( n71577 , n71574 , n71575 );
xor ( n71578 , n70399 , n70534 );
nor ( n71579 , n9527 , n71303 );
and ( n71580 , n71578 , n71579 );
xor ( n71581 , n71578 , n71579 );
xor ( n71582 , n70403 , n70532 );
nor ( n71583 , n9536 , n71303 );
and ( n71584 , n71582 , n71583 );
xor ( n71585 , n71582 , n71583 );
xor ( n71586 , n70407 , n70530 );
nor ( n71587 , n9545 , n71303 );
and ( n71588 , n71586 , n71587 );
xor ( n71589 , n71586 , n71587 );
xor ( n71590 , n70411 , n70528 );
nor ( n71591 , n9554 , n71303 );
and ( n71592 , n71590 , n71591 );
xor ( n71593 , n71590 , n71591 );
xor ( n71594 , n70415 , n70526 );
nor ( n71595 , n9563 , n71303 );
and ( n71596 , n71594 , n71595 );
xor ( n71597 , n71594 , n71595 );
xor ( n71598 , n70419 , n70524 );
nor ( n71599 , n9572 , n71303 );
and ( n71600 , n71598 , n71599 );
xor ( n71601 , n71598 , n71599 );
xor ( n71602 , n70423 , n70522 );
nor ( n71603 , n9581 , n71303 );
and ( n71604 , n71602 , n71603 );
xor ( n71605 , n71602 , n71603 );
xor ( n71606 , n70427 , n70520 );
nor ( n71607 , n9590 , n71303 );
and ( n71608 , n71606 , n71607 );
xor ( n71609 , n71606 , n71607 );
xor ( n71610 , n70431 , n70518 );
nor ( n71611 , n9599 , n71303 );
and ( n71612 , n71610 , n71611 );
xor ( n71613 , n71610 , n71611 );
xor ( n71614 , n70435 , n70516 );
nor ( n71615 , n9608 , n71303 );
and ( n71616 , n71614 , n71615 );
xor ( n71617 , n71614 , n71615 );
xor ( n71618 , n70439 , n70514 );
nor ( n71619 , n9617 , n71303 );
and ( n71620 , n71618 , n71619 );
xor ( n71621 , n71618 , n71619 );
xor ( n71622 , n70443 , n70512 );
nor ( n71623 , n9626 , n71303 );
and ( n71624 , n71622 , n71623 );
xor ( n71625 , n71622 , n71623 );
xor ( n71626 , n70447 , n70510 );
nor ( n71627 , n9635 , n71303 );
and ( n71628 , n71626 , n71627 );
xor ( n71629 , n71626 , n71627 );
xor ( n71630 , n70451 , n70508 );
nor ( n71631 , n9644 , n71303 );
and ( n71632 , n71630 , n71631 );
xor ( n71633 , n71630 , n71631 );
xor ( n71634 , n70455 , n70506 );
nor ( n71635 , n9653 , n71303 );
and ( n71636 , n71634 , n71635 );
xor ( n71637 , n71634 , n71635 );
xor ( n71638 , n70459 , n70504 );
nor ( n71639 , n9662 , n71303 );
and ( n71640 , n71638 , n71639 );
xor ( n71641 , n71638 , n71639 );
xor ( n71642 , n70463 , n70502 );
nor ( n71643 , n9671 , n71303 );
and ( n71644 , n71642 , n71643 );
xor ( n71645 , n71642 , n71643 );
xor ( n71646 , n70467 , n70500 );
nor ( n71647 , n9680 , n71303 );
and ( n71648 , n71646 , n71647 );
xor ( n71649 , n71646 , n71647 );
xor ( n71650 , n70471 , n70498 );
nor ( n71651 , n9689 , n71303 );
and ( n71652 , n71650 , n71651 );
xor ( n71653 , n71650 , n71651 );
xor ( n71654 , n70475 , n70496 );
nor ( n71655 , n9698 , n71303 );
and ( n71656 , n71654 , n71655 );
xor ( n71657 , n71654 , n71655 );
xor ( n71658 , n70479 , n70494 );
nor ( n71659 , n9707 , n71303 );
and ( n71660 , n71658 , n71659 );
xor ( n71661 , n71658 , n71659 );
xor ( n71662 , n70483 , n70492 );
nor ( n71663 , n9716 , n71303 );
and ( n71664 , n71662 , n71663 );
xor ( n71665 , n71662 , n71663 );
xor ( n71666 , n70487 , n70490 );
nor ( n71667 , n9725 , n71303 );
and ( n71668 , n71666 , n71667 );
xor ( n71669 , n71666 , n71667 );
xor ( n71670 , n70488 , n70489 );
nor ( n71671 , n9734 , n71303 );
and ( n71672 , n71670 , n71671 );
xor ( n71673 , n71670 , n71671 );
nor ( n71674 , n9752 , n70121 );
nor ( n71675 , n9743 , n71303 );
and ( n71676 , n71674 , n71675 );
and ( n71677 , n71673 , n71676 );
or ( n71678 , n71672 , n71677 );
and ( n71679 , n71669 , n71678 );
or ( n71680 , n71668 , n71679 );
and ( n71681 , n71665 , n71680 );
or ( n71682 , n71664 , n71681 );
and ( n71683 , n71661 , n71682 );
or ( n71684 , n71660 , n71683 );
and ( n71685 , n71657 , n71684 );
or ( n71686 , n71656 , n71685 );
and ( n71687 , n71653 , n71686 );
or ( n71688 , n71652 , n71687 );
and ( n71689 , n71649 , n71688 );
or ( n71690 , n71648 , n71689 );
and ( n71691 , n71645 , n71690 );
or ( n71692 , n71644 , n71691 );
and ( n71693 , n71641 , n71692 );
or ( n71694 , n71640 , n71693 );
and ( n71695 , n71637 , n71694 );
or ( n71696 , n71636 , n71695 );
and ( n71697 , n71633 , n71696 );
or ( n71698 , n71632 , n71697 );
and ( n71699 , n71629 , n71698 );
or ( n71700 , n71628 , n71699 );
and ( n71701 , n71625 , n71700 );
or ( n71702 , n71624 , n71701 );
and ( n71703 , n71621 , n71702 );
or ( n71704 , n71620 , n71703 );
and ( n71705 , n71617 , n71704 );
or ( n71706 , n71616 , n71705 );
and ( n71707 , n71613 , n71706 );
or ( n71708 , n71612 , n71707 );
and ( n71709 , n71609 , n71708 );
or ( n71710 , n71608 , n71709 );
and ( n71711 , n71605 , n71710 );
or ( n71712 , n71604 , n71711 );
and ( n71713 , n71601 , n71712 );
or ( n71714 , n71600 , n71713 );
and ( n71715 , n71597 , n71714 );
or ( n71716 , n71596 , n71715 );
and ( n71717 , n71593 , n71716 );
or ( n71718 , n71592 , n71717 );
and ( n71719 , n71589 , n71718 );
or ( n71720 , n71588 , n71719 );
and ( n71721 , n71585 , n71720 );
or ( n71722 , n71584 , n71721 );
and ( n71723 , n71581 , n71722 );
or ( n71724 , n71580 , n71723 );
and ( n71725 , n71577 , n71724 );
or ( n71726 , n71576 , n71725 );
and ( n71727 , n71573 , n71726 );
or ( n71728 , n71572 , n71727 );
and ( n71729 , n71569 , n71728 );
or ( n71730 , n71568 , n71729 );
and ( n71731 , n71565 , n71730 );
or ( n71732 , n71564 , n71731 );
and ( n71733 , n71561 , n71732 );
or ( n71734 , n71560 , n71733 );
and ( n71735 , n71557 , n71734 );
or ( n71736 , n71556 , n71735 );
and ( n71737 , n71553 , n71736 );
or ( n71738 , n71552 , n71737 );
and ( n71739 , n71549 , n71738 );
or ( n71740 , n71548 , n71739 );
and ( n71741 , n71545 , n71740 );
or ( n71742 , n71544 , n71741 );
and ( n71743 , n71541 , n71742 );
or ( n71744 , n71540 , n71743 );
and ( n71745 , n71537 , n71744 );
or ( n71746 , n71536 , n71745 );
and ( n71747 , n71533 , n71746 );
or ( n71748 , n71532 , n71747 );
and ( n71749 , n71529 , n71748 );
or ( n71750 , n71528 , n71749 );
and ( n71751 , n71525 , n71750 );
or ( n71752 , n71524 , n71751 );
and ( n71753 , n71521 , n71752 );
or ( n71754 , n71520 , n71753 );
and ( n71755 , n71517 , n71754 );
or ( n71756 , n71516 , n71755 );
and ( n71757 , n71513 , n71756 );
or ( n71758 , n71512 , n71757 );
and ( n71759 , n71509 , n71758 );
or ( n71760 , n71508 , n71759 );
and ( n71761 , n71505 , n71760 );
or ( n71762 , n71504 , n71761 );
and ( n71763 , n71501 , n71762 );
or ( n71764 , n71500 , n71763 );
and ( n71765 , n71497 , n71764 );
or ( n71766 , n71496 , n71765 );
and ( n71767 , n71493 , n71766 );
or ( n71768 , n71492 , n71767 );
and ( n71769 , n71489 , n71768 );
or ( n71770 , n71488 , n71769 );
and ( n71771 , n71485 , n71770 );
or ( n71772 , n71484 , n71771 );
and ( n71773 , n71481 , n71772 );
or ( n71774 , n71480 , n71773 );
and ( n71775 , n71477 , n71774 );
or ( n71776 , n71476 , n71775 );
and ( n71777 , n71473 , n71776 );
or ( n71778 , n71472 , n71777 );
and ( n71779 , n71469 , n71778 );
or ( n71780 , n71468 , n71779 );
and ( n71781 , n71465 , n71780 );
or ( n71782 , n71464 , n71781 );
and ( n71783 , n71461 , n71782 );
or ( n71784 , n71460 , n71783 );
and ( n71785 , n71457 , n71784 );
or ( n71786 , n71456 , n71785 );
and ( n71787 , n71453 , n71786 );
or ( n71788 , n71452 , n71787 );
and ( n71789 , n71449 , n71788 );
or ( n71790 , n71448 , n71789 );
and ( n71791 , n71445 , n71790 );
or ( n71792 , n71444 , n71791 );
and ( n71793 , n71441 , n71792 );
or ( n71794 , n71440 , n71793 );
and ( n71795 , n71437 , n71794 );
or ( n71796 , n71436 , n71795 );
and ( n71797 , n71433 , n71796 );
or ( n71798 , n71432 , n71797 );
and ( n71799 , n71429 , n71798 );
or ( n71800 , n71428 , n71799 );
and ( n71801 , n71425 , n71800 );
or ( n71802 , n71424 , n71801 );
and ( n71803 , n71421 , n71802 );
or ( n71804 , n71420 , n71803 );
and ( n71805 , n71417 , n71804 );
or ( n71806 , n71416 , n71805 );
and ( n71807 , n71413 , n71806 );
or ( n71808 , n71412 , n71807 );
and ( n71809 , n71409 , n71808 );
or ( n71810 , n71408 , n71809 );
and ( n71811 , n71405 , n71810 );
or ( n71812 , n71404 , n71811 );
and ( n71813 , n71401 , n71812 );
or ( n71814 , n71400 , n71813 );
and ( n71815 , n71397 , n71814 );
or ( n71816 , n71396 , n71815 );
and ( n71817 , n71393 , n71816 );
or ( n71818 , n71392 , n71817 );
and ( n71819 , n71389 , n71818 );
or ( n71820 , n71388 , n71819 );
and ( n71821 , n71385 , n71820 );
or ( n71822 , n71384 , n71821 );
and ( n71823 , n71381 , n71822 );
or ( n71824 , n71380 , n71823 );
and ( n71825 , n71377 , n71824 );
or ( n71826 , n71376 , n71825 );
and ( n71827 , n71373 , n71826 );
or ( n71828 , n71372 , n71827 );
and ( n71829 , n71369 , n71828 );
or ( n71830 , n71368 , n71829 );
and ( n71831 , n71365 , n71830 );
or ( n71832 , n71364 , n71831 );
and ( n71833 , n71361 , n71832 );
or ( n71834 , n71360 , n71833 );
and ( n71835 , n71357 , n71834 );
or ( n71836 , n71356 , n71835 );
and ( n71837 , n71353 , n71836 );
or ( n71838 , n71352 , n71837 );
and ( n71839 , n71349 , n71838 );
or ( n71840 , n71348 , n71839 );
and ( n71841 , n71345 , n71840 );
or ( n71842 , n71344 , n71841 );
and ( n71843 , n71341 , n71842 );
or ( n71844 , n71340 , n71843 );
and ( n71845 , n71337 , n71844 );
or ( n71846 , n71336 , n71845 );
and ( n71847 , n71333 , n71846 );
or ( n71848 , n71332 , n71847 );
and ( n71849 , n71329 , n71848 );
or ( n71850 , n71328 , n71849 );
and ( n71851 , n71325 , n71850 );
or ( n71852 , n71324 , n71851 );
and ( n71853 , n71321 , n71852 );
or ( n71854 , n71320 , n71853 );
and ( n71855 , n71317 , n71854 );
or ( n71856 , n71316 , n71855 );
and ( n71857 , n71313 , n71856 );
or ( n71858 , n71312 , n71857 );
and ( n71859 , n71309 , n71858 );
or ( n71860 , n71308 , n71859 );
xor ( n71861 , n71305 , n71860 );
and ( n71862 , n33403 , n6996 );
nor ( n71863 , n6997 , n71862 );
nor ( n71864 , n7413 , n32231 );
xor ( n71865 , n71863 , n71864 );
and ( n71866 , n70675 , n70676 );
and ( n71867 , n70677 , n70680 );
or ( n71868 , n71866 , n71867 );
xor ( n71869 , n71865 , n71868 );
nor ( n71870 , n7841 , n31083 );
xor ( n71871 , n71869 , n71870 );
and ( n71872 , n70681 , n70682 );
and ( n71873 , n70683 , n70686 );
or ( n71874 , n71872 , n71873 );
xor ( n71875 , n71871 , n71874 );
nor ( n71876 , n8281 , n29948 );
xor ( n71877 , n71875 , n71876 );
and ( n71878 , n70687 , n70688 );
and ( n71879 , n70689 , n70692 );
or ( n71880 , n71878 , n71879 );
xor ( n71881 , n71877 , n71880 );
nor ( n71882 , n8737 , n28833 );
xor ( n71883 , n71881 , n71882 );
and ( n71884 , n70693 , n70694 );
and ( n71885 , n70695 , n70698 );
or ( n71886 , n71884 , n71885 );
xor ( n71887 , n71883 , n71886 );
nor ( n71888 , n9420 , n27737 );
xor ( n71889 , n71887 , n71888 );
and ( n71890 , n70699 , n70700 );
and ( n71891 , n70701 , n70704 );
or ( n71892 , n71890 , n71891 );
xor ( n71893 , n71889 , n71892 );
nor ( n71894 , n10312 , n26660 );
xor ( n71895 , n71893 , n71894 );
and ( n71896 , n70705 , n70706 );
and ( n71897 , n70707 , n70710 );
or ( n71898 , n71896 , n71897 );
xor ( n71899 , n71895 , n71898 );
nor ( n71900 , n11041 , n25600 );
xor ( n71901 , n71899 , n71900 );
and ( n71902 , n70711 , n70712 );
and ( n71903 , n70713 , n70716 );
or ( n71904 , n71902 , n71903 );
xor ( n71905 , n71901 , n71904 );
nor ( n71906 , n11790 , n24564 );
xor ( n71907 , n71905 , n71906 );
and ( n71908 , n70717 , n70718 );
and ( n71909 , n70719 , n70722 );
or ( n71910 , n71908 , n71909 );
xor ( n71911 , n71907 , n71910 );
nor ( n71912 , n12555 , n23541 );
xor ( n71913 , n71911 , n71912 );
and ( n71914 , n70723 , n70724 );
and ( n71915 , n70725 , n70728 );
or ( n71916 , n71914 , n71915 );
xor ( n71917 , n71913 , n71916 );
nor ( n71918 , n13340 , n22541 );
xor ( n71919 , n71917 , n71918 );
and ( n71920 , n70729 , n70730 );
and ( n71921 , n70731 , n70734 );
or ( n71922 , n71920 , n71921 );
xor ( n71923 , n71919 , n71922 );
nor ( n71924 , n14138 , n21562 );
xor ( n71925 , n71923 , n71924 );
and ( n71926 , n70735 , n70736 );
and ( n71927 , n70737 , n70740 );
or ( n71928 , n71926 , n71927 );
xor ( n71929 , n71925 , n71928 );
nor ( n71930 , n14959 , n20601 );
xor ( n71931 , n71929 , n71930 );
and ( n71932 , n70741 , n70742 );
and ( n71933 , n70743 , n70746 );
or ( n71934 , n71932 , n71933 );
xor ( n71935 , n71931 , n71934 );
nor ( n71936 , n15800 , n19657 );
xor ( n71937 , n71935 , n71936 );
and ( n71938 , n70747 , n70748 );
and ( n71939 , n70749 , n70752 );
or ( n71940 , n71938 , n71939 );
xor ( n71941 , n71937 , n71940 );
nor ( n71942 , n16660 , n18734 );
xor ( n71943 , n71941 , n71942 );
and ( n71944 , n70753 , n70754 );
and ( n71945 , n70755 , n70758 );
or ( n71946 , n71944 , n71945 );
xor ( n71947 , n71943 , n71946 );
nor ( n71948 , n17539 , n17828 );
xor ( n71949 , n71947 , n71948 );
and ( n71950 , n70759 , n70760 );
and ( n71951 , n70761 , n70764 );
or ( n71952 , n71950 , n71951 );
xor ( n71953 , n71949 , n71952 );
nor ( n71954 , n18439 , n16943 );
xor ( n71955 , n71953 , n71954 );
and ( n71956 , n70765 , n70766 );
and ( n71957 , n70767 , n70770 );
or ( n71958 , n71956 , n71957 );
xor ( n71959 , n71955 , n71958 );
nor ( n71960 , n19356 , n16077 );
xor ( n71961 , n71959 , n71960 );
and ( n71962 , n70771 , n70772 );
and ( n71963 , n70773 , n70776 );
or ( n71964 , n71962 , n71963 );
xor ( n71965 , n71961 , n71964 );
nor ( n71966 , n20294 , n15230 );
xor ( n71967 , n71965 , n71966 );
and ( n71968 , n70777 , n70778 );
and ( n71969 , n70779 , n70782 );
or ( n71970 , n71968 , n71969 );
xor ( n71971 , n71967 , n71970 );
nor ( n71972 , n21249 , n14403 );
xor ( n71973 , n71971 , n71972 );
and ( n71974 , n70783 , n70784 );
and ( n71975 , n70785 , n70788 );
or ( n71976 , n71974 , n71975 );
xor ( n71977 , n71973 , n71976 );
nor ( n71978 , n22222 , n13599 );
xor ( n71979 , n71977 , n71978 );
and ( n71980 , n70789 , n70790 );
and ( n71981 , n70791 , n70794 );
or ( n71982 , n71980 , n71981 );
xor ( n71983 , n71979 , n71982 );
nor ( n71984 , n23216 , n12808 );
xor ( n71985 , n71983 , n71984 );
and ( n71986 , n70795 , n70796 );
and ( n71987 , n70797 , n70800 );
or ( n71988 , n71986 , n71987 );
xor ( n71989 , n71985 , n71988 );
nor ( n71990 , n24233 , n12037 );
xor ( n71991 , n71989 , n71990 );
and ( n71992 , n70801 , n70802 );
and ( n71993 , n70803 , n70806 );
or ( n71994 , n71992 , n71993 );
xor ( n71995 , n71991 , n71994 );
nor ( n71996 , n25263 , n11282 );
xor ( n71997 , n71995 , n71996 );
and ( n71998 , n70807 , n70808 );
and ( n71999 , n70809 , n70812 );
or ( n72000 , n71998 , n71999 );
xor ( n72001 , n71997 , n72000 );
nor ( n72002 , n26317 , n10547 );
xor ( n72003 , n72001 , n72002 );
and ( n72004 , n70813 , n70814 );
and ( n72005 , n70815 , n70818 );
or ( n72006 , n72004 , n72005 );
xor ( n72007 , n72003 , n72006 );
nor ( n72008 , n27388 , n9829 );
xor ( n72009 , n72007 , n72008 );
and ( n72010 , n70819 , n70820 );
and ( n72011 , n70821 , n70824 );
or ( n72012 , n72010 , n72011 );
xor ( n72013 , n72009 , n72012 );
nor ( n72014 , n28478 , n8955 );
xor ( n72015 , n72013 , n72014 );
and ( n72016 , n70825 , n70826 );
and ( n72017 , n70827 , n70830 );
or ( n72018 , n72016 , n72017 );
xor ( n72019 , n72015 , n72018 );
nor ( n72020 , n29587 , n603 );
xor ( n72021 , n72019 , n72020 );
and ( n72022 , n70831 , n70832 );
and ( n72023 , n70833 , n70836 );
or ( n72024 , n72022 , n72023 );
xor ( n72025 , n72021 , n72024 );
nor ( n72026 , n30716 , n652 );
xor ( n72027 , n72025 , n72026 );
and ( n72028 , n70837 , n70838 );
and ( n72029 , n70839 , n70842 );
or ( n72030 , n72028 , n72029 );
xor ( n72031 , n72027 , n72030 );
nor ( n72032 , n31858 , n624 );
xor ( n72033 , n72031 , n72032 );
and ( n72034 , n70843 , n70844 );
and ( n72035 , n70845 , n70848 );
or ( n72036 , n72034 , n72035 );
xor ( n72037 , n72033 , n72036 );
nor ( n72038 , n33024 , n648 );
xor ( n72039 , n72037 , n72038 );
and ( n72040 , n70849 , n70850 );
and ( n72041 , n70851 , n70854 );
or ( n72042 , n72040 , n72041 );
xor ( n72043 , n72039 , n72042 );
nor ( n72044 , n34215 , n686 );
xor ( n72045 , n72043 , n72044 );
and ( n72046 , n70855 , n70856 );
and ( n72047 , n70857 , n70860 );
or ( n72048 , n72046 , n72047 );
xor ( n72049 , n72045 , n72048 );
nor ( n72050 , n35410 , n735 );
xor ( n72051 , n72049 , n72050 );
and ( n72052 , n70861 , n70862 );
and ( n72053 , n70863 , n70866 );
or ( n72054 , n72052 , n72053 );
xor ( n72055 , n72051 , n72054 );
nor ( n72056 , n36611 , n798 );
xor ( n72057 , n72055 , n72056 );
and ( n72058 , n70867 , n70868 );
and ( n72059 , n70869 , n70872 );
or ( n72060 , n72058 , n72059 );
xor ( n72061 , n72057 , n72060 );
nor ( n72062 , n37816 , n870 );
xor ( n72063 , n72061 , n72062 );
and ( n72064 , n70873 , n70874 );
and ( n72065 , n70875 , n70878 );
or ( n72066 , n72064 , n72065 );
xor ( n72067 , n72063 , n72066 );
nor ( n72068 , n39018 , n960 );
xor ( n72069 , n72067 , n72068 );
and ( n72070 , n70879 , n70880 );
and ( n72071 , n70881 , n70884 );
or ( n72072 , n72070 , n72071 );
xor ( n72073 , n72069 , n72072 );
nor ( n72074 , n40223 , n1064 );
xor ( n72075 , n72073 , n72074 );
and ( n72076 , n70885 , n70886 );
and ( n72077 , n70887 , n70890 );
or ( n72078 , n72076 , n72077 );
xor ( n72079 , n72075 , n72078 );
nor ( n72080 , n41428 , n1178 );
xor ( n72081 , n72079 , n72080 );
and ( n72082 , n70891 , n70892 );
and ( n72083 , n70893 , n70896 );
or ( n72084 , n72082 , n72083 );
xor ( n72085 , n72081 , n72084 );
nor ( n72086 , n42632 , n1305 );
xor ( n72087 , n72085 , n72086 );
and ( n72088 , n70897 , n70898 );
and ( n72089 , n70899 , n70902 );
or ( n72090 , n72088 , n72089 );
xor ( n72091 , n72087 , n72090 );
nor ( n72092 , n43834 , n1447 );
xor ( n72093 , n72091 , n72092 );
and ( n72094 , n70903 , n70904 );
and ( n72095 , n70905 , n70908 );
or ( n72096 , n72094 , n72095 );
xor ( n72097 , n72093 , n72096 );
nor ( n72098 , n45038 , n1600 );
xor ( n72099 , n72097 , n72098 );
and ( n72100 , n70909 , n70910 );
and ( n72101 , n70911 , n70914 );
or ( n72102 , n72100 , n72101 );
xor ( n72103 , n72099 , n72102 );
nor ( n72104 , n46239 , n1768 );
xor ( n72105 , n72103 , n72104 );
and ( n72106 , n70915 , n70916 );
and ( n72107 , n70917 , n70920 );
or ( n72108 , n72106 , n72107 );
xor ( n72109 , n72105 , n72108 );
nor ( n72110 , n47440 , n1947 );
xor ( n72111 , n72109 , n72110 );
and ( n72112 , n70921 , n70922 );
and ( n72113 , n70923 , n70926 );
or ( n72114 , n72112 , n72113 );
xor ( n72115 , n72111 , n72114 );
nor ( n72116 , n48641 , n2139 );
xor ( n72117 , n72115 , n72116 );
and ( n72118 , n70927 , n70928 );
and ( n72119 , n70929 , n70932 );
or ( n72120 , n72118 , n72119 );
xor ( n72121 , n72117 , n72120 );
nor ( n72122 , n49841 , n2345 );
xor ( n72123 , n72121 , n72122 );
and ( n72124 , n70933 , n70934 );
and ( n72125 , n70935 , n70938 );
or ( n72126 , n72124 , n72125 );
xor ( n72127 , n72123 , n72126 );
nor ( n72128 , n51040 , n2568 );
xor ( n72129 , n72127 , n72128 );
and ( n72130 , n70939 , n70940 );
and ( n72131 , n70941 , n70944 );
or ( n72132 , n72130 , n72131 );
xor ( n72133 , n72129 , n72132 );
nor ( n72134 , n52238 , n2799 );
xor ( n72135 , n72133 , n72134 );
and ( n72136 , n70945 , n70946 );
and ( n72137 , n70947 , n70950 );
or ( n72138 , n72136 , n72137 );
xor ( n72139 , n72135 , n72138 );
nor ( n72140 , n53432 , n3045 );
xor ( n72141 , n72139 , n72140 );
and ( n72142 , n70951 , n70952 );
and ( n72143 , n70953 , n70956 );
or ( n72144 , n72142 , n72143 );
xor ( n72145 , n72141 , n72144 );
nor ( n72146 , n54629 , n3302 );
xor ( n72147 , n72145 , n72146 );
and ( n72148 , n70957 , n70958 );
and ( n72149 , n70959 , n70962 );
or ( n72150 , n72148 , n72149 );
xor ( n72151 , n72147 , n72150 );
nor ( n72152 , n55826 , n3572 );
xor ( n72153 , n72151 , n72152 );
and ( n72154 , n70963 , n70964 );
and ( n72155 , n70965 , n70968 );
or ( n72156 , n72154 , n72155 );
xor ( n72157 , n72153 , n72156 );
nor ( n72158 , n57022 , n3855 );
xor ( n72159 , n72157 , n72158 );
and ( n72160 , n70969 , n70970 );
and ( n72161 , n70971 , n70974 );
or ( n72162 , n72160 , n72161 );
xor ( n72163 , n72159 , n72162 );
nor ( n72164 , n58217 , n4153 );
xor ( n72165 , n72163 , n72164 );
and ( n72166 , n70975 , n70976 );
and ( n72167 , n70977 , n70980 );
or ( n72168 , n72166 , n72167 );
xor ( n72169 , n72165 , n72168 );
nor ( n72170 , n59412 , n4460 );
xor ( n72171 , n72169 , n72170 );
and ( n72172 , n70981 , n70982 );
and ( n72173 , n70983 , n70986 );
or ( n72174 , n72172 , n72173 );
xor ( n72175 , n72171 , n72174 );
nor ( n72176 , n60600 , n4788 );
xor ( n72177 , n72175 , n72176 );
and ( n72178 , n70987 , n70988 );
and ( n72179 , n70989 , n70992 );
or ( n72180 , n72178 , n72179 );
xor ( n72181 , n72177 , n72180 );
nor ( n72182 , n61791 , n5128 );
xor ( n72183 , n72181 , n72182 );
and ( n72184 , n70993 , n70994 );
and ( n72185 , n70995 , n70998 );
or ( n72186 , n72184 , n72185 );
xor ( n72187 , n72183 , n72186 );
nor ( n72188 , n62982 , n5479 );
xor ( n72189 , n72187 , n72188 );
and ( n72190 , n70999 , n71000 );
and ( n72191 , n71001 , n71004 );
or ( n72192 , n72190 , n72191 );
xor ( n72193 , n72189 , n72192 );
nor ( n72194 , n64172 , n5840 );
xor ( n72195 , n72193 , n72194 );
and ( n72196 , n71005 , n71006 );
and ( n72197 , n71007 , n71010 );
or ( n72198 , n72196 , n72197 );
xor ( n72199 , n72195 , n72198 );
nor ( n72200 , n65360 , n6214 );
xor ( n72201 , n72199 , n72200 );
and ( n72202 , n71011 , n71012 );
and ( n72203 , n71013 , n71016 );
or ( n72204 , n72202 , n72203 );
xor ( n72205 , n72201 , n72204 );
nor ( n72206 , n66550 , n6598 );
xor ( n72207 , n72205 , n72206 );
and ( n72208 , n71017 , n71018 );
and ( n72209 , n71019 , n71022 );
or ( n72210 , n72208 , n72209 );
xor ( n72211 , n72207 , n72210 );
nor ( n72212 , n67736 , n6999 );
xor ( n72213 , n72211 , n72212 );
and ( n72214 , n71023 , n71024 );
and ( n72215 , n71025 , n71028 );
or ( n72216 , n72214 , n72215 );
xor ( n72217 , n72213 , n72216 );
nor ( n72218 , n68924 , n7415 );
xor ( n72219 , n72217 , n72218 );
and ( n72220 , n71029 , n71030 );
and ( n72221 , n71031 , n71034 );
or ( n72222 , n72220 , n72221 );
xor ( n72223 , n72219 , n72222 );
nor ( n72224 , n70110 , n7843 );
xor ( n72225 , n72223 , n72224 );
and ( n72226 , n71035 , n71036 );
and ( n72227 , n71037 , n71040 );
or ( n72228 , n72226 , n72227 );
xor ( n72229 , n72225 , n72228 );
nor ( n72230 , n71292 , n8283 );
xor ( n72231 , n72229 , n72230 );
and ( n72232 , n71041 , n71042 );
and ( n72233 , n71043 , n71046 );
or ( n72234 , n72232 , n72233 );
xor ( n72235 , n72231 , n72234 );
and ( n72236 , n71059 , n71063 );
and ( n72237 , n71063 , n71278 );
and ( n72238 , n71059 , n71278 );
or ( n72239 , n72236 , n72237 , n72238 );
and ( n72240 , n33774 , n6971 );
not ( n72241 , n6971 );
nor ( n72242 , n72240 , n72241 );
xor ( n72243 , n72239 , n72242 );
and ( n72244 , n71069 , n71070 );
and ( n72245 , n71070 , n71138 );
and ( n72246 , n71069 , n71138 );
or ( n72247 , n72244 , n72245 , n72246 );
and ( n72248 , n71065 , n71139 );
and ( n72249 , n71139 , n71277 );
and ( n72250 , n71065 , n71277 );
or ( n72251 , n72248 , n72249 , n72250 );
xor ( n72252 , n72247 , n72251 );
and ( n72253 , n71161 , n71276 );
and ( n72254 , n71075 , n71079 );
and ( n72255 , n71079 , n71137 );
and ( n72256 , n71075 , n71137 );
or ( n72257 , n72254 , n72255 , n72256 );
and ( n72258 , n71165 , n71275 );
xor ( n72259 , n72257 , n72258 );
and ( n72260 , n71106 , n71110 );
and ( n72261 , n71110 , n71116 );
and ( n72262 , n71106 , n71116 );
or ( n72263 , n72260 , n72261 , n72262 );
and ( n72264 , n71084 , n71088 );
and ( n72265 , n71088 , n71136 );
and ( n72266 , n71084 , n71136 );
or ( n72267 , n72264 , n72265 , n72266 );
xor ( n72268 , n72263 , n72267 );
and ( n72269 , n71093 , n71097 );
and ( n72270 , n71097 , n71135 );
and ( n72271 , n71093 , n71135 );
or ( n72272 , n72269 , n72270 , n72271 );
and ( n72273 , n71173 , n71198 );
and ( n72274 , n71198 , n71236 );
and ( n72275 , n71173 , n71236 );
or ( n72276 , n72273 , n72274 , n72275 );
xor ( n72277 , n72272 , n72276 );
and ( n72278 , n71102 , n71117 );
and ( n72279 , n71117 , n71134 );
and ( n72280 , n71102 , n71134 );
or ( n72281 , n72278 , n72279 , n72280 );
and ( n72282 , n71177 , n71181 );
and ( n72283 , n71181 , n71197 );
and ( n72284 , n71177 , n71197 );
or ( n72285 , n72282 , n72283 , n72284 );
xor ( n72286 , n72281 , n72285 );
and ( n72287 , n71122 , n71127 );
and ( n72288 , n71127 , n71133 );
and ( n72289 , n71122 , n71133 );
or ( n72290 , n72287 , n72288 , n72289 );
and ( n72291 , n71112 , n71113 );
and ( n72292 , n71113 , n71115 );
and ( n72293 , n71112 , n71115 );
or ( n72294 , n72291 , n72292 , n72293 );
and ( n72295 , n71123 , n71124 );
and ( n72296 , n71124 , n71126 );
and ( n72297 , n71123 , n71126 );
or ( n72298 , n72295 , n72296 , n72297 );
xor ( n72299 , n72294 , n72298 );
and ( n72300 , n30695 , n8243 );
and ( n72301 , n31836 , n7662 );
xor ( n72302 , n72300 , n72301 );
and ( n72303 , n32649 , n7310 );
xor ( n72304 , n72302 , n72303 );
xor ( n72305 , n72299 , n72304 );
xor ( n72306 , n72290 , n72305 );
and ( n72307 , n71129 , n71130 );
and ( n72308 , n71130 , n71132 );
and ( n72309 , n71129 , n71132 );
or ( n72310 , n72307 , n72308 , n72309 );
and ( n72311 , n27361 , n10239 );
and ( n72312 , n28456 , n9348 );
xor ( n72313 , n72311 , n72312 );
and ( n72314 , n29559 , n8669 );
xor ( n72315 , n72313 , n72314 );
xor ( n72316 , n72310 , n72315 );
and ( n72317 , n24214 , n12531 );
and ( n72318 , n25243 , n11718 );
xor ( n72319 , n72317 , n72318 );
and ( n72320 , n26296 , n10977 );
xor ( n72321 , n72319 , n72320 );
xor ( n72322 , n72316 , n72321 );
xor ( n72323 , n72306 , n72322 );
xor ( n72324 , n72286 , n72323 );
xor ( n72325 , n72277 , n72324 );
xor ( n72326 , n72268 , n72325 );
xor ( n72327 , n72259 , n72326 );
xor ( n72328 , n72253 , n72327 );
not ( n72329 , n6816 );
and ( n72330 , n34193 , n6816 );
nor ( n72331 , n72329 , n72330 );
and ( n72332 , n71150 , n71151 );
and ( n72333 , n71151 , n71153 );
and ( n72334 , n71150 , n71153 );
or ( n72335 , n72332 , n72333 , n72334 );
and ( n72336 , n71158 , n71159 );
xor ( n72337 , n72335 , n72336 );
and ( n72338 , n7385 , n32999 );
and ( n72339 , n7808 , n31761 );
xor ( n72340 , n72338 , n72339 );
and ( n72341 , n8079 , n30629 );
xor ( n72342 , n72340 , n72341 );
xor ( n72343 , n72337 , n72342 );
xor ( n72344 , n72331 , n72343 );
and ( n72345 , n71169 , n71237 );
and ( n72346 , n71237 , n71274 );
and ( n72347 , n71169 , n71274 );
or ( n72348 , n72345 , n72346 , n72347 );
and ( n72349 , n71242 , n71246 );
and ( n72350 , n71246 , n71273 );
and ( n72351 , n71242 , n71273 );
or ( n72352 , n72349 , n72350 , n72351 );
and ( n72353 , n71203 , n71219 );
and ( n72354 , n71219 , n71235 );
and ( n72355 , n71203 , n71235 );
or ( n72356 , n72353 , n72354 , n72355 );
and ( n72357 , n71186 , n71190 );
and ( n72358 , n71190 , n71196 );
and ( n72359 , n71186 , n71196 );
or ( n72360 , n72357 , n72358 , n72359 );
and ( n72361 , n71207 , n71212 );
and ( n72362 , n71212 , n71218 );
and ( n72363 , n71207 , n71218 );
or ( n72364 , n72361 , n72362 , n72363 );
xor ( n72365 , n72360 , n72364 );
and ( n72366 , n71192 , n71193 );
and ( n72367 , n71193 , n71195 );
and ( n72368 , n71192 , n71195 );
or ( n72369 , n72366 , n72367 , n72368 );
and ( n72370 , n71208 , n71209 );
and ( n72371 , n71209 , n71211 );
and ( n72372 , n71208 , n71211 );
or ( n72373 , n72370 , n72371 , n72372 );
xor ( n72374 , n72369 , n72373 );
and ( n72375 , n21216 , n14838 );
and ( n72376 , n22186 , n14044 );
xor ( n72377 , n72375 , n72376 );
and ( n72378 , n22892 , n13256 );
xor ( n72379 , n72377 , n72378 );
xor ( n72380 , n72374 , n72379 );
xor ( n72381 , n72365 , n72380 );
xor ( n72382 , n72356 , n72381 );
and ( n72383 , n71224 , n71228 );
and ( n72384 , n71228 , n71234 );
and ( n72385 , n71224 , n71234 );
or ( n72386 , n72383 , n72384 , n72385 );
and ( n72387 , n71214 , n71215 );
and ( n72388 , n71215 , n71217 );
and ( n72389 , n71214 , n71217 );
or ( n72390 , n72387 , n72388 , n72389 );
and ( n72391 , n18144 , n17422 );
and ( n72392 , n19324 , n16550 );
xor ( n72393 , n72391 , n72392 );
and ( n72394 , n20233 , n15691 );
xor ( n72395 , n72393 , n72394 );
xor ( n72396 , n72390 , n72395 );
and ( n72397 , n15758 , n20156 );
and ( n72398 , n16637 , n19222 );
xor ( n72399 , n72397 , n72398 );
and ( n72400 , n17512 , n18407 );
xor ( n72401 , n72399 , n72400 );
xor ( n72402 , n72396 , n72401 );
xor ( n72403 , n72386 , n72402 );
and ( n72404 , n71230 , n71231 );
and ( n72405 , n71231 , n71233 );
and ( n72406 , n71230 , n71233 );
or ( n72407 , n72404 , n72405 , n72406 );
and ( n72408 , n71261 , n71262 );
and ( n72409 , n71262 , n71264 );
and ( n72410 , n71261 , n71264 );
or ( n72411 , n72408 , n72409 , n72410 );
xor ( n72412 , n72407 , n72411 );
and ( n72413 , n13322 , n23075 );
and ( n72414 , n14118 , n22065 );
xor ( n72415 , n72413 , n72414 );
and ( n72416 , n14938 , n20976 );
xor ( n72417 , n72415 , n72416 );
xor ( n72418 , n72412 , n72417 );
xor ( n72419 , n72403 , n72418 );
xor ( n72420 , n72382 , n72419 );
xor ( n72421 , n72352 , n72420 );
and ( n72422 , n71251 , n71255 );
and ( n72423 , n71255 , n71272 );
and ( n72424 , n71251 , n71272 );
or ( n72425 , n72422 , n72423 , n72424 );
and ( n72426 , n71155 , n71160 );
xor ( n72427 , n72425 , n72426 );
and ( n72428 , n71144 , n71148 );
and ( n72429 , n71148 , n71154 );
and ( n72430 , n71144 , n71154 );
or ( n72431 , n72428 , n72429 , n72430 );
and ( n72432 , n71260 , n71265 );
and ( n72433 , n71265 , n71271 );
and ( n72434 , n71260 , n71271 );
or ( n72435 , n72432 , n72433 , n72434 );
xor ( n72436 , n72431 , n72435 );
and ( n72437 , n71267 , n71268 );
and ( n72438 , n71268 , n71270 );
and ( n72439 , n71267 , n71270 );
or ( n72440 , n72437 , n72438 , n72439 );
and ( n72441 , n11015 , n26216 );
and ( n72442 , n11769 , n25163 );
xor ( n72443 , n72441 , n72442 );
and ( n72444 , n12320 , n24137 );
xor ( n72445 , n72443 , n72444 );
xor ( n72446 , n72440 , n72445 );
and ( n72447 , n8718 , n29508 );
and ( n72448 , n9400 , n28406 );
xor ( n72449 , n72447 , n72448 );
and ( n72450 , n10291 , n27296 );
xor ( n72451 , n72449 , n72450 );
xor ( n72452 , n72446 , n72451 );
xor ( n72453 , n72436 , n72452 );
xor ( n72454 , n72427 , n72453 );
xor ( n72455 , n72421 , n72454 );
xor ( n72456 , n72348 , n72455 );
xor ( n72457 , n72344 , n72456 );
xor ( n72458 , n72328 , n72457 );
xor ( n72459 , n72252 , n72458 );
xor ( n72460 , n72243 , n72459 );
and ( n72461 , n71051 , n71054 );
and ( n72462 , n71054 , n71279 );
and ( n72463 , n71051 , n71279 );
or ( n72464 , n72461 , n72462 , n72463 );
xor ( n72465 , n72460 , n72464 );
and ( n72466 , n71280 , n71284 );
and ( n72467 , n71285 , n71288 );
or ( n72468 , n72466 , n72467 );
xor ( n72469 , n72465 , n72468 );
buf ( n72470 , n72469 );
buf ( n72471 , n72470 );
not ( n72472 , n72471 );
nor ( n72473 , n72472 , n8739 );
xor ( n72474 , n72235 , n72473 );
and ( n72475 , n71047 , n71293 );
and ( n72476 , n71294 , n71297 );
or ( n72477 , n72475 , n72476 );
xor ( n72478 , n72474 , n72477 );
buf ( n72479 , n72478 );
buf ( n72480 , n72479 );
not ( n72481 , n72480 );
buf ( n72482 , n594 );
not ( n72483 , n72482 );
nor ( n72484 , n72481 , n72483 );
xor ( n72485 , n71861 , n72484 );
xor ( n72486 , n71309 , n71858 );
nor ( n72487 , n71301 , n72483 );
and ( n72488 , n72486 , n72487 );
xor ( n72489 , n72486 , n72487 );
xor ( n72490 , n71313 , n71856 );
nor ( n72491 , n70119 , n72483 );
and ( n72492 , n72490 , n72491 );
xor ( n72493 , n72490 , n72491 );
xor ( n72494 , n71317 , n71854 );
nor ( n72495 , n68933 , n72483 );
and ( n72496 , n72494 , n72495 );
xor ( n72497 , n72494 , n72495 );
xor ( n72498 , n71321 , n71852 );
nor ( n72499 , n67745 , n72483 );
and ( n72500 , n72498 , n72499 );
xor ( n72501 , n72498 , n72499 );
xor ( n72502 , n71325 , n71850 );
nor ( n72503 , n66559 , n72483 );
and ( n72504 , n72502 , n72503 );
xor ( n72505 , n72502 , n72503 );
xor ( n72506 , n71329 , n71848 );
nor ( n72507 , n65369 , n72483 );
and ( n72508 , n72506 , n72507 );
xor ( n72509 , n72506 , n72507 );
xor ( n72510 , n71333 , n71846 );
nor ( n72511 , n64181 , n72483 );
and ( n72512 , n72510 , n72511 );
xor ( n72513 , n72510 , n72511 );
xor ( n72514 , n71337 , n71844 );
nor ( n72515 , n62991 , n72483 );
and ( n72516 , n72514 , n72515 );
xor ( n72517 , n72514 , n72515 );
xor ( n72518 , n71341 , n71842 );
nor ( n72519 , n61800 , n72483 );
and ( n72520 , n72518 , n72519 );
xor ( n72521 , n72518 , n72519 );
xor ( n72522 , n71345 , n71840 );
nor ( n72523 , n60609 , n72483 );
and ( n72524 , n72522 , n72523 );
xor ( n72525 , n72522 , n72523 );
xor ( n72526 , n71349 , n71838 );
nor ( n72527 , n59421 , n72483 );
and ( n72528 , n72526 , n72527 );
xor ( n72529 , n72526 , n72527 );
xor ( n72530 , n71353 , n71836 );
nor ( n72531 , n58226 , n72483 );
and ( n72532 , n72530 , n72531 );
xor ( n72533 , n72530 , n72531 );
xor ( n72534 , n71357 , n71834 );
nor ( n72535 , n57031 , n72483 );
and ( n72536 , n72534 , n72535 );
xor ( n72537 , n72534 , n72535 );
xor ( n72538 , n71361 , n71832 );
nor ( n72539 , n55835 , n72483 );
and ( n72540 , n72538 , n72539 );
xor ( n72541 , n72538 , n72539 );
xor ( n72542 , n71365 , n71830 );
nor ( n72543 , n54638 , n72483 );
and ( n72544 , n72542 , n72543 );
xor ( n72545 , n72542 , n72543 );
xor ( n72546 , n71369 , n71828 );
nor ( n72547 , n53441 , n72483 );
and ( n72548 , n72546 , n72547 );
xor ( n72549 , n72546 , n72547 );
xor ( n72550 , n71373 , n71826 );
nor ( n72551 , n52247 , n72483 );
and ( n72552 , n72550 , n72551 );
xor ( n72553 , n72550 , n72551 );
xor ( n72554 , n71377 , n71824 );
nor ( n72555 , n51049 , n72483 );
and ( n72556 , n72554 , n72555 );
xor ( n72557 , n72554 , n72555 );
xor ( n72558 , n71381 , n71822 );
nor ( n72559 , n49850 , n72483 );
and ( n72560 , n72558 , n72559 );
xor ( n72561 , n72558 , n72559 );
xor ( n72562 , n71385 , n71820 );
nor ( n72563 , n48650 , n72483 );
and ( n72564 , n72562 , n72563 );
xor ( n72565 , n72562 , n72563 );
xor ( n72566 , n71389 , n71818 );
nor ( n72567 , n47449 , n72483 );
and ( n72568 , n72566 , n72567 );
xor ( n72569 , n72566 , n72567 );
xor ( n72570 , n71393 , n71816 );
nor ( n72571 , n46248 , n72483 );
and ( n72572 , n72570 , n72571 );
xor ( n72573 , n72570 , n72571 );
xor ( n72574 , n71397 , n71814 );
nor ( n72575 , n45047 , n72483 );
and ( n72576 , n72574 , n72575 );
xor ( n72577 , n72574 , n72575 );
xor ( n72578 , n71401 , n71812 );
nor ( n72579 , n43843 , n72483 );
and ( n72580 , n72578 , n72579 );
xor ( n72581 , n72578 , n72579 );
xor ( n72582 , n71405 , n71810 );
nor ( n72583 , n42641 , n72483 );
and ( n72584 , n72582 , n72583 );
xor ( n72585 , n72582 , n72583 );
xor ( n72586 , n71409 , n71808 );
nor ( n72587 , n41437 , n72483 );
and ( n72588 , n72586 , n72587 );
xor ( n72589 , n72586 , n72587 );
xor ( n72590 , n71413 , n71806 );
nor ( n72591 , n40232 , n72483 );
and ( n72592 , n72590 , n72591 );
xor ( n72593 , n72590 , n72591 );
xor ( n72594 , n71417 , n71804 );
nor ( n72595 , n39027 , n72483 );
and ( n72596 , n72594 , n72595 );
xor ( n72597 , n72594 , n72595 );
xor ( n72598 , n71421 , n71802 );
nor ( n72599 , n37825 , n72483 );
and ( n72600 , n72598 , n72599 );
xor ( n72601 , n72598 , n72599 );
xor ( n72602 , n71425 , n71800 );
nor ( n72603 , n36620 , n72483 );
and ( n72604 , n72602 , n72603 );
xor ( n72605 , n72602 , n72603 );
xor ( n72606 , n71429 , n71798 );
nor ( n72607 , n35419 , n72483 );
and ( n72608 , n72606 , n72607 );
xor ( n72609 , n72606 , n72607 );
xor ( n72610 , n71433 , n71796 );
nor ( n72611 , n34224 , n72483 );
and ( n72612 , n72610 , n72611 );
xor ( n72613 , n72610 , n72611 );
xor ( n72614 , n71437 , n71794 );
nor ( n72615 , n33033 , n72483 );
and ( n72616 , n72614 , n72615 );
xor ( n72617 , n72614 , n72615 );
xor ( n72618 , n71441 , n71792 );
nor ( n72619 , n31867 , n72483 );
and ( n72620 , n72618 , n72619 );
xor ( n72621 , n72618 , n72619 );
xor ( n72622 , n71445 , n71790 );
nor ( n72623 , n30725 , n72483 );
and ( n72624 , n72622 , n72623 );
xor ( n72625 , n72622 , n72623 );
xor ( n72626 , n71449 , n71788 );
nor ( n72627 , n29596 , n72483 );
and ( n72628 , n72626 , n72627 );
xor ( n72629 , n72626 , n72627 );
xor ( n72630 , n71453 , n71786 );
nor ( n72631 , n28487 , n72483 );
and ( n72632 , n72630 , n72631 );
xor ( n72633 , n72630 , n72631 );
xor ( n72634 , n71457 , n71784 );
nor ( n72635 , n27397 , n72483 );
and ( n72636 , n72634 , n72635 );
xor ( n72637 , n72634 , n72635 );
xor ( n72638 , n71461 , n71782 );
nor ( n72639 , n26326 , n72483 );
and ( n72640 , n72638 , n72639 );
xor ( n72641 , n72638 , n72639 );
xor ( n72642 , n71465 , n71780 );
nor ( n72643 , n25272 , n72483 );
and ( n72644 , n72642 , n72643 );
xor ( n72645 , n72642 , n72643 );
xor ( n72646 , n71469 , n71778 );
nor ( n72647 , n24242 , n72483 );
and ( n72648 , n72646 , n72647 );
xor ( n72649 , n72646 , n72647 );
xor ( n72650 , n71473 , n71776 );
nor ( n72651 , n23225 , n72483 );
and ( n72652 , n72650 , n72651 );
xor ( n72653 , n72650 , n72651 );
xor ( n72654 , n71477 , n71774 );
nor ( n72655 , n22231 , n72483 );
and ( n72656 , n72654 , n72655 );
xor ( n72657 , n72654 , n72655 );
xor ( n72658 , n71481 , n71772 );
nor ( n72659 , n21258 , n72483 );
and ( n72660 , n72658 , n72659 );
xor ( n72661 , n72658 , n72659 );
xor ( n72662 , n71485 , n71770 );
nor ( n72663 , n20303 , n72483 );
and ( n72664 , n72662 , n72663 );
xor ( n72665 , n72662 , n72663 );
xor ( n72666 , n71489 , n71768 );
nor ( n72667 , n19365 , n72483 );
and ( n72668 , n72666 , n72667 );
xor ( n72669 , n72666 , n72667 );
xor ( n72670 , n71493 , n71766 );
nor ( n72671 , n18448 , n72483 );
and ( n72672 , n72670 , n72671 );
xor ( n72673 , n72670 , n72671 );
xor ( n72674 , n71497 , n71764 );
nor ( n72675 , n17548 , n72483 );
and ( n72676 , n72674 , n72675 );
xor ( n72677 , n72674 , n72675 );
xor ( n72678 , n71501 , n71762 );
nor ( n72679 , n16669 , n72483 );
and ( n72680 , n72678 , n72679 );
xor ( n72681 , n72678 , n72679 );
xor ( n72682 , n71505 , n71760 );
nor ( n72683 , n15809 , n72483 );
and ( n72684 , n72682 , n72683 );
xor ( n72685 , n72682 , n72683 );
xor ( n72686 , n71509 , n71758 );
nor ( n72687 , n14968 , n72483 );
and ( n72688 , n72686 , n72687 );
xor ( n72689 , n72686 , n72687 );
xor ( n72690 , n71513 , n71756 );
nor ( n72691 , n14147 , n72483 );
and ( n72692 , n72690 , n72691 );
xor ( n72693 , n72690 , n72691 );
xor ( n72694 , n71517 , n71754 );
nor ( n72695 , n13349 , n72483 );
and ( n72696 , n72694 , n72695 );
xor ( n72697 , n72694 , n72695 );
xor ( n72698 , n71521 , n71752 );
nor ( n72699 , n12564 , n72483 );
and ( n72700 , n72698 , n72699 );
xor ( n72701 , n72698 , n72699 );
xor ( n72702 , n71525 , n71750 );
nor ( n72703 , n11799 , n72483 );
and ( n72704 , n72702 , n72703 );
xor ( n72705 , n72702 , n72703 );
xor ( n72706 , n71529 , n71748 );
nor ( n72707 , n11050 , n72483 );
and ( n72708 , n72706 , n72707 );
xor ( n72709 , n72706 , n72707 );
xor ( n72710 , n71533 , n71746 );
nor ( n72711 , n10321 , n72483 );
and ( n72712 , n72710 , n72711 );
xor ( n72713 , n72710 , n72711 );
xor ( n72714 , n71537 , n71744 );
nor ( n72715 , n9429 , n72483 );
and ( n72716 , n72714 , n72715 );
xor ( n72717 , n72714 , n72715 );
xor ( n72718 , n71541 , n71742 );
nor ( n72719 , n8949 , n72483 );
and ( n72720 , n72718 , n72719 );
xor ( n72721 , n72718 , n72719 );
xor ( n72722 , n71545 , n71740 );
nor ( n72723 , n9437 , n72483 );
and ( n72724 , n72722 , n72723 );
xor ( n72725 , n72722 , n72723 );
xor ( n72726 , n71549 , n71738 );
nor ( n72727 , n9446 , n72483 );
and ( n72728 , n72726 , n72727 );
xor ( n72729 , n72726 , n72727 );
xor ( n72730 , n71553 , n71736 );
nor ( n72731 , n9455 , n72483 );
and ( n72732 , n72730 , n72731 );
xor ( n72733 , n72730 , n72731 );
xor ( n72734 , n71557 , n71734 );
nor ( n72735 , n9464 , n72483 );
and ( n72736 , n72734 , n72735 );
xor ( n72737 , n72734 , n72735 );
xor ( n72738 , n71561 , n71732 );
nor ( n72739 , n9473 , n72483 );
and ( n72740 , n72738 , n72739 );
xor ( n72741 , n72738 , n72739 );
xor ( n72742 , n71565 , n71730 );
nor ( n72743 , n9482 , n72483 );
and ( n72744 , n72742 , n72743 );
xor ( n72745 , n72742 , n72743 );
xor ( n72746 , n71569 , n71728 );
nor ( n72747 , n9491 , n72483 );
and ( n72748 , n72746 , n72747 );
xor ( n72749 , n72746 , n72747 );
xor ( n72750 , n71573 , n71726 );
nor ( n72751 , n9500 , n72483 );
and ( n72752 , n72750 , n72751 );
xor ( n72753 , n72750 , n72751 );
xor ( n72754 , n71577 , n71724 );
nor ( n72755 , n9509 , n72483 );
and ( n72756 , n72754 , n72755 );
xor ( n72757 , n72754 , n72755 );
xor ( n72758 , n71581 , n71722 );
nor ( n72759 , n9518 , n72483 );
and ( n72760 , n72758 , n72759 );
xor ( n72761 , n72758 , n72759 );
xor ( n72762 , n71585 , n71720 );
nor ( n72763 , n9527 , n72483 );
and ( n72764 , n72762 , n72763 );
xor ( n72765 , n72762 , n72763 );
xor ( n72766 , n71589 , n71718 );
nor ( n72767 , n9536 , n72483 );
and ( n72768 , n72766 , n72767 );
xor ( n72769 , n72766 , n72767 );
xor ( n72770 , n71593 , n71716 );
nor ( n72771 , n9545 , n72483 );
and ( n72772 , n72770 , n72771 );
xor ( n72773 , n72770 , n72771 );
xor ( n72774 , n71597 , n71714 );
nor ( n72775 , n9554 , n72483 );
and ( n72776 , n72774 , n72775 );
xor ( n72777 , n72774 , n72775 );
xor ( n72778 , n71601 , n71712 );
nor ( n72779 , n9563 , n72483 );
and ( n72780 , n72778 , n72779 );
xor ( n72781 , n72778 , n72779 );
xor ( n72782 , n71605 , n71710 );
nor ( n72783 , n9572 , n72483 );
and ( n72784 , n72782 , n72783 );
xor ( n72785 , n72782 , n72783 );
xor ( n72786 , n71609 , n71708 );
nor ( n72787 , n9581 , n72483 );
and ( n72788 , n72786 , n72787 );
xor ( n72789 , n72786 , n72787 );
xor ( n72790 , n71613 , n71706 );
nor ( n72791 , n9590 , n72483 );
and ( n72792 , n72790 , n72791 );
xor ( n72793 , n72790 , n72791 );
xor ( n72794 , n71617 , n71704 );
nor ( n72795 , n9599 , n72483 );
and ( n72796 , n72794 , n72795 );
xor ( n72797 , n72794 , n72795 );
xor ( n72798 , n71621 , n71702 );
nor ( n72799 , n9608 , n72483 );
and ( n72800 , n72798 , n72799 );
xor ( n72801 , n72798 , n72799 );
xor ( n72802 , n71625 , n71700 );
nor ( n72803 , n9617 , n72483 );
and ( n72804 , n72802 , n72803 );
xor ( n72805 , n72802 , n72803 );
xor ( n72806 , n71629 , n71698 );
nor ( n72807 , n9626 , n72483 );
and ( n72808 , n72806 , n72807 );
xor ( n72809 , n72806 , n72807 );
xor ( n72810 , n71633 , n71696 );
nor ( n72811 , n9635 , n72483 );
and ( n72812 , n72810 , n72811 );
xor ( n72813 , n72810 , n72811 );
xor ( n72814 , n71637 , n71694 );
nor ( n72815 , n9644 , n72483 );
and ( n72816 , n72814 , n72815 );
xor ( n72817 , n72814 , n72815 );
xor ( n72818 , n71641 , n71692 );
nor ( n72819 , n9653 , n72483 );
and ( n72820 , n72818 , n72819 );
xor ( n72821 , n72818 , n72819 );
xor ( n72822 , n71645 , n71690 );
nor ( n72823 , n9662 , n72483 );
and ( n72824 , n72822 , n72823 );
xor ( n72825 , n72822 , n72823 );
xor ( n72826 , n71649 , n71688 );
nor ( n72827 , n9671 , n72483 );
and ( n72828 , n72826 , n72827 );
xor ( n72829 , n72826 , n72827 );
xor ( n72830 , n71653 , n71686 );
nor ( n72831 , n9680 , n72483 );
and ( n72832 , n72830 , n72831 );
xor ( n72833 , n72830 , n72831 );
xor ( n72834 , n71657 , n71684 );
nor ( n72835 , n9689 , n72483 );
and ( n72836 , n72834 , n72835 );
xor ( n72837 , n72834 , n72835 );
xor ( n72838 , n71661 , n71682 );
nor ( n72839 , n9698 , n72483 );
and ( n72840 , n72838 , n72839 );
xor ( n72841 , n72838 , n72839 );
xor ( n72842 , n71665 , n71680 );
nor ( n72843 , n9707 , n72483 );
and ( n72844 , n72842 , n72843 );
xor ( n72845 , n72842 , n72843 );
xor ( n72846 , n71669 , n71678 );
nor ( n72847 , n9716 , n72483 );
and ( n72848 , n72846 , n72847 );
xor ( n72849 , n72846 , n72847 );
xor ( n72850 , n71673 , n71676 );
nor ( n72851 , n9725 , n72483 );
and ( n72852 , n72850 , n72851 );
xor ( n72853 , n72850 , n72851 );
xor ( n72854 , n71674 , n71675 );
nor ( n72855 , n9734 , n72483 );
and ( n72856 , n72854 , n72855 );
xor ( n72857 , n72854 , n72855 );
nor ( n72858 , n9752 , n71303 );
nor ( n72859 , n9743 , n72483 );
and ( n72860 , n72858 , n72859 );
and ( n72861 , n72857 , n72860 );
or ( n72862 , n72856 , n72861 );
and ( n72863 , n72853 , n72862 );
or ( n72864 , n72852 , n72863 );
and ( n72865 , n72849 , n72864 );
or ( n72866 , n72848 , n72865 );
and ( n72867 , n72845 , n72866 );
or ( n72868 , n72844 , n72867 );
and ( n72869 , n72841 , n72868 );
or ( n72870 , n72840 , n72869 );
and ( n72871 , n72837 , n72870 );
or ( n72872 , n72836 , n72871 );
and ( n72873 , n72833 , n72872 );
or ( n72874 , n72832 , n72873 );
and ( n72875 , n72829 , n72874 );
or ( n72876 , n72828 , n72875 );
and ( n72877 , n72825 , n72876 );
or ( n72878 , n72824 , n72877 );
and ( n72879 , n72821 , n72878 );
or ( n72880 , n72820 , n72879 );
and ( n72881 , n72817 , n72880 );
or ( n72882 , n72816 , n72881 );
and ( n72883 , n72813 , n72882 );
or ( n72884 , n72812 , n72883 );
and ( n72885 , n72809 , n72884 );
or ( n72886 , n72808 , n72885 );
and ( n72887 , n72805 , n72886 );
or ( n72888 , n72804 , n72887 );
and ( n72889 , n72801 , n72888 );
or ( n72890 , n72800 , n72889 );
and ( n72891 , n72797 , n72890 );
or ( n72892 , n72796 , n72891 );
and ( n72893 , n72793 , n72892 );
or ( n72894 , n72792 , n72893 );
and ( n72895 , n72789 , n72894 );
or ( n72896 , n72788 , n72895 );
and ( n72897 , n72785 , n72896 );
or ( n72898 , n72784 , n72897 );
and ( n72899 , n72781 , n72898 );
or ( n72900 , n72780 , n72899 );
and ( n72901 , n72777 , n72900 );
or ( n72902 , n72776 , n72901 );
and ( n72903 , n72773 , n72902 );
or ( n72904 , n72772 , n72903 );
and ( n72905 , n72769 , n72904 );
or ( n72906 , n72768 , n72905 );
and ( n72907 , n72765 , n72906 );
or ( n72908 , n72764 , n72907 );
and ( n72909 , n72761 , n72908 );
or ( n72910 , n72760 , n72909 );
and ( n72911 , n72757 , n72910 );
or ( n72912 , n72756 , n72911 );
and ( n72913 , n72753 , n72912 );
or ( n72914 , n72752 , n72913 );
and ( n72915 , n72749 , n72914 );
or ( n72916 , n72748 , n72915 );
and ( n72917 , n72745 , n72916 );
or ( n72918 , n72744 , n72917 );
and ( n72919 , n72741 , n72918 );
or ( n72920 , n72740 , n72919 );
and ( n72921 , n72737 , n72920 );
or ( n72922 , n72736 , n72921 );
and ( n72923 , n72733 , n72922 );
or ( n72924 , n72732 , n72923 );
and ( n72925 , n72729 , n72924 );
or ( n72926 , n72728 , n72925 );
and ( n72927 , n72725 , n72926 );
or ( n72928 , n72724 , n72927 );
and ( n72929 , n72721 , n72928 );
or ( n72930 , n72720 , n72929 );
and ( n72931 , n72717 , n72930 );
or ( n72932 , n72716 , n72931 );
and ( n72933 , n72713 , n72932 );
or ( n72934 , n72712 , n72933 );
and ( n72935 , n72709 , n72934 );
or ( n72936 , n72708 , n72935 );
and ( n72937 , n72705 , n72936 );
or ( n72938 , n72704 , n72937 );
and ( n72939 , n72701 , n72938 );
or ( n72940 , n72700 , n72939 );
and ( n72941 , n72697 , n72940 );
or ( n72942 , n72696 , n72941 );
and ( n72943 , n72693 , n72942 );
or ( n72944 , n72692 , n72943 );
and ( n72945 , n72689 , n72944 );
or ( n72946 , n72688 , n72945 );
and ( n72947 , n72685 , n72946 );
or ( n72948 , n72684 , n72947 );
and ( n72949 , n72681 , n72948 );
or ( n72950 , n72680 , n72949 );
and ( n72951 , n72677 , n72950 );
or ( n72952 , n72676 , n72951 );
and ( n72953 , n72673 , n72952 );
or ( n72954 , n72672 , n72953 );
and ( n72955 , n72669 , n72954 );
or ( n72956 , n72668 , n72955 );
and ( n72957 , n72665 , n72956 );
or ( n72958 , n72664 , n72957 );
and ( n72959 , n72661 , n72958 );
or ( n72960 , n72660 , n72959 );
and ( n72961 , n72657 , n72960 );
or ( n72962 , n72656 , n72961 );
and ( n72963 , n72653 , n72962 );
or ( n72964 , n72652 , n72963 );
and ( n72965 , n72649 , n72964 );
or ( n72966 , n72648 , n72965 );
and ( n72967 , n72645 , n72966 );
or ( n72968 , n72644 , n72967 );
and ( n72969 , n72641 , n72968 );
or ( n72970 , n72640 , n72969 );
and ( n72971 , n72637 , n72970 );
or ( n72972 , n72636 , n72971 );
and ( n72973 , n72633 , n72972 );
or ( n72974 , n72632 , n72973 );
and ( n72975 , n72629 , n72974 );
or ( n72976 , n72628 , n72975 );
and ( n72977 , n72625 , n72976 );
or ( n72978 , n72624 , n72977 );
and ( n72979 , n72621 , n72978 );
or ( n72980 , n72620 , n72979 );
and ( n72981 , n72617 , n72980 );
or ( n72982 , n72616 , n72981 );
and ( n72983 , n72613 , n72982 );
or ( n72984 , n72612 , n72983 );
and ( n72985 , n72609 , n72984 );
or ( n72986 , n72608 , n72985 );
and ( n72987 , n72605 , n72986 );
or ( n72988 , n72604 , n72987 );
and ( n72989 , n72601 , n72988 );
or ( n72990 , n72600 , n72989 );
and ( n72991 , n72597 , n72990 );
or ( n72992 , n72596 , n72991 );
and ( n72993 , n72593 , n72992 );
or ( n72994 , n72592 , n72993 );
and ( n72995 , n72589 , n72994 );
or ( n72996 , n72588 , n72995 );
and ( n72997 , n72585 , n72996 );
or ( n72998 , n72584 , n72997 );
and ( n72999 , n72581 , n72998 );
or ( n73000 , n72580 , n72999 );
and ( n73001 , n72577 , n73000 );
or ( n73002 , n72576 , n73001 );
and ( n73003 , n72573 , n73002 );
or ( n73004 , n72572 , n73003 );
and ( n73005 , n72569 , n73004 );
or ( n73006 , n72568 , n73005 );
and ( n73007 , n72565 , n73006 );
or ( n73008 , n72564 , n73007 );
and ( n73009 , n72561 , n73008 );
or ( n73010 , n72560 , n73009 );
and ( n73011 , n72557 , n73010 );
or ( n73012 , n72556 , n73011 );
and ( n73013 , n72553 , n73012 );
or ( n73014 , n72552 , n73013 );
and ( n73015 , n72549 , n73014 );
or ( n73016 , n72548 , n73015 );
and ( n73017 , n72545 , n73016 );
or ( n73018 , n72544 , n73017 );
and ( n73019 , n72541 , n73018 );
or ( n73020 , n72540 , n73019 );
and ( n73021 , n72537 , n73020 );
or ( n73022 , n72536 , n73021 );
and ( n73023 , n72533 , n73022 );
or ( n73024 , n72532 , n73023 );
and ( n73025 , n72529 , n73024 );
or ( n73026 , n72528 , n73025 );
and ( n73027 , n72525 , n73026 );
or ( n73028 , n72524 , n73027 );
and ( n73029 , n72521 , n73028 );
or ( n73030 , n72520 , n73029 );
and ( n73031 , n72517 , n73030 );
or ( n73032 , n72516 , n73031 );
and ( n73033 , n72513 , n73032 );
or ( n73034 , n72512 , n73033 );
and ( n73035 , n72509 , n73034 );
or ( n73036 , n72508 , n73035 );
and ( n73037 , n72505 , n73036 );
or ( n73038 , n72504 , n73037 );
and ( n73039 , n72501 , n73038 );
or ( n73040 , n72500 , n73039 );
and ( n73041 , n72497 , n73040 );
or ( n73042 , n72496 , n73041 );
and ( n73043 , n72493 , n73042 );
or ( n73044 , n72492 , n73043 );
and ( n73045 , n72489 , n73044 );
or ( n73046 , n72488 , n73045 );
xor ( n73047 , n72485 , n73046 );
and ( n73048 , n33403 , n7412 );
nor ( n73049 , n7413 , n73048 );
nor ( n73050 , n7841 , n32231 );
xor ( n73051 , n73049 , n73050 );
and ( n73052 , n71863 , n71864 );
and ( n73053 , n71865 , n71868 );
or ( n73054 , n73052 , n73053 );
xor ( n73055 , n73051 , n73054 );
nor ( n73056 , n8281 , n31083 );
xor ( n73057 , n73055 , n73056 );
and ( n73058 , n71869 , n71870 );
and ( n73059 , n71871 , n71874 );
or ( n73060 , n73058 , n73059 );
xor ( n73061 , n73057 , n73060 );
nor ( n73062 , n8737 , n29948 );
xor ( n73063 , n73061 , n73062 );
and ( n73064 , n71875 , n71876 );
and ( n73065 , n71877 , n71880 );
or ( n73066 , n73064 , n73065 );
xor ( n73067 , n73063 , n73066 );
nor ( n73068 , n9420 , n28833 );
xor ( n73069 , n73067 , n73068 );
and ( n73070 , n71881 , n71882 );
and ( n73071 , n71883 , n71886 );
or ( n73072 , n73070 , n73071 );
xor ( n73073 , n73069 , n73072 );
nor ( n73074 , n10312 , n27737 );
xor ( n73075 , n73073 , n73074 );
and ( n73076 , n71887 , n71888 );
and ( n73077 , n71889 , n71892 );
or ( n73078 , n73076 , n73077 );
xor ( n73079 , n73075 , n73078 );
nor ( n73080 , n11041 , n26660 );
xor ( n73081 , n73079 , n73080 );
and ( n73082 , n71893 , n71894 );
and ( n73083 , n71895 , n71898 );
or ( n73084 , n73082 , n73083 );
xor ( n73085 , n73081 , n73084 );
nor ( n73086 , n11790 , n25600 );
xor ( n73087 , n73085 , n73086 );
and ( n73088 , n71899 , n71900 );
and ( n73089 , n71901 , n71904 );
or ( n73090 , n73088 , n73089 );
xor ( n73091 , n73087 , n73090 );
nor ( n73092 , n12555 , n24564 );
xor ( n73093 , n73091 , n73092 );
and ( n73094 , n71905 , n71906 );
and ( n73095 , n71907 , n71910 );
or ( n73096 , n73094 , n73095 );
xor ( n73097 , n73093 , n73096 );
nor ( n73098 , n13340 , n23541 );
xor ( n73099 , n73097 , n73098 );
and ( n73100 , n71911 , n71912 );
and ( n73101 , n71913 , n71916 );
or ( n73102 , n73100 , n73101 );
xor ( n73103 , n73099 , n73102 );
nor ( n73104 , n14138 , n22541 );
xor ( n73105 , n73103 , n73104 );
and ( n73106 , n71917 , n71918 );
and ( n73107 , n71919 , n71922 );
or ( n73108 , n73106 , n73107 );
xor ( n73109 , n73105 , n73108 );
nor ( n73110 , n14959 , n21562 );
xor ( n73111 , n73109 , n73110 );
and ( n73112 , n71923 , n71924 );
and ( n73113 , n71925 , n71928 );
or ( n73114 , n73112 , n73113 );
xor ( n73115 , n73111 , n73114 );
nor ( n73116 , n15800 , n20601 );
xor ( n73117 , n73115 , n73116 );
and ( n73118 , n71929 , n71930 );
and ( n73119 , n71931 , n71934 );
or ( n73120 , n73118 , n73119 );
xor ( n73121 , n73117 , n73120 );
nor ( n73122 , n16660 , n19657 );
xor ( n73123 , n73121 , n73122 );
and ( n73124 , n71935 , n71936 );
and ( n73125 , n71937 , n71940 );
or ( n73126 , n73124 , n73125 );
xor ( n73127 , n73123 , n73126 );
nor ( n73128 , n17539 , n18734 );
xor ( n73129 , n73127 , n73128 );
and ( n73130 , n71941 , n71942 );
and ( n73131 , n71943 , n71946 );
or ( n73132 , n73130 , n73131 );
xor ( n73133 , n73129 , n73132 );
nor ( n73134 , n18439 , n17828 );
xor ( n73135 , n73133 , n73134 );
and ( n73136 , n71947 , n71948 );
and ( n73137 , n71949 , n71952 );
or ( n73138 , n73136 , n73137 );
xor ( n73139 , n73135 , n73138 );
nor ( n73140 , n19356 , n16943 );
xor ( n73141 , n73139 , n73140 );
and ( n73142 , n71953 , n71954 );
and ( n73143 , n71955 , n71958 );
or ( n73144 , n73142 , n73143 );
xor ( n73145 , n73141 , n73144 );
nor ( n73146 , n20294 , n16077 );
xor ( n73147 , n73145 , n73146 );
and ( n73148 , n71959 , n71960 );
and ( n73149 , n71961 , n71964 );
or ( n73150 , n73148 , n73149 );
xor ( n73151 , n73147 , n73150 );
nor ( n73152 , n21249 , n15230 );
xor ( n73153 , n73151 , n73152 );
and ( n73154 , n71965 , n71966 );
and ( n73155 , n71967 , n71970 );
or ( n73156 , n73154 , n73155 );
xor ( n73157 , n73153 , n73156 );
nor ( n73158 , n22222 , n14403 );
xor ( n73159 , n73157 , n73158 );
and ( n73160 , n71971 , n71972 );
and ( n73161 , n71973 , n71976 );
or ( n73162 , n73160 , n73161 );
xor ( n73163 , n73159 , n73162 );
nor ( n73164 , n23216 , n13599 );
xor ( n73165 , n73163 , n73164 );
and ( n73166 , n71977 , n71978 );
and ( n73167 , n71979 , n71982 );
or ( n73168 , n73166 , n73167 );
xor ( n73169 , n73165 , n73168 );
nor ( n73170 , n24233 , n12808 );
xor ( n73171 , n73169 , n73170 );
and ( n73172 , n71983 , n71984 );
and ( n73173 , n71985 , n71988 );
or ( n73174 , n73172 , n73173 );
xor ( n73175 , n73171 , n73174 );
nor ( n73176 , n25263 , n12037 );
xor ( n73177 , n73175 , n73176 );
and ( n73178 , n71989 , n71990 );
and ( n73179 , n71991 , n71994 );
or ( n73180 , n73178 , n73179 );
xor ( n73181 , n73177 , n73180 );
nor ( n73182 , n26317 , n11282 );
xor ( n73183 , n73181 , n73182 );
and ( n73184 , n71995 , n71996 );
and ( n73185 , n71997 , n72000 );
or ( n73186 , n73184 , n73185 );
xor ( n73187 , n73183 , n73186 );
nor ( n73188 , n27388 , n10547 );
xor ( n73189 , n73187 , n73188 );
and ( n73190 , n72001 , n72002 );
and ( n73191 , n72003 , n72006 );
or ( n73192 , n73190 , n73191 );
xor ( n73193 , n73189 , n73192 );
nor ( n73194 , n28478 , n9829 );
xor ( n73195 , n73193 , n73194 );
and ( n73196 , n72007 , n72008 );
and ( n73197 , n72009 , n72012 );
or ( n73198 , n73196 , n73197 );
xor ( n73199 , n73195 , n73198 );
nor ( n73200 , n29587 , n8955 );
xor ( n73201 , n73199 , n73200 );
and ( n73202 , n72013 , n72014 );
and ( n73203 , n72015 , n72018 );
or ( n73204 , n73202 , n73203 );
xor ( n73205 , n73201 , n73204 );
nor ( n73206 , n30716 , n603 );
xor ( n73207 , n73205 , n73206 );
and ( n73208 , n72019 , n72020 );
and ( n73209 , n72021 , n72024 );
or ( n73210 , n73208 , n73209 );
xor ( n73211 , n73207 , n73210 );
nor ( n73212 , n31858 , n652 );
xor ( n73213 , n73211 , n73212 );
and ( n73214 , n72025 , n72026 );
and ( n73215 , n72027 , n72030 );
or ( n73216 , n73214 , n73215 );
xor ( n73217 , n73213 , n73216 );
nor ( n73218 , n33024 , n624 );
xor ( n73219 , n73217 , n73218 );
and ( n73220 , n72031 , n72032 );
and ( n73221 , n72033 , n72036 );
or ( n73222 , n73220 , n73221 );
xor ( n73223 , n73219 , n73222 );
nor ( n73224 , n34215 , n648 );
xor ( n73225 , n73223 , n73224 );
and ( n73226 , n72037 , n72038 );
and ( n73227 , n72039 , n72042 );
or ( n73228 , n73226 , n73227 );
xor ( n73229 , n73225 , n73228 );
nor ( n73230 , n35410 , n686 );
xor ( n73231 , n73229 , n73230 );
and ( n73232 , n72043 , n72044 );
and ( n73233 , n72045 , n72048 );
or ( n73234 , n73232 , n73233 );
xor ( n73235 , n73231 , n73234 );
nor ( n73236 , n36611 , n735 );
xor ( n73237 , n73235 , n73236 );
and ( n73238 , n72049 , n72050 );
and ( n73239 , n72051 , n72054 );
or ( n73240 , n73238 , n73239 );
xor ( n73241 , n73237 , n73240 );
nor ( n73242 , n37816 , n798 );
xor ( n73243 , n73241 , n73242 );
and ( n73244 , n72055 , n72056 );
and ( n73245 , n72057 , n72060 );
or ( n73246 , n73244 , n73245 );
xor ( n73247 , n73243 , n73246 );
nor ( n73248 , n39018 , n870 );
xor ( n73249 , n73247 , n73248 );
and ( n73250 , n72061 , n72062 );
and ( n73251 , n72063 , n72066 );
or ( n73252 , n73250 , n73251 );
xor ( n73253 , n73249 , n73252 );
nor ( n73254 , n40223 , n960 );
xor ( n73255 , n73253 , n73254 );
and ( n73256 , n72067 , n72068 );
and ( n73257 , n72069 , n72072 );
or ( n73258 , n73256 , n73257 );
xor ( n73259 , n73255 , n73258 );
nor ( n73260 , n41428 , n1064 );
xor ( n73261 , n73259 , n73260 );
and ( n73262 , n72073 , n72074 );
and ( n73263 , n72075 , n72078 );
or ( n73264 , n73262 , n73263 );
xor ( n73265 , n73261 , n73264 );
nor ( n73266 , n42632 , n1178 );
xor ( n73267 , n73265 , n73266 );
and ( n73268 , n72079 , n72080 );
and ( n73269 , n72081 , n72084 );
or ( n73270 , n73268 , n73269 );
xor ( n73271 , n73267 , n73270 );
nor ( n73272 , n43834 , n1305 );
xor ( n73273 , n73271 , n73272 );
and ( n73274 , n72085 , n72086 );
and ( n73275 , n72087 , n72090 );
or ( n73276 , n73274 , n73275 );
xor ( n73277 , n73273 , n73276 );
nor ( n73278 , n45038 , n1447 );
xor ( n73279 , n73277 , n73278 );
and ( n73280 , n72091 , n72092 );
and ( n73281 , n72093 , n72096 );
or ( n73282 , n73280 , n73281 );
xor ( n73283 , n73279 , n73282 );
nor ( n73284 , n46239 , n1600 );
xor ( n73285 , n73283 , n73284 );
and ( n73286 , n72097 , n72098 );
and ( n73287 , n72099 , n72102 );
or ( n73288 , n73286 , n73287 );
xor ( n73289 , n73285 , n73288 );
nor ( n73290 , n47440 , n1768 );
xor ( n73291 , n73289 , n73290 );
and ( n73292 , n72103 , n72104 );
and ( n73293 , n72105 , n72108 );
or ( n73294 , n73292 , n73293 );
xor ( n73295 , n73291 , n73294 );
nor ( n73296 , n48641 , n1947 );
xor ( n73297 , n73295 , n73296 );
and ( n73298 , n72109 , n72110 );
and ( n73299 , n72111 , n72114 );
or ( n73300 , n73298 , n73299 );
xor ( n73301 , n73297 , n73300 );
nor ( n73302 , n49841 , n2139 );
xor ( n73303 , n73301 , n73302 );
and ( n73304 , n72115 , n72116 );
and ( n73305 , n72117 , n72120 );
or ( n73306 , n73304 , n73305 );
xor ( n73307 , n73303 , n73306 );
nor ( n73308 , n51040 , n2345 );
xor ( n73309 , n73307 , n73308 );
and ( n73310 , n72121 , n72122 );
and ( n73311 , n72123 , n72126 );
or ( n73312 , n73310 , n73311 );
xor ( n73313 , n73309 , n73312 );
nor ( n73314 , n52238 , n2568 );
xor ( n73315 , n73313 , n73314 );
and ( n73316 , n72127 , n72128 );
and ( n73317 , n72129 , n72132 );
or ( n73318 , n73316 , n73317 );
xor ( n73319 , n73315 , n73318 );
nor ( n73320 , n53432 , n2799 );
xor ( n73321 , n73319 , n73320 );
and ( n73322 , n72133 , n72134 );
and ( n73323 , n72135 , n72138 );
or ( n73324 , n73322 , n73323 );
xor ( n73325 , n73321 , n73324 );
nor ( n73326 , n54629 , n3045 );
xor ( n73327 , n73325 , n73326 );
and ( n73328 , n72139 , n72140 );
and ( n73329 , n72141 , n72144 );
or ( n73330 , n73328 , n73329 );
xor ( n73331 , n73327 , n73330 );
nor ( n73332 , n55826 , n3302 );
xor ( n73333 , n73331 , n73332 );
and ( n73334 , n72145 , n72146 );
and ( n73335 , n72147 , n72150 );
or ( n73336 , n73334 , n73335 );
xor ( n73337 , n73333 , n73336 );
nor ( n73338 , n57022 , n3572 );
xor ( n73339 , n73337 , n73338 );
and ( n73340 , n72151 , n72152 );
and ( n73341 , n72153 , n72156 );
or ( n73342 , n73340 , n73341 );
xor ( n73343 , n73339 , n73342 );
nor ( n73344 , n58217 , n3855 );
xor ( n73345 , n73343 , n73344 );
and ( n73346 , n72157 , n72158 );
and ( n73347 , n72159 , n72162 );
or ( n73348 , n73346 , n73347 );
xor ( n73349 , n73345 , n73348 );
nor ( n73350 , n59412 , n4153 );
xor ( n73351 , n73349 , n73350 );
and ( n73352 , n72163 , n72164 );
and ( n73353 , n72165 , n72168 );
or ( n73354 , n73352 , n73353 );
xor ( n73355 , n73351 , n73354 );
nor ( n73356 , n60600 , n4460 );
xor ( n73357 , n73355 , n73356 );
and ( n73358 , n72169 , n72170 );
and ( n73359 , n72171 , n72174 );
or ( n73360 , n73358 , n73359 );
xor ( n73361 , n73357 , n73360 );
nor ( n73362 , n61791 , n4788 );
xor ( n73363 , n73361 , n73362 );
and ( n73364 , n72175 , n72176 );
and ( n73365 , n72177 , n72180 );
or ( n73366 , n73364 , n73365 );
xor ( n73367 , n73363 , n73366 );
nor ( n73368 , n62982 , n5128 );
xor ( n73369 , n73367 , n73368 );
and ( n73370 , n72181 , n72182 );
and ( n73371 , n72183 , n72186 );
or ( n73372 , n73370 , n73371 );
xor ( n73373 , n73369 , n73372 );
nor ( n73374 , n64172 , n5479 );
xor ( n73375 , n73373 , n73374 );
and ( n73376 , n72187 , n72188 );
and ( n73377 , n72189 , n72192 );
or ( n73378 , n73376 , n73377 );
xor ( n73379 , n73375 , n73378 );
nor ( n73380 , n65360 , n5840 );
xor ( n73381 , n73379 , n73380 );
and ( n73382 , n72193 , n72194 );
and ( n73383 , n72195 , n72198 );
or ( n73384 , n73382 , n73383 );
xor ( n73385 , n73381 , n73384 );
nor ( n73386 , n66550 , n6214 );
xor ( n73387 , n73385 , n73386 );
and ( n73388 , n72199 , n72200 );
and ( n73389 , n72201 , n72204 );
or ( n73390 , n73388 , n73389 );
xor ( n73391 , n73387 , n73390 );
nor ( n73392 , n67736 , n6598 );
xor ( n73393 , n73391 , n73392 );
and ( n73394 , n72205 , n72206 );
and ( n73395 , n72207 , n72210 );
or ( n73396 , n73394 , n73395 );
xor ( n73397 , n73393 , n73396 );
nor ( n73398 , n68924 , n6999 );
xor ( n73399 , n73397 , n73398 );
and ( n73400 , n72211 , n72212 );
and ( n73401 , n72213 , n72216 );
or ( n73402 , n73400 , n73401 );
xor ( n73403 , n73399 , n73402 );
nor ( n73404 , n70110 , n7415 );
xor ( n73405 , n73403 , n73404 );
and ( n73406 , n72217 , n72218 );
and ( n73407 , n72219 , n72222 );
or ( n73408 , n73406 , n73407 );
xor ( n73409 , n73405 , n73408 );
nor ( n73410 , n71292 , n7843 );
xor ( n73411 , n73409 , n73410 );
and ( n73412 , n72223 , n72224 );
and ( n73413 , n72225 , n72228 );
or ( n73414 , n73412 , n73413 );
xor ( n73415 , n73411 , n73414 );
nor ( n73416 , n72472 , n8283 );
xor ( n73417 , n73415 , n73416 );
and ( n73418 , n72229 , n72230 );
and ( n73419 , n72231 , n72234 );
or ( n73420 , n73418 , n73419 );
xor ( n73421 , n73417 , n73420 );
and ( n73422 , n72247 , n72251 );
and ( n73423 , n72251 , n72458 );
and ( n73424 , n72247 , n72458 );
or ( n73425 , n73422 , n73423 , n73424 );
and ( n73426 , n33774 , n7310 );
not ( n73427 , n7310 );
nor ( n73428 , n73426 , n73427 );
xor ( n73429 , n73425 , n73428 );
and ( n73430 , n72257 , n72258 );
and ( n73431 , n72258 , n72326 );
and ( n73432 , n72257 , n72326 );
or ( n73433 , n73430 , n73431 , n73432 );
and ( n73434 , n72253 , n72327 );
and ( n73435 , n72327 , n72457 );
and ( n73436 , n72253 , n72457 );
or ( n73437 , n73434 , n73435 , n73436 );
xor ( n73438 , n73433 , n73437 );
and ( n73439 , n72344 , n72456 );
and ( n73440 , n72263 , n72267 );
and ( n73441 , n72267 , n72325 );
and ( n73442 , n72263 , n72325 );
or ( n73443 , n73440 , n73441 , n73442 );
and ( n73444 , n72348 , n72455 );
xor ( n73445 , n73443 , n73444 );
and ( n73446 , n72294 , n72298 );
and ( n73447 , n72298 , n72304 );
and ( n73448 , n72294 , n72304 );
or ( n73449 , n73446 , n73447 , n73448 );
and ( n73450 , n72272 , n72276 );
and ( n73451 , n72276 , n72324 );
and ( n73452 , n72272 , n72324 );
or ( n73453 , n73450 , n73451 , n73452 );
xor ( n73454 , n73449 , n73453 );
and ( n73455 , n72281 , n72285 );
and ( n73456 , n72285 , n72323 );
and ( n73457 , n72281 , n72323 );
or ( n73458 , n73455 , n73456 , n73457 );
and ( n73459 , n72356 , n72381 );
and ( n73460 , n72381 , n72419 );
and ( n73461 , n72356 , n72419 );
or ( n73462 , n73459 , n73460 , n73461 );
xor ( n73463 , n73458 , n73462 );
and ( n73464 , n72290 , n72305 );
and ( n73465 , n72305 , n72322 );
and ( n73466 , n72290 , n72322 );
or ( n73467 , n73464 , n73465 , n73466 );
and ( n73468 , n72360 , n72364 );
and ( n73469 , n72364 , n72380 );
and ( n73470 , n72360 , n72380 );
or ( n73471 , n73468 , n73469 , n73470 );
xor ( n73472 , n73467 , n73471 );
and ( n73473 , n72310 , n72315 );
and ( n73474 , n72315 , n72321 );
and ( n73475 , n72310 , n72321 );
or ( n73476 , n73473 , n73474 , n73475 );
and ( n73477 , n72300 , n72301 );
and ( n73478 , n72301 , n72303 );
and ( n73479 , n72300 , n72303 );
or ( n73480 , n73477 , n73478 , n73479 );
and ( n73481 , n72311 , n72312 );
and ( n73482 , n72312 , n72314 );
and ( n73483 , n72311 , n72314 );
or ( n73484 , n73481 , n73482 , n73483 );
xor ( n73485 , n73480 , n73484 );
and ( n73486 , n30695 , n8669 );
and ( n73487 , n31836 , n8243 );
xor ( n73488 , n73486 , n73487 );
and ( n73489 , n32649 , n7662 );
xor ( n73490 , n73488 , n73489 );
xor ( n73491 , n73485 , n73490 );
xor ( n73492 , n73476 , n73491 );
and ( n73493 , n72317 , n72318 );
and ( n73494 , n72318 , n72320 );
and ( n73495 , n72317 , n72320 );
or ( n73496 , n73493 , n73494 , n73495 );
and ( n73497 , n27361 , n10977 );
and ( n73498 , n28456 , n10239 );
xor ( n73499 , n73497 , n73498 );
and ( n73500 , n29559 , n9348 );
xor ( n73501 , n73499 , n73500 );
xor ( n73502 , n73496 , n73501 );
and ( n73503 , n24214 , n13256 );
and ( n73504 , n25243 , n12531 );
xor ( n73505 , n73503 , n73504 );
and ( n73506 , n26296 , n11718 );
xor ( n73507 , n73505 , n73506 );
xor ( n73508 , n73502 , n73507 );
xor ( n73509 , n73492 , n73508 );
xor ( n73510 , n73472 , n73509 );
xor ( n73511 , n73463 , n73510 );
xor ( n73512 , n73454 , n73511 );
xor ( n73513 , n73445 , n73512 );
xor ( n73514 , n73439 , n73513 );
and ( n73515 , n72338 , n72339 );
and ( n73516 , n72339 , n72341 );
and ( n73517 , n72338 , n72341 );
or ( n73518 , n73515 , n73516 , n73517 );
not ( n73519 , n7385 );
and ( n73520 , n34193 , n7385 );
nor ( n73521 , n73519 , n73520 );
and ( n73522 , n7808 , n32999 );
xor ( n73523 , n73521 , n73522 );
and ( n73524 , n8079 , n31761 );
xor ( n73525 , n73523 , n73524 );
xor ( n73526 , n73518 , n73525 );
and ( n73527 , n72352 , n72420 );
and ( n73528 , n72420 , n72454 );
and ( n73529 , n72352 , n72454 );
or ( n73530 , n73527 , n73528 , n73529 );
and ( n73531 , n72425 , n72426 );
and ( n73532 , n72426 , n72453 );
and ( n73533 , n72425 , n72453 );
or ( n73534 , n73531 , n73532 , n73533 );
and ( n73535 , n72386 , n72402 );
and ( n73536 , n72402 , n72418 );
and ( n73537 , n72386 , n72418 );
or ( n73538 , n73535 , n73536 , n73537 );
and ( n73539 , n72369 , n72373 );
and ( n73540 , n72373 , n72379 );
and ( n73541 , n72369 , n72379 );
or ( n73542 , n73539 , n73540 , n73541 );
and ( n73543 , n72390 , n72395 );
and ( n73544 , n72395 , n72401 );
and ( n73545 , n72390 , n72401 );
or ( n73546 , n73543 , n73544 , n73545 );
xor ( n73547 , n73542 , n73546 );
and ( n73548 , n72375 , n72376 );
and ( n73549 , n72376 , n72378 );
and ( n73550 , n72375 , n72378 );
or ( n73551 , n73548 , n73549 , n73550 );
and ( n73552 , n72391 , n72392 );
and ( n73553 , n72392 , n72394 );
and ( n73554 , n72391 , n72394 );
or ( n73555 , n73552 , n73553 , n73554 );
xor ( n73556 , n73551 , n73555 );
and ( n73557 , n21216 , n15691 );
and ( n73558 , n22186 , n14838 );
xor ( n73559 , n73557 , n73558 );
and ( n73560 , n22892 , n14044 );
xor ( n73561 , n73559 , n73560 );
xor ( n73562 , n73556 , n73561 );
xor ( n73563 , n73547 , n73562 );
xor ( n73564 , n73538 , n73563 );
and ( n73565 , n72407 , n72411 );
and ( n73566 , n72411 , n72417 );
and ( n73567 , n72407 , n72417 );
or ( n73568 , n73565 , n73566 , n73567 );
and ( n73569 , n72397 , n72398 );
and ( n73570 , n72398 , n72400 );
and ( n73571 , n72397 , n72400 );
or ( n73572 , n73569 , n73570 , n73571 );
buf ( n73573 , n18144 );
and ( n73574 , n19324 , n17422 );
xor ( n73575 , n73573 , n73574 );
and ( n73576 , n20233 , n16550 );
xor ( n73577 , n73575 , n73576 );
xor ( n73578 , n73572 , n73577 );
and ( n73579 , n15758 , n20976 );
and ( n73580 , n16637 , n20156 );
xor ( n73581 , n73579 , n73580 );
and ( n73582 , n17512 , n19222 );
xor ( n73583 , n73581 , n73582 );
xor ( n73584 , n73578 , n73583 );
xor ( n73585 , n73568 , n73584 );
and ( n73586 , n72413 , n72414 );
and ( n73587 , n72414 , n72416 );
and ( n73588 , n72413 , n72416 );
or ( n73589 , n73586 , n73587 , n73588 );
and ( n73590 , n72441 , n72442 );
and ( n73591 , n72442 , n72444 );
and ( n73592 , n72441 , n72444 );
or ( n73593 , n73590 , n73591 , n73592 );
xor ( n73594 , n73589 , n73593 );
and ( n73595 , n13322 , n24137 );
and ( n73596 , n14118 , n23075 );
xor ( n73597 , n73595 , n73596 );
and ( n73598 , n14938 , n22065 );
xor ( n73599 , n73597 , n73598 );
xor ( n73600 , n73594 , n73599 );
xor ( n73601 , n73585 , n73600 );
xor ( n73602 , n73564 , n73601 );
xor ( n73603 , n73534 , n73602 );
and ( n73604 , n72431 , n72435 );
and ( n73605 , n72435 , n72452 );
and ( n73606 , n72431 , n72452 );
or ( n73607 , n73604 , n73605 , n73606 );
and ( n73608 , n72331 , n72343 );
xor ( n73609 , n73607 , n73608 );
and ( n73610 , n72335 , n72336 );
and ( n73611 , n72336 , n72342 );
and ( n73612 , n72335 , n72342 );
or ( n73613 , n73610 , n73611 , n73612 );
and ( n73614 , n72440 , n72445 );
and ( n73615 , n72445 , n72451 );
and ( n73616 , n72440 , n72451 );
or ( n73617 , n73614 , n73615 , n73616 );
xor ( n73618 , n73613 , n73617 );
and ( n73619 , n72447 , n72448 );
and ( n73620 , n72448 , n72450 );
and ( n73621 , n72447 , n72450 );
or ( n73622 , n73619 , n73620 , n73621 );
and ( n73623 , n11015 , n27296 );
and ( n73624 , n11769 , n26216 );
xor ( n73625 , n73623 , n73624 );
and ( n73626 , n12320 , n25163 );
xor ( n73627 , n73625 , n73626 );
xor ( n73628 , n73622 , n73627 );
and ( n73629 , n8718 , n30629 );
and ( n73630 , n9400 , n29508 );
xor ( n73631 , n73629 , n73630 );
and ( n73632 , n10291 , n28406 );
xor ( n73633 , n73631 , n73632 );
xor ( n73634 , n73628 , n73633 );
xor ( n73635 , n73618 , n73634 );
xor ( n73636 , n73609 , n73635 );
xor ( n73637 , n73603 , n73636 );
xor ( n73638 , n73530 , n73637 );
xor ( n73639 , n73526 , n73638 );
xor ( n73640 , n73514 , n73639 );
xor ( n73641 , n73438 , n73640 );
xor ( n73642 , n73429 , n73641 );
and ( n73643 , n72239 , n72242 );
and ( n73644 , n72242 , n72459 );
and ( n73645 , n72239 , n72459 );
or ( n73646 , n73643 , n73644 , n73645 );
xor ( n73647 , n73642 , n73646 );
and ( n73648 , n72460 , n72464 );
and ( n73649 , n72465 , n72468 );
or ( n73650 , n73648 , n73649 );
xor ( n73651 , n73647 , n73650 );
buf ( n73652 , n73651 );
buf ( n73653 , n73652 );
not ( n73654 , n73653 );
nor ( n73655 , n73654 , n8739 );
xor ( n73656 , n73421 , n73655 );
and ( n73657 , n72235 , n72473 );
and ( n73658 , n72474 , n72477 );
or ( n73659 , n73657 , n73658 );
xor ( n73660 , n73656 , n73659 );
buf ( n73661 , n73660 );
buf ( n73662 , n73661 );
not ( n73663 , n73662 );
buf ( n73664 , n595 );
not ( n73665 , n73664 );
nor ( n73666 , n73663 , n73665 );
xor ( n73667 , n73047 , n73666 );
xor ( n73668 , n72489 , n73044 );
nor ( n73669 , n72481 , n73665 );
and ( n73670 , n73668 , n73669 );
xor ( n73671 , n73668 , n73669 );
xor ( n73672 , n72493 , n73042 );
nor ( n73673 , n71301 , n73665 );
and ( n73674 , n73672 , n73673 );
xor ( n73675 , n73672 , n73673 );
xor ( n73676 , n72497 , n73040 );
nor ( n73677 , n70119 , n73665 );
and ( n73678 , n73676 , n73677 );
xor ( n73679 , n73676 , n73677 );
xor ( n73680 , n72501 , n73038 );
nor ( n73681 , n68933 , n73665 );
and ( n73682 , n73680 , n73681 );
xor ( n73683 , n73680 , n73681 );
xor ( n73684 , n72505 , n73036 );
nor ( n73685 , n67745 , n73665 );
and ( n73686 , n73684 , n73685 );
xor ( n73687 , n73684 , n73685 );
xor ( n73688 , n72509 , n73034 );
nor ( n73689 , n66559 , n73665 );
and ( n73690 , n73688 , n73689 );
xor ( n73691 , n73688 , n73689 );
xor ( n73692 , n72513 , n73032 );
nor ( n73693 , n65369 , n73665 );
and ( n73694 , n73692 , n73693 );
xor ( n73695 , n73692 , n73693 );
xor ( n73696 , n72517 , n73030 );
nor ( n73697 , n64181 , n73665 );
and ( n73698 , n73696 , n73697 );
xor ( n73699 , n73696 , n73697 );
xor ( n73700 , n72521 , n73028 );
nor ( n73701 , n62991 , n73665 );
and ( n73702 , n73700 , n73701 );
xor ( n73703 , n73700 , n73701 );
xor ( n73704 , n72525 , n73026 );
nor ( n73705 , n61800 , n73665 );
and ( n73706 , n73704 , n73705 );
xor ( n73707 , n73704 , n73705 );
xor ( n73708 , n72529 , n73024 );
nor ( n73709 , n60609 , n73665 );
and ( n73710 , n73708 , n73709 );
xor ( n73711 , n73708 , n73709 );
xor ( n73712 , n72533 , n73022 );
nor ( n73713 , n59421 , n73665 );
and ( n73714 , n73712 , n73713 );
xor ( n73715 , n73712 , n73713 );
xor ( n73716 , n72537 , n73020 );
nor ( n73717 , n58226 , n73665 );
and ( n73718 , n73716 , n73717 );
xor ( n73719 , n73716 , n73717 );
xor ( n73720 , n72541 , n73018 );
nor ( n73721 , n57031 , n73665 );
and ( n73722 , n73720 , n73721 );
xor ( n73723 , n73720 , n73721 );
xor ( n73724 , n72545 , n73016 );
nor ( n73725 , n55835 , n73665 );
and ( n73726 , n73724 , n73725 );
xor ( n73727 , n73724 , n73725 );
xor ( n73728 , n72549 , n73014 );
nor ( n73729 , n54638 , n73665 );
and ( n73730 , n73728 , n73729 );
xor ( n73731 , n73728 , n73729 );
xor ( n73732 , n72553 , n73012 );
nor ( n73733 , n53441 , n73665 );
and ( n73734 , n73732 , n73733 );
xor ( n73735 , n73732 , n73733 );
xor ( n73736 , n72557 , n73010 );
nor ( n73737 , n52247 , n73665 );
and ( n73738 , n73736 , n73737 );
xor ( n73739 , n73736 , n73737 );
xor ( n73740 , n72561 , n73008 );
nor ( n73741 , n51049 , n73665 );
and ( n73742 , n73740 , n73741 );
xor ( n73743 , n73740 , n73741 );
xor ( n73744 , n72565 , n73006 );
nor ( n73745 , n49850 , n73665 );
and ( n73746 , n73744 , n73745 );
xor ( n73747 , n73744 , n73745 );
xor ( n73748 , n72569 , n73004 );
nor ( n73749 , n48650 , n73665 );
and ( n73750 , n73748 , n73749 );
xor ( n73751 , n73748 , n73749 );
xor ( n73752 , n72573 , n73002 );
nor ( n73753 , n47449 , n73665 );
and ( n73754 , n73752 , n73753 );
xor ( n73755 , n73752 , n73753 );
xor ( n73756 , n72577 , n73000 );
nor ( n73757 , n46248 , n73665 );
and ( n73758 , n73756 , n73757 );
xor ( n73759 , n73756 , n73757 );
xor ( n73760 , n72581 , n72998 );
nor ( n73761 , n45047 , n73665 );
and ( n73762 , n73760 , n73761 );
xor ( n73763 , n73760 , n73761 );
xor ( n73764 , n72585 , n72996 );
nor ( n73765 , n43843 , n73665 );
and ( n73766 , n73764 , n73765 );
xor ( n73767 , n73764 , n73765 );
xor ( n73768 , n72589 , n72994 );
nor ( n73769 , n42641 , n73665 );
and ( n73770 , n73768 , n73769 );
xor ( n73771 , n73768 , n73769 );
xor ( n73772 , n72593 , n72992 );
nor ( n73773 , n41437 , n73665 );
and ( n73774 , n73772 , n73773 );
xor ( n73775 , n73772 , n73773 );
xor ( n73776 , n72597 , n72990 );
nor ( n73777 , n40232 , n73665 );
and ( n73778 , n73776 , n73777 );
xor ( n73779 , n73776 , n73777 );
xor ( n73780 , n72601 , n72988 );
nor ( n73781 , n39027 , n73665 );
and ( n73782 , n73780 , n73781 );
xor ( n73783 , n73780 , n73781 );
xor ( n73784 , n72605 , n72986 );
nor ( n73785 , n37825 , n73665 );
and ( n73786 , n73784 , n73785 );
xor ( n73787 , n73784 , n73785 );
xor ( n73788 , n72609 , n72984 );
nor ( n73789 , n36620 , n73665 );
and ( n73790 , n73788 , n73789 );
xor ( n73791 , n73788 , n73789 );
xor ( n73792 , n72613 , n72982 );
nor ( n73793 , n35419 , n73665 );
and ( n73794 , n73792 , n73793 );
xor ( n73795 , n73792 , n73793 );
xor ( n73796 , n72617 , n72980 );
nor ( n73797 , n34224 , n73665 );
and ( n73798 , n73796 , n73797 );
xor ( n73799 , n73796 , n73797 );
xor ( n73800 , n72621 , n72978 );
nor ( n73801 , n33033 , n73665 );
and ( n73802 , n73800 , n73801 );
xor ( n73803 , n73800 , n73801 );
xor ( n73804 , n72625 , n72976 );
nor ( n73805 , n31867 , n73665 );
and ( n73806 , n73804 , n73805 );
xor ( n73807 , n73804 , n73805 );
xor ( n73808 , n72629 , n72974 );
nor ( n73809 , n30725 , n73665 );
and ( n73810 , n73808 , n73809 );
xor ( n73811 , n73808 , n73809 );
xor ( n73812 , n72633 , n72972 );
nor ( n73813 , n29596 , n73665 );
and ( n73814 , n73812 , n73813 );
xor ( n73815 , n73812 , n73813 );
xor ( n73816 , n72637 , n72970 );
nor ( n73817 , n28487 , n73665 );
and ( n73818 , n73816 , n73817 );
xor ( n73819 , n73816 , n73817 );
xor ( n73820 , n72641 , n72968 );
nor ( n73821 , n27397 , n73665 );
and ( n73822 , n73820 , n73821 );
xor ( n73823 , n73820 , n73821 );
xor ( n73824 , n72645 , n72966 );
nor ( n73825 , n26326 , n73665 );
and ( n73826 , n73824 , n73825 );
xor ( n73827 , n73824 , n73825 );
xor ( n73828 , n72649 , n72964 );
nor ( n73829 , n25272 , n73665 );
and ( n73830 , n73828 , n73829 );
xor ( n73831 , n73828 , n73829 );
xor ( n73832 , n72653 , n72962 );
nor ( n73833 , n24242 , n73665 );
and ( n73834 , n73832 , n73833 );
xor ( n73835 , n73832 , n73833 );
xor ( n73836 , n72657 , n72960 );
nor ( n73837 , n23225 , n73665 );
and ( n73838 , n73836 , n73837 );
xor ( n73839 , n73836 , n73837 );
xor ( n73840 , n72661 , n72958 );
nor ( n73841 , n22231 , n73665 );
and ( n73842 , n73840 , n73841 );
xor ( n73843 , n73840 , n73841 );
xor ( n73844 , n72665 , n72956 );
nor ( n73845 , n21258 , n73665 );
and ( n73846 , n73844 , n73845 );
xor ( n73847 , n73844 , n73845 );
xor ( n73848 , n72669 , n72954 );
nor ( n73849 , n20303 , n73665 );
and ( n73850 , n73848 , n73849 );
xor ( n73851 , n73848 , n73849 );
xor ( n73852 , n72673 , n72952 );
nor ( n73853 , n19365 , n73665 );
and ( n73854 , n73852 , n73853 );
xor ( n73855 , n73852 , n73853 );
xor ( n73856 , n72677 , n72950 );
nor ( n73857 , n18448 , n73665 );
and ( n73858 , n73856 , n73857 );
xor ( n73859 , n73856 , n73857 );
xor ( n73860 , n72681 , n72948 );
nor ( n73861 , n17548 , n73665 );
and ( n73862 , n73860 , n73861 );
xor ( n73863 , n73860 , n73861 );
xor ( n73864 , n72685 , n72946 );
nor ( n73865 , n16669 , n73665 );
and ( n73866 , n73864 , n73865 );
xor ( n73867 , n73864 , n73865 );
xor ( n73868 , n72689 , n72944 );
nor ( n73869 , n15809 , n73665 );
and ( n73870 , n73868 , n73869 );
xor ( n73871 , n73868 , n73869 );
xor ( n73872 , n72693 , n72942 );
nor ( n73873 , n14968 , n73665 );
and ( n73874 , n73872 , n73873 );
xor ( n73875 , n73872 , n73873 );
xor ( n73876 , n72697 , n72940 );
nor ( n73877 , n14147 , n73665 );
and ( n73878 , n73876 , n73877 );
xor ( n73879 , n73876 , n73877 );
xor ( n73880 , n72701 , n72938 );
nor ( n73881 , n13349 , n73665 );
and ( n73882 , n73880 , n73881 );
xor ( n73883 , n73880 , n73881 );
xor ( n73884 , n72705 , n72936 );
nor ( n73885 , n12564 , n73665 );
and ( n73886 , n73884 , n73885 );
xor ( n73887 , n73884 , n73885 );
xor ( n73888 , n72709 , n72934 );
nor ( n73889 , n11799 , n73665 );
and ( n73890 , n73888 , n73889 );
xor ( n73891 , n73888 , n73889 );
xor ( n73892 , n72713 , n72932 );
nor ( n73893 , n11050 , n73665 );
and ( n73894 , n73892 , n73893 );
xor ( n73895 , n73892 , n73893 );
xor ( n73896 , n72717 , n72930 );
nor ( n73897 , n10321 , n73665 );
and ( n73898 , n73896 , n73897 );
xor ( n73899 , n73896 , n73897 );
xor ( n73900 , n72721 , n72928 );
nor ( n73901 , n9429 , n73665 );
and ( n73902 , n73900 , n73901 );
xor ( n73903 , n73900 , n73901 );
xor ( n73904 , n72725 , n72926 );
nor ( n73905 , n8949 , n73665 );
and ( n73906 , n73904 , n73905 );
xor ( n73907 , n73904 , n73905 );
xor ( n73908 , n72729 , n72924 );
nor ( n73909 , n9437 , n73665 );
and ( n73910 , n73908 , n73909 );
xor ( n73911 , n73908 , n73909 );
xor ( n73912 , n72733 , n72922 );
nor ( n73913 , n9446 , n73665 );
and ( n73914 , n73912 , n73913 );
xor ( n73915 , n73912 , n73913 );
xor ( n73916 , n72737 , n72920 );
nor ( n73917 , n9455 , n73665 );
and ( n73918 , n73916 , n73917 );
xor ( n73919 , n73916 , n73917 );
xor ( n73920 , n72741 , n72918 );
nor ( n73921 , n9464 , n73665 );
and ( n73922 , n73920 , n73921 );
xor ( n73923 , n73920 , n73921 );
xor ( n73924 , n72745 , n72916 );
nor ( n73925 , n9473 , n73665 );
and ( n73926 , n73924 , n73925 );
xor ( n73927 , n73924 , n73925 );
xor ( n73928 , n72749 , n72914 );
nor ( n73929 , n9482 , n73665 );
and ( n73930 , n73928 , n73929 );
xor ( n73931 , n73928 , n73929 );
xor ( n73932 , n72753 , n72912 );
nor ( n73933 , n9491 , n73665 );
and ( n73934 , n73932 , n73933 );
xor ( n73935 , n73932 , n73933 );
xor ( n73936 , n72757 , n72910 );
nor ( n73937 , n9500 , n73665 );
and ( n73938 , n73936 , n73937 );
xor ( n73939 , n73936 , n73937 );
xor ( n73940 , n72761 , n72908 );
nor ( n73941 , n9509 , n73665 );
and ( n73942 , n73940 , n73941 );
xor ( n73943 , n73940 , n73941 );
xor ( n73944 , n72765 , n72906 );
nor ( n73945 , n9518 , n73665 );
and ( n73946 , n73944 , n73945 );
xor ( n73947 , n73944 , n73945 );
xor ( n73948 , n72769 , n72904 );
nor ( n73949 , n9527 , n73665 );
and ( n73950 , n73948 , n73949 );
xor ( n73951 , n73948 , n73949 );
xor ( n73952 , n72773 , n72902 );
nor ( n73953 , n9536 , n73665 );
and ( n73954 , n73952 , n73953 );
xor ( n73955 , n73952 , n73953 );
xor ( n73956 , n72777 , n72900 );
nor ( n73957 , n9545 , n73665 );
and ( n73958 , n73956 , n73957 );
xor ( n73959 , n73956 , n73957 );
xor ( n73960 , n72781 , n72898 );
nor ( n73961 , n9554 , n73665 );
and ( n73962 , n73960 , n73961 );
xor ( n73963 , n73960 , n73961 );
xor ( n73964 , n72785 , n72896 );
nor ( n73965 , n9563 , n73665 );
and ( n73966 , n73964 , n73965 );
xor ( n73967 , n73964 , n73965 );
xor ( n73968 , n72789 , n72894 );
nor ( n73969 , n9572 , n73665 );
and ( n73970 , n73968 , n73969 );
xor ( n73971 , n73968 , n73969 );
xor ( n73972 , n72793 , n72892 );
nor ( n73973 , n9581 , n73665 );
and ( n73974 , n73972 , n73973 );
xor ( n73975 , n73972 , n73973 );
xor ( n73976 , n72797 , n72890 );
nor ( n73977 , n9590 , n73665 );
and ( n73978 , n73976 , n73977 );
xor ( n73979 , n73976 , n73977 );
xor ( n73980 , n72801 , n72888 );
nor ( n73981 , n9599 , n73665 );
and ( n73982 , n73980 , n73981 );
xor ( n73983 , n73980 , n73981 );
xor ( n73984 , n72805 , n72886 );
nor ( n73985 , n9608 , n73665 );
and ( n73986 , n73984 , n73985 );
xor ( n73987 , n73984 , n73985 );
xor ( n73988 , n72809 , n72884 );
nor ( n73989 , n9617 , n73665 );
and ( n73990 , n73988 , n73989 );
xor ( n73991 , n73988 , n73989 );
xor ( n73992 , n72813 , n72882 );
nor ( n73993 , n9626 , n73665 );
and ( n73994 , n73992 , n73993 );
xor ( n73995 , n73992 , n73993 );
xor ( n73996 , n72817 , n72880 );
nor ( n73997 , n9635 , n73665 );
and ( n73998 , n73996 , n73997 );
xor ( n73999 , n73996 , n73997 );
xor ( n74000 , n72821 , n72878 );
nor ( n74001 , n9644 , n73665 );
and ( n74002 , n74000 , n74001 );
xor ( n74003 , n74000 , n74001 );
xor ( n74004 , n72825 , n72876 );
nor ( n74005 , n9653 , n73665 );
and ( n74006 , n74004 , n74005 );
xor ( n74007 , n74004 , n74005 );
xor ( n74008 , n72829 , n72874 );
nor ( n74009 , n9662 , n73665 );
and ( n74010 , n74008 , n74009 );
xor ( n74011 , n74008 , n74009 );
xor ( n74012 , n72833 , n72872 );
nor ( n74013 , n9671 , n73665 );
and ( n74014 , n74012 , n74013 );
xor ( n74015 , n74012 , n74013 );
xor ( n74016 , n72837 , n72870 );
nor ( n74017 , n9680 , n73665 );
and ( n74018 , n74016 , n74017 );
xor ( n74019 , n74016 , n74017 );
xor ( n74020 , n72841 , n72868 );
nor ( n74021 , n9689 , n73665 );
and ( n74022 , n74020 , n74021 );
xor ( n74023 , n74020 , n74021 );
xor ( n74024 , n72845 , n72866 );
nor ( n74025 , n9698 , n73665 );
and ( n74026 , n74024 , n74025 );
xor ( n74027 , n74024 , n74025 );
xor ( n74028 , n72849 , n72864 );
nor ( n74029 , n9707 , n73665 );
and ( n74030 , n74028 , n74029 );
xor ( n74031 , n74028 , n74029 );
xor ( n74032 , n72853 , n72862 );
nor ( n74033 , n9716 , n73665 );
and ( n74034 , n74032 , n74033 );
xor ( n74035 , n74032 , n74033 );
xor ( n74036 , n72857 , n72860 );
nor ( n74037 , n9725 , n73665 );
and ( n74038 , n74036 , n74037 );
xor ( n74039 , n74036 , n74037 );
xor ( n74040 , n72858 , n72859 );
nor ( n74041 , n9734 , n73665 );
and ( n74042 , n74040 , n74041 );
xor ( n74043 , n74040 , n74041 );
nor ( n74044 , n9752 , n72483 );
nor ( n74045 , n9743 , n73665 );
and ( n74046 , n74044 , n74045 );
and ( n74047 , n74043 , n74046 );
or ( n74048 , n74042 , n74047 );
and ( n74049 , n74039 , n74048 );
or ( n74050 , n74038 , n74049 );
and ( n74051 , n74035 , n74050 );
or ( n74052 , n74034 , n74051 );
and ( n74053 , n74031 , n74052 );
or ( n74054 , n74030 , n74053 );
and ( n74055 , n74027 , n74054 );
or ( n74056 , n74026 , n74055 );
and ( n74057 , n74023 , n74056 );
or ( n74058 , n74022 , n74057 );
and ( n74059 , n74019 , n74058 );
or ( n74060 , n74018 , n74059 );
and ( n74061 , n74015 , n74060 );
or ( n74062 , n74014 , n74061 );
and ( n74063 , n74011 , n74062 );
or ( n74064 , n74010 , n74063 );
and ( n74065 , n74007 , n74064 );
or ( n74066 , n74006 , n74065 );
and ( n74067 , n74003 , n74066 );
or ( n74068 , n74002 , n74067 );
and ( n74069 , n73999 , n74068 );
or ( n74070 , n73998 , n74069 );
and ( n74071 , n73995 , n74070 );
or ( n74072 , n73994 , n74071 );
and ( n74073 , n73991 , n74072 );
or ( n74074 , n73990 , n74073 );
and ( n74075 , n73987 , n74074 );
or ( n74076 , n73986 , n74075 );
and ( n74077 , n73983 , n74076 );
or ( n74078 , n73982 , n74077 );
and ( n74079 , n73979 , n74078 );
or ( n74080 , n73978 , n74079 );
and ( n74081 , n73975 , n74080 );
or ( n74082 , n73974 , n74081 );
and ( n74083 , n73971 , n74082 );
or ( n74084 , n73970 , n74083 );
and ( n74085 , n73967 , n74084 );
or ( n74086 , n73966 , n74085 );
and ( n74087 , n73963 , n74086 );
or ( n74088 , n73962 , n74087 );
and ( n74089 , n73959 , n74088 );
or ( n74090 , n73958 , n74089 );
and ( n74091 , n73955 , n74090 );
or ( n74092 , n73954 , n74091 );
and ( n74093 , n73951 , n74092 );
or ( n74094 , n73950 , n74093 );
and ( n74095 , n73947 , n74094 );
or ( n74096 , n73946 , n74095 );
and ( n74097 , n73943 , n74096 );
or ( n74098 , n73942 , n74097 );
and ( n74099 , n73939 , n74098 );
or ( n74100 , n73938 , n74099 );
and ( n74101 , n73935 , n74100 );
or ( n74102 , n73934 , n74101 );
and ( n74103 , n73931 , n74102 );
or ( n74104 , n73930 , n74103 );
and ( n74105 , n73927 , n74104 );
or ( n74106 , n73926 , n74105 );
and ( n74107 , n73923 , n74106 );
or ( n74108 , n73922 , n74107 );
and ( n74109 , n73919 , n74108 );
or ( n74110 , n73918 , n74109 );
and ( n74111 , n73915 , n74110 );
or ( n74112 , n73914 , n74111 );
and ( n74113 , n73911 , n74112 );
or ( n74114 , n73910 , n74113 );
and ( n74115 , n73907 , n74114 );
or ( n74116 , n73906 , n74115 );
and ( n74117 , n73903 , n74116 );
or ( n74118 , n73902 , n74117 );
and ( n74119 , n73899 , n74118 );
or ( n74120 , n73898 , n74119 );
and ( n74121 , n73895 , n74120 );
or ( n74122 , n73894 , n74121 );
and ( n74123 , n73891 , n74122 );
or ( n74124 , n73890 , n74123 );
and ( n74125 , n73887 , n74124 );
or ( n74126 , n73886 , n74125 );
and ( n74127 , n73883 , n74126 );
or ( n74128 , n73882 , n74127 );
and ( n74129 , n73879 , n74128 );
or ( n74130 , n73878 , n74129 );
and ( n74131 , n73875 , n74130 );
or ( n74132 , n73874 , n74131 );
and ( n74133 , n73871 , n74132 );
or ( n74134 , n73870 , n74133 );
and ( n74135 , n73867 , n74134 );
or ( n74136 , n73866 , n74135 );
and ( n74137 , n73863 , n74136 );
or ( n74138 , n73862 , n74137 );
and ( n74139 , n73859 , n74138 );
or ( n74140 , n73858 , n74139 );
and ( n74141 , n73855 , n74140 );
or ( n74142 , n73854 , n74141 );
and ( n74143 , n73851 , n74142 );
or ( n74144 , n73850 , n74143 );
and ( n74145 , n73847 , n74144 );
or ( n74146 , n73846 , n74145 );
and ( n74147 , n73843 , n74146 );
or ( n74148 , n73842 , n74147 );
and ( n74149 , n73839 , n74148 );
or ( n74150 , n73838 , n74149 );
and ( n74151 , n73835 , n74150 );
or ( n74152 , n73834 , n74151 );
and ( n74153 , n73831 , n74152 );
or ( n74154 , n73830 , n74153 );
and ( n74155 , n73827 , n74154 );
or ( n74156 , n73826 , n74155 );
and ( n74157 , n73823 , n74156 );
or ( n74158 , n73822 , n74157 );
and ( n74159 , n73819 , n74158 );
or ( n74160 , n73818 , n74159 );
and ( n74161 , n73815 , n74160 );
or ( n74162 , n73814 , n74161 );
and ( n74163 , n73811 , n74162 );
or ( n74164 , n73810 , n74163 );
and ( n74165 , n73807 , n74164 );
or ( n74166 , n73806 , n74165 );
and ( n74167 , n73803 , n74166 );
or ( n74168 , n73802 , n74167 );
and ( n74169 , n73799 , n74168 );
or ( n74170 , n73798 , n74169 );
and ( n74171 , n73795 , n74170 );
or ( n74172 , n73794 , n74171 );
and ( n74173 , n73791 , n74172 );
or ( n74174 , n73790 , n74173 );
and ( n74175 , n73787 , n74174 );
or ( n74176 , n73786 , n74175 );
and ( n74177 , n73783 , n74176 );
or ( n74178 , n73782 , n74177 );
and ( n74179 , n73779 , n74178 );
or ( n74180 , n73778 , n74179 );
and ( n74181 , n73775 , n74180 );
or ( n74182 , n73774 , n74181 );
and ( n74183 , n73771 , n74182 );
or ( n74184 , n73770 , n74183 );
and ( n74185 , n73767 , n74184 );
or ( n74186 , n73766 , n74185 );
and ( n74187 , n73763 , n74186 );
or ( n74188 , n73762 , n74187 );
and ( n74189 , n73759 , n74188 );
or ( n74190 , n73758 , n74189 );
and ( n74191 , n73755 , n74190 );
or ( n74192 , n73754 , n74191 );
and ( n74193 , n73751 , n74192 );
or ( n74194 , n73750 , n74193 );
and ( n74195 , n73747 , n74194 );
or ( n74196 , n73746 , n74195 );
and ( n74197 , n73743 , n74196 );
or ( n74198 , n73742 , n74197 );
and ( n74199 , n73739 , n74198 );
or ( n74200 , n73738 , n74199 );
and ( n74201 , n73735 , n74200 );
or ( n74202 , n73734 , n74201 );
and ( n74203 , n73731 , n74202 );
or ( n74204 , n73730 , n74203 );
and ( n74205 , n73727 , n74204 );
or ( n74206 , n73726 , n74205 );
and ( n74207 , n73723 , n74206 );
or ( n74208 , n73722 , n74207 );
and ( n74209 , n73719 , n74208 );
or ( n74210 , n73718 , n74209 );
and ( n74211 , n73715 , n74210 );
or ( n74212 , n73714 , n74211 );
and ( n74213 , n73711 , n74212 );
or ( n74214 , n73710 , n74213 );
and ( n74215 , n73707 , n74214 );
or ( n74216 , n73706 , n74215 );
and ( n74217 , n73703 , n74216 );
or ( n74218 , n73702 , n74217 );
and ( n74219 , n73699 , n74218 );
or ( n74220 , n73698 , n74219 );
and ( n74221 , n73695 , n74220 );
or ( n74222 , n73694 , n74221 );
and ( n74223 , n73691 , n74222 );
or ( n74224 , n73690 , n74223 );
and ( n74225 , n73687 , n74224 );
or ( n74226 , n73686 , n74225 );
and ( n74227 , n73683 , n74226 );
or ( n74228 , n73682 , n74227 );
and ( n74229 , n73679 , n74228 );
or ( n74230 , n73678 , n74229 );
and ( n74231 , n73675 , n74230 );
or ( n74232 , n73674 , n74231 );
and ( n74233 , n73671 , n74232 );
or ( n74234 , n73670 , n74233 );
xor ( n74235 , n73667 , n74234 );
and ( n74236 , n33403 , n7840 );
nor ( n74237 , n7841 , n74236 );
nor ( n74238 , n8281 , n32231 );
xor ( n74239 , n74237 , n74238 );
and ( n74240 , n73049 , n73050 );
and ( n74241 , n73051 , n73054 );
or ( n74242 , n74240 , n74241 );
xor ( n74243 , n74239 , n74242 );
nor ( n74244 , n8737 , n31083 );
xor ( n74245 , n74243 , n74244 );
and ( n74246 , n73055 , n73056 );
and ( n74247 , n73057 , n73060 );
or ( n74248 , n74246 , n74247 );
xor ( n74249 , n74245 , n74248 );
nor ( n74250 , n9420 , n29948 );
xor ( n74251 , n74249 , n74250 );
and ( n74252 , n73061 , n73062 );
and ( n74253 , n73063 , n73066 );
or ( n74254 , n74252 , n74253 );
xor ( n74255 , n74251 , n74254 );
nor ( n74256 , n10312 , n28833 );
xor ( n74257 , n74255 , n74256 );
and ( n74258 , n73067 , n73068 );
and ( n74259 , n73069 , n73072 );
or ( n74260 , n74258 , n74259 );
xor ( n74261 , n74257 , n74260 );
nor ( n74262 , n11041 , n27737 );
xor ( n74263 , n74261 , n74262 );
and ( n74264 , n73073 , n73074 );
and ( n74265 , n73075 , n73078 );
or ( n74266 , n74264 , n74265 );
xor ( n74267 , n74263 , n74266 );
nor ( n74268 , n11790 , n26660 );
xor ( n74269 , n74267 , n74268 );
and ( n74270 , n73079 , n73080 );
and ( n74271 , n73081 , n73084 );
or ( n74272 , n74270 , n74271 );
xor ( n74273 , n74269 , n74272 );
nor ( n74274 , n12555 , n25600 );
xor ( n74275 , n74273 , n74274 );
and ( n74276 , n73085 , n73086 );
and ( n74277 , n73087 , n73090 );
or ( n74278 , n74276 , n74277 );
xor ( n74279 , n74275 , n74278 );
nor ( n74280 , n13340 , n24564 );
xor ( n74281 , n74279 , n74280 );
and ( n74282 , n73091 , n73092 );
and ( n74283 , n73093 , n73096 );
or ( n74284 , n74282 , n74283 );
xor ( n74285 , n74281 , n74284 );
nor ( n74286 , n14138 , n23541 );
xor ( n74287 , n74285 , n74286 );
and ( n74288 , n73097 , n73098 );
and ( n74289 , n73099 , n73102 );
or ( n74290 , n74288 , n74289 );
xor ( n74291 , n74287 , n74290 );
nor ( n74292 , n14959 , n22541 );
xor ( n74293 , n74291 , n74292 );
and ( n74294 , n73103 , n73104 );
and ( n74295 , n73105 , n73108 );
or ( n74296 , n74294 , n74295 );
xor ( n74297 , n74293 , n74296 );
nor ( n74298 , n15800 , n21562 );
xor ( n74299 , n74297 , n74298 );
and ( n74300 , n73109 , n73110 );
and ( n74301 , n73111 , n73114 );
or ( n74302 , n74300 , n74301 );
xor ( n74303 , n74299 , n74302 );
nor ( n74304 , n16660 , n20601 );
xor ( n74305 , n74303 , n74304 );
and ( n74306 , n73115 , n73116 );
and ( n74307 , n73117 , n73120 );
or ( n74308 , n74306 , n74307 );
xor ( n74309 , n74305 , n74308 );
nor ( n74310 , n17539 , n19657 );
xor ( n74311 , n74309 , n74310 );
and ( n74312 , n73121 , n73122 );
and ( n74313 , n73123 , n73126 );
or ( n74314 , n74312 , n74313 );
xor ( n74315 , n74311 , n74314 );
nor ( n74316 , n18439 , n18734 );
xor ( n74317 , n74315 , n74316 );
and ( n74318 , n73127 , n73128 );
and ( n74319 , n73129 , n73132 );
or ( n74320 , n74318 , n74319 );
xor ( n74321 , n74317 , n74320 );
nor ( n74322 , n19356 , n17828 );
xor ( n74323 , n74321 , n74322 );
and ( n74324 , n73133 , n73134 );
and ( n74325 , n73135 , n73138 );
or ( n74326 , n74324 , n74325 );
xor ( n74327 , n74323 , n74326 );
nor ( n74328 , n20294 , n16943 );
xor ( n74329 , n74327 , n74328 );
and ( n74330 , n73139 , n73140 );
and ( n74331 , n73141 , n73144 );
or ( n74332 , n74330 , n74331 );
xor ( n74333 , n74329 , n74332 );
nor ( n74334 , n21249 , n16077 );
xor ( n74335 , n74333 , n74334 );
and ( n74336 , n73145 , n73146 );
and ( n74337 , n73147 , n73150 );
or ( n74338 , n74336 , n74337 );
xor ( n74339 , n74335 , n74338 );
nor ( n74340 , n22222 , n15230 );
xor ( n74341 , n74339 , n74340 );
and ( n74342 , n73151 , n73152 );
and ( n74343 , n73153 , n73156 );
or ( n74344 , n74342 , n74343 );
xor ( n74345 , n74341 , n74344 );
nor ( n74346 , n23216 , n14403 );
xor ( n74347 , n74345 , n74346 );
and ( n74348 , n73157 , n73158 );
and ( n74349 , n73159 , n73162 );
or ( n74350 , n74348 , n74349 );
xor ( n74351 , n74347 , n74350 );
nor ( n74352 , n24233 , n13599 );
xor ( n74353 , n74351 , n74352 );
and ( n74354 , n73163 , n73164 );
and ( n74355 , n73165 , n73168 );
or ( n74356 , n74354 , n74355 );
xor ( n74357 , n74353 , n74356 );
nor ( n74358 , n25263 , n12808 );
xor ( n74359 , n74357 , n74358 );
and ( n74360 , n73169 , n73170 );
and ( n74361 , n73171 , n73174 );
or ( n74362 , n74360 , n74361 );
xor ( n74363 , n74359 , n74362 );
nor ( n74364 , n26317 , n12037 );
xor ( n74365 , n74363 , n74364 );
and ( n74366 , n73175 , n73176 );
and ( n74367 , n73177 , n73180 );
or ( n74368 , n74366 , n74367 );
xor ( n74369 , n74365 , n74368 );
nor ( n74370 , n27388 , n11282 );
xor ( n74371 , n74369 , n74370 );
and ( n74372 , n73181 , n73182 );
and ( n74373 , n73183 , n73186 );
or ( n74374 , n74372 , n74373 );
xor ( n74375 , n74371 , n74374 );
nor ( n74376 , n28478 , n10547 );
xor ( n74377 , n74375 , n74376 );
and ( n74378 , n73187 , n73188 );
and ( n74379 , n73189 , n73192 );
or ( n74380 , n74378 , n74379 );
xor ( n74381 , n74377 , n74380 );
nor ( n74382 , n29587 , n9829 );
xor ( n74383 , n74381 , n74382 );
and ( n74384 , n73193 , n73194 );
and ( n74385 , n73195 , n73198 );
or ( n74386 , n74384 , n74385 );
xor ( n74387 , n74383 , n74386 );
nor ( n74388 , n30716 , n8955 );
xor ( n74389 , n74387 , n74388 );
and ( n74390 , n73199 , n73200 );
and ( n74391 , n73201 , n73204 );
or ( n74392 , n74390 , n74391 );
xor ( n74393 , n74389 , n74392 );
nor ( n74394 , n31858 , n603 );
xor ( n74395 , n74393 , n74394 );
and ( n74396 , n73205 , n73206 );
and ( n74397 , n73207 , n73210 );
or ( n74398 , n74396 , n74397 );
xor ( n74399 , n74395 , n74398 );
nor ( n74400 , n33024 , n652 );
xor ( n74401 , n74399 , n74400 );
and ( n74402 , n73211 , n73212 );
and ( n74403 , n73213 , n73216 );
or ( n74404 , n74402 , n74403 );
xor ( n74405 , n74401 , n74404 );
nor ( n74406 , n34215 , n624 );
xor ( n74407 , n74405 , n74406 );
and ( n74408 , n73217 , n73218 );
and ( n74409 , n73219 , n73222 );
or ( n74410 , n74408 , n74409 );
xor ( n74411 , n74407 , n74410 );
nor ( n74412 , n35410 , n648 );
xor ( n74413 , n74411 , n74412 );
and ( n74414 , n73223 , n73224 );
and ( n74415 , n73225 , n73228 );
or ( n74416 , n74414 , n74415 );
xor ( n74417 , n74413 , n74416 );
nor ( n74418 , n36611 , n686 );
xor ( n74419 , n74417 , n74418 );
and ( n74420 , n73229 , n73230 );
and ( n74421 , n73231 , n73234 );
or ( n74422 , n74420 , n74421 );
xor ( n74423 , n74419 , n74422 );
nor ( n74424 , n37816 , n735 );
xor ( n74425 , n74423 , n74424 );
and ( n74426 , n73235 , n73236 );
and ( n74427 , n73237 , n73240 );
or ( n74428 , n74426 , n74427 );
xor ( n74429 , n74425 , n74428 );
nor ( n74430 , n39018 , n798 );
xor ( n74431 , n74429 , n74430 );
and ( n74432 , n73241 , n73242 );
and ( n74433 , n73243 , n73246 );
or ( n74434 , n74432 , n74433 );
xor ( n74435 , n74431 , n74434 );
nor ( n74436 , n40223 , n870 );
xor ( n74437 , n74435 , n74436 );
and ( n74438 , n73247 , n73248 );
and ( n74439 , n73249 , n73252 );
or ( n74440 , n74438 , n74439 );
xor ( n74441 , n74437 , n74440 );
nor ( n74442 , n41428 , n960 );
xor ( n74443 , n74441 , n74442 );
and ( n74444 , n73253 , n73254 );
and ( n74445 , n73255 , n73258 );
or ( n74446 , n74444 , n74445 );
xor ( n74447 , n74443 , n74446 );
nor ( n74448 , n42632 , n1064 );
xor ( n74449 , n74447 , n74448 );
and ( n74450 , n73259 , n73260 );
and ( n74451 , n73261 , n73264 );
or ( n74452 , n74450 , n74451 );
xor ( n74453 , n74449 , n74452 );
nor ( n74454 , n43834 , n1178 );
xor ( n74455 , n74453 , n74454 );
and ( n74456 , n73265 , n73266 );
and ( n74457 , n73267 , n73270 );
or ( n74458 , n74456 , n74457 );
xor ( n74459 , n74455 , n74458 );
nor ( n74460 , n45038 , n1305 );
xor ( n74461 , n74459 , n74460 );
and ( n74462 , n73271 , n73272 );
and ( n74463 , n73273 , n73276 );
or ( n74464 , n74462 , n74463 );
xor ( n74465 , n74461 , n74464 );
nor ( n74466 , n46239 , n1447 );
xor ( n74467 , n74465 , n74466 );
and ( n74468 , n73277 , n73278 );
and ( n74469 , n73279 , n73282 );
or ( n74470 , n74468 , n74469 );
xor ( n74471 , n74467 , n74470 );
nor ( n74472 , n47440 , n1600 );
xor ( n74473 , n74471 , n74472 );
and ( n74474 , n73283 , n73284 );
and ( n74475 , n73285 , n73288 );
or ( n74476 , n74474 , n74475 );
xor ( n74477 , n74473 , n74476 );
nor ( n74478 , n48641 , n1768 );
xor ( n74479 , n74477 , n74478 );
and ( n74480 , n73289 , n73290 );
and ( n74481 , n73291 , n73294 );
or ( n74482 , n74480 , n74481 );
xor ( n74483 , n74479 , n74482 );
nor ( n74484 , n49841 , n1947 );
xor ( n74485 , n74483 , n74484 );
and ( n74486 , n73295 , n73296 );
and ( n74487 , n73297 , n73300 );
or ( n74488 , n74486 , n74487 );
xor ( n74489 , n74485 , n74488 );
nor ( n74490 , n51040 , n2139 );
xor ( n74491 , n74489 , n74490 );
and ( n74492 , n73301 , n73302 );
and ( n74493 , n73303 , n73306 );
or ( n74494 , n74492 , n74493 );
xor ( n74495 , n74491 , n74494 );
nor ( n74496 , n52238 , n2345 );
xor ( n74497 , n74495 , n74496 );
and ( n74498 , n73307 , n73308 );
and ( n74499 , n73309 , n73312 );
or ( n74500 , n74498 , n74499 );
xor ( n74501 , n74497 , n74500 );
nor ( n74502 , n53432 , n2568 );
xor ( n74503 , n74501 , n74502 );
and ( n74504 , n73313 , n73314 );
and ( n74505 , n73315 , n73318 );
or ( n74506 , n74504 , n74505 );
xor ( n74507 , n74503 , n74506 );
nor ( n74508 , n54629 , n2799 );
xor ( n74509 , n74507 , n74508 );
and ( n74510 , n73319 , n73320 );
and ( n74511 , n73321 , n73324 );
or ( n74512 , n74510 , n74511 );
xor ( n74513 , n74509 , n74512 );
nor ( n74514 , n55826 , n3045 );
xor ( n74515 , n74513 , n74514 );
and ( n74516 , n73325 , n73326 );
and ( n74517 , n73327 , n73330 );
or ( n74518 , n74516 , n74517 );
xor ( n74519 , n74515 , n74518 );
nor ( n74520 , n57022 , n3302 );
xor ( n74521 , n74519 , n74520 );
and ( n74522 , n73331 , n73332 );
and ( n74523 , n73333 , n73336 );
or ( n74524 , n74522 , n74523 );
xor ( n74525 , n74521 , n74524 );
nor ( n74526 , n58217 , n3572 );
xor ( n74527 , n74525 , n74526 );
and ( n74528 , n73337 , n73338 );
and ( n74529 , n73339 , n73342 );
or ( n74530 , n74528 , n74529 );
xor ( n74531 , n74527 , n74530 );
nor ( n74532 , n59412 , n3855 );
xor ( n74533 , n74531 , n74532 );
and ( n74534 , n73343 , n73344 );
and ( n74535 , n73345 , n73348 );
or ( n74536 , n74534 , n74535 );
xor ( n74537 , n74533 , n74536 );
nor ( n74538 , n60600 , n4153 );
xor ( n74539 , n74537 , n74538 );
and ( n74540 , n73349 , n73350 );
and ( n74541 , n73351 , n73354 );
or ( n74542 , n74540 , n74541 );
xor ( n74543 , n74539 , n74542 );
nor ( n74544 , n61791 , n4460 );
xor ( n74545 , n74543 , n74544 );
and ( n74546 , n73355 , n73356 );
and ( n74547 , n73357 , n73360 );
or ( n74548 , n74546 , n74547 );
xor ( n74549 , n74545 , n74548 );
nor ( n74550 , n62982 , n4788 );
xor ( n74551 , n74549 , n74550 );
and ( n74552 , n73361 , n73362 );
and ( n74553 , n73363 , n73366 );
or ( n74554 , n74552 , n74553 );
xor ( n74555 , n74551 , n74554 );
nor ( n74556 , n64172 , n5128 );
xor ( n74557 , n74555 , n74556 );
and ( n74558 , n73367 , n73368 );
and ( n74559 , n73369 , n73372 );
or ( n74560 , n74558 , n74559 );
xor ( n74561 , n74557 , n74560 );
nor ( n74562 , n65360 , n5479 );
xor ( n74563 , n74561 , n74562 );
and ( n74564 , n73373 , n73374 );
and ( n74565 , n73375 , n73378 );
or ( n74566 , n74564 , n74565 );
xor ( n74567 , n74563 , n74566 );
nor ( n74568 , n66550 , n5840 );
xor ( n74569 , n74567 , n74568 );
and ( n74570 , n73379 , n73380 );
and ( n74571 , n73381 , n73384 );
or ( n74572 , n74570 , n74571 );
xor ( n74573 , n74569 , n74572 );
nor ( n74574 , n67736 , n6214 );
xor ( n74575 , n74573 , n74574 );
and ( n74576 , n73385 , n73386 );
and ( n74577 , n73387 , n73390 );
or ( n74578 , n74576 , n74577 );
xor ( n74579 , n74575 , n74578 );
nor ( n74580 , n68924 , n6598 );
xor ( n74581 , n74579 , n74580 );
and ( n74582 , n73391 , n73392 );
and ( n74583 , n73393 , n73396 );
or ( n74584 , n74582 , n74583 );
xor ( n74585 , n74581 , n74584 );
nor ( n74586 , n70110 , n6999 );
xor ( n74587 , n74585 , n74586 );
and ( n74588 , n73397 , n73398 );
and ( n74589 , n73399 , n73402 );
or ( n74590 , n74588 , n74589 );
xor ( n74591 , n74587 , n74590 );
nor ( n74592 , n71292 , n7415 );
xor ( n74593 , n74591 , n74592 );
and ( n74594 , n73403 , n73404 );
and ( n74595 , n73405 , n73408 );
or ( n74596 , n74594 , n74595 );
xor ( n74597 , n74593 , n74596 );
nor ( n74598 , n72472 , n7843 );
xor ( n74599 , n74597 , n74598 );
and ( n74600 , n73409 , n73410 );
and ( n74601 , n73411 , n73414 );
or ( n74602 , n74600 , n74601 );
xor ( n74603 , n74599 , n74602 );
nor ( n74604 , n73654 , n8283 );
xor ( n74605 , n74603 , n74604 );
and ( n74606 , n73415 , n73416 );
and ( n74607 , n73417 , n73420 );
or ( n74608 , n74606 , n74607 );
xor ( n74609 , n74605 , n74608 );
and ( n74610 , n73433 , n73437 );
and ( n74611 , n73437 , n73640 );
and ( n74612 , n73433 , n73640 );
or ( n74613 , n74610 , n74611 , n74612 );
and ( n74614 , n33774 , n7662 );
not ( n74615 , n7662 );
nor ( n74616 , n74614 , n74615 );
xor ( n74617 , n74613 , n74616 );
and ( n74618 , n73443 , n73444 );
and ( n74619 , n73444 , n73512 );
and ( n74620 , n73443 , n73512 );
or ( n74621 , n74618 , n74619 , n74620 );
and ( n74622 , n73439 , n73513 );
and ( n74623 , n73513 , n73639 );
and ( n74624 , n73439 , n73639 );
or ( n74625 , n74622 , n74623 , n74624 );
xor ( n74626 , n74621 , n74625 );
and ( n74627 , n73526 , n73638 );
and ( n74628 , n73449 , n73453 );
and ( n74629 , n73453 , n73511 );
and ( n74630 , n73449 , n73511 );
or ( n74631 , n74628 , n74629 , n74630 );
and ( n74632 , n73530 , n73637 );
xor ( n74633 , n74631 , n74632 );
and ( n74634 , n73480 , n73484 );
and ( n74635 , n73484 , n73490 );
and ( n74636 , n73480 , n73490 );
or ( n74637 , n74634 , n74635 , n74636 );
and ( n74638 , n73458 , n73462 );
and ( n74639 , n73462 , n73510 );
and ( n74640 , n73458 , n73510 );
or ( n74641 , n74638 , n74639 , n74640 );
xor ( n74642 , n74637 , n74641 );
and ( n74643 , n73467 , n73471 );
and ( n74644 , n73471 , n73509 );
and ( n74645 , n73467 , n73509 );
or ( n74646 , n74643 , n74644 , n74645 );
and ( n74647 , n73538 , n73563 );
and ( n74648 , n73563 , n73601 );
and ( n74649 , n73538 , n73601 );
or ( n74650 , n74647 , n74648 , n74649 );
xor ( n74651 , n74646 , n74650 );
and ( n74652 , n73476 , n73491 );
and ( n74653 , n73491 , n73508 );
and ( n74654 , n73476 , n73508 );
or ( n74655 , n74652 , n74653 , n74654 );
and ( n74656 , n73542 , n73546 );
and ( n74657 , n73546 , n73562 );
and ( n74658 , n73542 , n73562 );
or ( n74659 , n74656 , n74657 , n74658 );
xor ( n74660 , n74655 , n74659 );
and ( n74661 , n73496 , n73501 );
and ( n74662 , n73501 , n73507 );
and ( n74663 , n73496 , n73507 );
or ( n74664 , n74661 , n74662 , n74663 );
and ( n74665 , n73486 , n73487 );
and ( n74666 , n73487 , n73489 );
and ( n74667 , n73486 , n73489 );
or ( n74668 , n74665 , n74666 , n74667 );
and ( n74669 , n73497 , n73498 );
and ( n74670 , n73498 , n73500 );
and ( n74671 , n73497 , n73500 );
or ( n74672 , n74669 , n74670 , n74671 );
xor ( n74673 , n74668 , n74672 );
and ( n74674 , n30695 , n9348 );
and ( n74675 , n31836 , n8669 );
xor ( n74676 , n74674 , n74675 );
and ( n74677 , n32649 , n8243 );
xor ( n74678 , n74676 , n74677 );
xor ( n74679 , n74673 , n74678 );
xor ( n74680 , n74664 , n74679 );
and ( n74681 , n73503 , n73504 );
and ( n74682 , n73504 , n73506 );
and ( n74683 , n73503 , n73506 );
or ( n74684 , n74681 , n74682 , n74683 );
and ( n74685 , n27361 , n11718 );
and ( n74686 , n28456 , n10977 );
xor ( n74687 , n74685 , n74686 );
and ( n74688 , n29559 , n10239 );
xor ( n74689 , n74687 , n74688 );
xor ( n74690 , n74684 , n74689 );
and ( n74691 , n24214 , n14044 );
and ( n74692 , n25243 , n13256 );
xor ( n74693 , n74691 , n74692 );
and ( n74694 , n26296 , n12531 );
xor ( n74695 , n74693 , n74694 );
xor ( n74696 , n74690 , n74695 );
xor ( n74697 , n74680 , n74696 );
xor ( n74698 , n74660 , n74697 );
xor ( n74699 , n74651 , n74698 );
xor ( n74700 , n74642 , n74699 );
xor ( n74701 , n74633 , n74700 );
xor ( n74702 , n74627 , n74701 );
and ( n74703 , n73521 , n73522 );
and ( n74704 , n73522 , n73524 );
and ( n74705 , n73521 , n73524 );
or ( n74706 , n74703 , n74704 , n74705 );
not ( n74707 , n7808 );
and ( n74708 , n34193 , n7808 );
nor ( n74709 , n74707 , n74708 );
and ( n74710 , n8079 , n32999 );
xor ( n74711 , n74709 , n74710 );
xor ( n74712 , n74706 , n74711 );
and ( n74713 , n73534 , n73602 );
and ( n74714 , n73602 , n73636 );
and ( n74715 , n73534 , n73636 );
or ( n74716 , n74713 , n74714 , n74715 );
and ( n74717 , n73607 , n73608 );
and ( n74718 , n73608 , n73635 );
and ( n74719 , n73607 , n73635 );
or ( n74720 , n74717 , n74718 , n74719 );
and ( n74721 , n73568 , n73584 );
and ( n74722 , n73584 , n73600 );
and ( n74723 , n73568 , n73600 );
or ( n74724 , n74721 , n74722 , n74723 );
and ( n74725 , n73551 , n73555 );
and ( n74726 , n73555 , n73561 );
and ( n74727 , n73551 , n73561 );
or ( n74728 , n74725 , n74726 , n74727 );
and ( n74729 , n73572 , n73577 );
and ( n74730 , n73577 , n73583 );
and ( n74731 , n73572 , n73583 );
or ( n74732 , n74729 , n74730 , n74731 );
xor ( n74733 , n74728 , n74732 );
and ( n74734 , n73557 , n73558 );
and ( n74735 , n73558 , n73560 );
and ( n74736 , n73557 , n73560 );
or ( n74737 , n74734 , n74735 , n74736 );
and ( n74738 , n73573 , n73574 );
and ( n74739 , n73574 , n73576 );
and ( n74740 , n73573 , n73576 );
or ( n74741 , n74738 , n74739 , n74740 );
xor ( n74742 , n74737 , n74741 );
and ( n74743 , n21216 , n16550 );
and ( n74744 , n22186 , n15691 );
xor ( n74745 , n74743 , n74744 );
and ( n74746 , n22892 , n14838 );
xor ( n74747 , n74745 , n74746 );
xor ( n74748 , n74742 , n74747 );
xor ( n74749 , n74733 , n74748 );
xor ( n74750 , n74724 , n74749 );
and ( n74751 , n73589 , n73593 );
and ( n74752 , n73593 , n73599 );
and ( n74753 , n73589 , n73599 );
or ( n74754 , n74751 , n74752 , n74753 );
and ( n74755 , n73579 , n73580 );
and ( n74756 , n73580 , n73582 );
and ( n74757 , n73579 , n73582 );
or ( n74758 , n74755 , n74756 , n74757 );
and ( n74759 , n15758 , n22065 );
and ( n74760 , n16637 , n20976 );
xor ( n74761 , n74759 , n74760 );
and ( n74762 , n17512 , n20156 );
xor ( n74763 , n74761 , n74762 );
xor ( n74764 , n74758 , n74763 );
and ( n74765 , n20233 , n17422 );
buf ( n74766 , n74765 );
xor ( n74767 , n74764 , n74766 );
xor ( n74768 , n74754 , n74767 );
and ( n74769 , n73595 , n73596 );
and ( n74770 , n73596 , n73598 );
and ( n74771 , n73595 , n73598 );
or ( n74772 , n74769 , n74770 , n74771 );
and ( n74773 , n73623 , n73624 );
and ( n74774 , n73624 , n73626 );
and ( n74775 , n73623 , n73626 );
or ( n74776 , n74773 , n74774 , n74775 );
xor ( n74777 , n74772 , n74776 );
and ( n74778 , n13322 , n25163 );
and ( n74779 , n14118 , n24137 );
xor ( n74780 , n74778 , n74779 );
and ( n74781 , n14938 , n23075 );
xor ( n74782 , n74780 , n74781 );
xor ( n74783 , n74777 , n74782 );
xor ( n74784 , n74768 , n74783 );
xor ( n74785 , n74750 , n74784 );
xor ( n74786 , n74720 , n74785 );
and ( n74787 , n73613 , n73617 );
and ( n74788 , n73617 , n73634 );
and ( n74789 , n73613 , n73634 );
or ( n74790 , n74787 , n74788 , n74789 );
and ( n74791 , n73622 , n73627 );
and ( n74792 , n73627 , n73633 );
and ( n74793 , n73622 , n73633 );
or ( n74794 , n74791 , n74792 , n74793 );
and ( n74795 , n73518 , n73525 );
xor ( n74796 , n74794 , n74795 );
and ( n74797 , n73629 , n73630 );
and ( n74798 , n73630 , n73632 );
and ( n74799 , n73629 , n73632 );
or ( n74800 , n74797 , n74798 , n74799 );
and ( n74801 , n8718 , n31761 );
and ( n74802 , n9400 , n30629 );
xor ( n74803 , n74801 , n74802 );
and ( n74804 , n10291 , n29508 );
xor ( n74805 , n74803 , n74804 );
xor ( n74806 , n74800 , n74805 );
and ( n74807 , n11015 , n28406 );
and ( n74808 , n11769 , n27296 );
xor ( n74809 , n74807 , n74808 );
and ( n74810 , n12320 , n26216 );
xor ( n74811 , n74809 , n74810 );
xor ( n74812 , n74806 , n74811 );
xor ( n74813 , n74796 , n74812 );
xor ( n74814 , n74790 , n74813 );
xor ( n74815 , n74786 , n74814 );
xor ( n74816 , n74716 , n74815 );
xor ( n74817 , n74712 , n74816 );
xor ( n74818 , n74702 , n74817 );
xor ( n74819 , n74626 , n74818 );
xor ( n74820 , n74617 , n74819 );
and ( n74821 , n73425 , n73428 );
and ( n74822 , n73428 , n73641 );
and ( n74823 , n73425 , n73641 );
or ( n74824 , n74821 , n74822 , n74823 );
xor ( n74825 , n74820 , n74824 );
and ( n74826 , n73642 , n73646 );
and ( n74827 , n73647 , n73650 );
or ( n74828 , n74826 , n74827 );
xor ( n74829 , n74825 , n74828 );
buf ( n74830 , n74829 );
buf ( n74831 , n74830 );
not ( n74832 , n74831 );
nor ( n74833 , n74832 , n8739 );
xor ( n74834 , n74609 , n74833 );
and ( n74835 , n73421 , n73655 );
and ( n74836 , n73656 , n73659 );
or ( n74837 , n74835 , n74836 );
xor ( n74838 , n74834 , n74837 );
buf ( n74839 , n74838 );
buf ( n74840 , n74839 );
not ( n74841 , n74840 );
buf ( n74842 , n596 );
not ( n74843 , n74842 );
nor ( n74844 , n74841 , n74843 );
xor ( n74845 , n74235 , n74844 );
xor ( n74846 , n73671 , n74232 );
nor ( n74847 , n73663 , n74843 );
and ( n74848 , n74846 , n74847 );
xor ( n74849 , n74846 , n74847 );
xor ( n74850 , n73675 , n74230 );
nor ( n74851 , n72481 , n74843 );
and ( n74852 , n74850 , n74851 );
xor ( n74853 , n74850 , n74851 );
xor ( n74854 , n73679 , n74228 );
nor ( n74855 , n71301 , n74843 );
and ( n74856 , n74854 , n74855 );
xor ( n74857 , n74854 , n74855 );
xor ( n74858 , n73683 , n74226 );
nor ( n74859 , n70119 , n74843 );
and ( n74860 , n74858 , n74859 );
xor ( n74861 , n74858 , n74859 );
xor ( n74862 , n73687 , n74224 );
nor ( n74863 , n68933 , n74843 );
and ( n74864 , n74862 , n74863 );
xor ( n74865 , n74862 , n74863 );
xor ( n74866 , n73691 , n74222 );
nor ( n74867 , n67745 , n74843 );
and ( n74868 , n74866 , n74867 );
xor ( n74869 , n74866 , n74867 );
xor ( n74870 , n73695 , n74220 );
nor ( n74871 , n66559 , n74843 );
and ( n74872 , n74870 , n74871 );
xor ( n74873 , n74870 , n74871 );
xor ( n74874 , n73699 , n74218 );
nor ( n74875 , n65369 , n74843 );
and ( n74876 , n74874 , n74875 );
xor ( n74877 , n74874 , n74875 );
xor ( n74878 , n73703 , n74216 );
nor ( n74879 , n64181 , n74843 );
and ( n74880 , n74878 , n74879 );
xor ( n74881 , n74878 , n74879 );
xor ( n74882 , n73707 , n74214 );
nor ( n74883 , n62991 , n74843 );
and ( n74884 , n74882 , n74883 );
xor ( n74885 , n74882 , n74883 );
xor ( n74886 , n73711 , n74212 );
nor ( n74887 , n61800 , n74843 );
and ( n74888 , n74886 , n74887 );
xor ( n74889 , n74886 , n74887 );
xor ( n74890 , n73715 , n74210 );
nor ( n74891 , n60609 , n74843 );
and ( n74892 , n74890 , n74891 );
xor ( n74893 , n74890 , n74891 );
xor ( n74894 , n73719 , n74208 );
nor ( n74895 , n59421 , n74843 );
and ( n74896 , n74894 , n74895 );
xor ( n74897 , n74894 , n74895 );
xor ( n74898 , n73723 , n74206 );
nor ( n74899 , n58226 , n74843 );
and ( n74900 , n74898 , n74899 );
xor ( n74901 , n74898 , n74899 );
xor ( n74902 , n73727 , n74204 );
nor ( n74903 , n57031 , n74843 );
and ( n74904 , n74902 , n74903 );
xor ( n74905 , n74902 , n74903 );
xor ( n74906 , n73731 , n74202 );
nor ( n74907 , n55835 , n74843 );
and ( n74908 , n74906 , n74907 );
xor ( n74909 , n74906 , n74907 );
xor ( n74910 , n73735 , n74200 );
nor ( n74911 , n54638 , n74843 );
and ( n74912 , n74910 , n74911 );
xor ( n74913 , n74910 , n74911 );
xor ( n74914 , n73739 , n74198 );
nor ( n74915 , n53441 , n74843 );
and ( n74916 , n74914 , n74915 );
xor ( n74917 , n74914 , n74915 );
xor ( n74918 , n73743 , n74196 );
nor ( n74919 , n52247 , n74843 );
and ( n74920 , n74918 , n74919 );
xor ( n74921 , n74918 , n74919 );
xor ( n74922 , n73747 , n74194 );
nor ( n74923 , n51049 , n74843 );
and ( n74924 , n74922 , n74923 );
xor ( n74925 , n74922 , n74923 );
xor ( n74926 , n73751 , n74192 );
nor ( n74927 , n49850 , n74843 );
and ( n74928 , n74926 , n74927 );
xor ( n74929 , n74926 , n74927 );
xor ( n74930 , n73755 , n74190 );
nor ( n74931 , n48650 , n74843 );
and ( n74932 , n74930 , n74931 );
xor ( n74933 , n74930 , n74931 );
xor ( n74934 , n73759 , n74188 );
nor ( n74935 , n47449 , n74843 );
and ( n74936 , n74934 , n74935 );
xor ( n74937 , n74934 , n74935 );
xor ( n74938 , n73763 , n74186 );
nor ( n74939 , n46248 , n74843 );
and ( n74940 , n74938 , n74939 );
xor ( n74941 , n74938 , n74939 );
xor ( n74942 , n73767 , n74184 );
nor ( n74943 , n45047 , n74843 );
and ( n74944 , n74942 , n74943 );
xor ( n74945 , n74942 , n74943 );
xor ( n74946 , n73771 , n74182 );
nor ( n74947 , n43843 , n74843 );
and ( n74948 , n74946 , n74947 );
xor ( n74949 , n74946 , n74947 );
xor ( n74950 , n73775 , n74180 );
nor ( n74951 , n42641 , n74843 );
and ( n74952 , n74950 , n74951 );
xor ( n74953 , n74950 , n74951 );
xor ( n74954 , n73779 , n74178 );
nor ( n74955 , n41437 , n74843 );
and ( n74956 , n74954 , n74955 );
xor ( n74957 , n74954 , n74955 );
xor ( n74958 , n73783 , n74176 );
nor ( n74959 , n40232 , n74843 );
and ( n74960 , n74958 , n74959 );
xor ( n74961 , n74958 , n74959 );
xor ( n74962 , n73787 , n74174 );
nor ( n74963 , n39027 , n74843 );
and ( n74964 , n74962 , n74963 );
xor ( n74965 , n74962 , n74963 );
xor ( n74966 , n73791 , n74172 );
nor ( n74967 , n37825 , n74843 );
and ( n74968 , n74966 , n74967 );
xor ( n74969 , n74966 , n74967 );
xor ( n74970 , n73795 , n74170 );
nor ( n74971 , n36620 , n74843 );
and ( n74972 , n74970 , n74971 );
xor ( n74973 , n74970 , n74971 );
xor ( n74974 , n73799 , n74168 );
nor ( n74975 , n35419 , n74843 );
and ( n74976 , n74974 , n74975 );
xor ( n74977 , n74974 , n74975 );
xor ( n74978 , n73803 , n74166 );
nor ( n74979 , n34224 , n74843 );
and ( n74980 , n74978 , n74979 );
xor ( n74981 , n74978 , n74979 );
xor ( n74982 , n73807 , n74164 );
nor ( n74983 , n33033 , n74843 );
and ( n74984 , n74982 , n74983 );
xor ( n74985 , n74982 , n74983 );
xor ( n74986 , n73811 , n74162 );
nor ( n74987 , n31867 , n74843 );
and ( n74988 , n74986 , n74987 );
xor ( n74989 , n74986 , n74987 );
xor ( n74990 , n73815 , n74160 );
nor ( n74991 , n30725 , n74843 );
and ( n74992 , n74990 , n74991 );
xor ( n74993 , n74990 , n74991 );
xor ( n74994 , n73819 , n74158 );
nor ( n74995 , n29596 , n74843 );
and ( n74996 , n74994 , n74995 );
xor ( n74997 , n74994 , n74995 );
xor ( n74998 , n73823 , n74156 );
nor ( n74999 , n28487 , n74843 );
and ( n75000 , n74998 , n74999 );
xor ( n75001 , n74998 , n74999 );
xor ( n75002 , n73827 , n74154 );
nor ( n75003 , n27397 , n74843 );
and ( n75004 , n75002 , n75003 );
xor ( n75005 , n75002 , n75003 );
xor ( n75006 , n73831 , n74152 );
nor ( n75007 , n26326 , n74843 );
and ( n75008 , n75006 , n75007 );
xor ( n75009 , n75006 , n75007 );
xor ( n75010 , n73835 , n74150 );
nor ( n75011 , n25272 , n74843 );
and ( n75012 , n75010 , n75011 );
xor ( n75013 , n75010 , n75011 );
xor ( n75014 , n73839 , n74148 );
nor ( n75015 , n24242 , n74843 );
and ( n75016 , n75014 , n75015 );
xor ( n75017 , n75014 , n75015 );
xor ( n75018 , n73843 , n74146 );
nor ( n75019 , n23225 , n74843 );
and ( n75020 , n75018 , n75019 );
xor ( n75021 , n75018 , n75019 );
xor ( n75022 , n73847 , n74144 );
nor ( n75023 , n22231 , n74843 );
and ( n75024 , n75022 , n75023 );
xor ( n75025 , n75022 , n75023 );
xor ( n75026 , n73851 , n74142 );
nor ( n75027 , n21258 , n74843 );
and ( n75028 , n75026 , n75027 );
xor ( n75029 , n75026 , n75027 );
xor ( n75030 , n73855 , n74140 );
nor ( n75031 , n20303 , n74843 );
and ( n75032 , n75030 , n75031 );
xor ( n75033 , n75030 , n75031 );
xor ( n75034 , n73859 , n74138 );
nor ( n75035 , n19365 , n74843 );
and ( n75036 , n75034 , n75035 );
xor ( n75037 , n75034 , n75035 );
xor ( n75038 , n73863 , n74136 );
nor ( n75039 , n18448 , n74843 );
and ( n75040 , n75038 , n75039 );
xor ( n75041 , n75038 , n75039 );
xor ( n75042 , n73867 , n74134 );
nor ( n75043 , n17548 , n74843 );
and ( n75044 , n75042 , n75043 );
xor ( n75045 , n75042 , n75043 );
xor ( n75046 , n73871 , n74132 );
nor ( n75047 , n16669 , n74843 );
and ( n75048 , n75046 , n75047 );
xor ( n75049 , n75046 , n75047 );
xor ( n75050 , n73875 , n74130 );
nor ( n75051 , n15809 , n74843 );
and ( n75052 , n75050 , n75051 );
xor ( n75053 , n75050 , n75051 );
xor ( n75054 , n73879 , n74128 );
nor ( n75055 , n14968 , n74843 );
and ( n75056 , n75054 , n75055 );
xor ( n75057 , n75054 , n75055 );
xor ( n75058 , n73883 , n74126 );
nor ( n75059 , n14147 , n74843 );
and ( n75060 , n75058 , n75059 );
xor ( n75061 , n75058 , n75059 );
xor ( n75062 , n73887 , n74124 );
nor ( n75063 , n13349 , n74843 );
and ( n75064 , n75062 , n75063 );
xor ( n75065 , n75062 , n75063 );
xor ( n75066 , n73891 , n74122 );
nor ( n75067 , n12564 , n74843 );
and ( n75068 , n75066 , n75067 );
xor ( n75069 , n75066 , n75067 );
xor ( n75070 , n73895 , n74120 );
nor ( n75071 , n11799 , n74843 );
and ( n75072 , n75070 , n75071 );
xor ( n75073 , n75070 , n75071 );
xor ( n75074 , n73899 , n74118 );
nor ( n75075 , n11050 , n74843 );
and ( n75076 , n75074 , n75075 );
xor ( n75077 , n75074 , n75075 );
xor ( n75078 , n73903 , n74116 );
nor ( n75079 , n10321 , n74843 );
and ( n75080 , n75078 , n75079 );
xor ( n75081 , n75078 , n75079 );
xor ( n75082 , n73907 , n74114 );
nor ( n75083 , n9429 , n74843 );
and ( n75084 , n75082 , n75083 );
xor ( n75085 , n75082 , n75083 );
xor ( n75086 , n73911 , n74112 );
nor ( n75087 , n8949 , n74843 );
and ( n75088 , n75086 , n75087 );
xor ( n75089 , n75086 , n75087 );
xor ( n75090 , n73915 , n74110 );
nor ( n75091 , n9437 , n74843 );
and ( n75092 , n75090 , n75091 );
xor ( n75093 , n75090 , n75091 );
xor ( n75094 , n73919 , n74108 );
nor ( n75095 , n9446 , n74843 );
and ( n75096 , n75094 , n75095 );
xor ( n75097 , n75094 , n75095 );
xor ( n75098 , n73923 , n74106 );
nor ( n75099 , n9455 , n74843 );
and ( n75100 , n75098 , n75099 );
xor ( n75101 , n75098 , n75099 );
xor ( n75102 , n73927 , n74104 );
nor ( n75103 , n9464 , n74843 );
and ( n75104 , n75102 , n75103 );
xor ( n75105 , n75102 , n75103 );
xor ( n75106 , n73931 , n74102 );
nor ( n75107 , n9473 , n74843 );
and ( n75108 , n75106 , n75107 );
xor ( n75109 , n75106 , n75107 );
xor ( n75110 , n73935 , n74100 );
nor ( n75111 , n9482 , n74843 );
and ( n75112 , n75110 , n75111 );
xor ( n75113 , n75110 , n75111 );
xor ( n75114 , n73939 , n74098 );
nor ( n75115 , n9491 , n74843 );
and ( n75116 , n75114 , n75115 );
xor ( n75117 , n75114 , n75115 );
xor ( n75118 , n73943 , n74096 );
nor ( n75119 , n9500 , n74843 );
and ( n75120 , n75118 , n75119 );
xor ( n75121 , n75118 , n75119 );
xor ( n75122 , n73947 , n74094 );
nor ( n75123 , n9509 , n74843 );
and ( n75124 , n75122 , n75123 );
xor ( n75125 , n75122 , n75123 );
xor ( n75126 , n73951 , n74092 );
nor ( n75127 , n9518 , n74843 );
and ( n75128 , n75126 , n75127 );
xor ( n75129 , n75126 , n75127 );
xor ( n75130 , n73955 , n74090 );
nor ( n75131 , n9527 , n74843 );
and ( n75132 , n75130 , n75131 );
xor ( n75133 , n75130 , n75131 );
xor ( n75134 , n73959 , n74088 );
nor ( n75135 , n9536 , n74843 );
and ( n75136 , n75134 , n75135 );
xor ( n75137 , n75134 , n75135 );
xor ( n75138 , n73963 , n74086 );
nor ( n75139 , n9545 , n74843 );
and ( n75140 , n75138 , n75139 );
xor ( n75141 , n75138 , n75139 );
xor ( n75142 , n73967 , n74084 );
nor ( n75143 , n9554 , n74843 );
and ( n75144 , n75142 , n75143 );
xor ( n75145 , n75142 , n75143 );
xor ( n75146 , n73971 , n74082 );
nor ( n75147 , n9563 , n74843 );
and ( n75148 , n75146 , n75147 );
xor ( n75149 , n75146 , n75147 );
xor ( n75150 , n73975 , n74080 );
nor ( n75151 , n9572 , n74843 );
and ( n75152 , n75150 , n75151 );
xor ( n75153 , n75150 , n75151 );
xor ( n75154 , n73979 , n74078 );
nor ( n75155 , n9581 , n74843 );
and ( n75156 , n75154 , n75155 );
xor ( n75157 , n75154 , n75155 );
xor ( n75158 , n73983 , n74076 );
nor ( n75159 , n9590 , n74843 );
and ( n75160 , n75158 , n75159 );
xor ( n75161 , n75158 , n75159 );
xor ( n75162 , n73987 , n74074 );
nor ( n75163 , n9599 , n74843 );
and ( n75164 , n75162 , n75163 );
xor ( n75165 , n75162 , n75163 );
xor ( n75166 , n73991 , n74072 );
nor ( n75167 , n9608 , n74843 );
and ( n75168 , n75166 , n75167 );
xor ( n75169 , n75166 , n75167 );
xor ( n75170 , n73995 , n74070 );
nor ( n75171 , n9617 , n74843 );
and ( n75172 , n75170 , n75171 );
xor ( n75173 , n75170 , n75171 );
xor ( n75174 , n73999 , n74068 );
nor ( n75175 , n9626 , n74843 );
and ( n75176 , n75174 , n75175 );
xor ( n75177 , n75174 , n75175 );
xor ( n75178 , n74003 , n74066 );
nor ( n75179 , n9635 , n74843 );
and ( n75180 , n75178 , n75179 );
xor ( n75181 , n75178 , n75179 );
xor ( n75182 , n74007 , n74064 );
nor ( n75183 , n9644 , n74843 );
and ( n75184 , n75182 , n75183 );
xor ( n75185 , n75182 , n75183 );
xor ( n75186 , n74011 , n74062 );
nor ( n75187 , n9653 , n74843 );
and ( n75188 , n75186 , n75187 );
xor ( n75189 , n75186 , n75187 );
xor ( n75190 , n74015 , n74060 );
nor ( n75191 , n9662 , n74843 );
and ( n75192 , n75190 , n75191 );
xor ( n75193 , n75190 , n75191 );
xor ( n75194 , n74019 , n74058 );
nor ( n75195 , n9671 , n74843 );
and ( n75196 , n75194 , n75195 );
xor ( n75197 , n75194 , n75195 );
xor ( n75198 , n74023 , n74056 );
nor ( n75199 , n9680 , n74843 );
and ( n75200 , n75198 , n75199 );
xor ( n75201 , n75198 , n75199 );
xor ( n75202 , n74027 , n74054 );
nor ( n75203 , n9689 , n74843 );
and ( n75204 , n75202 , n75203 );
xor ( n75205 , n75202 , n75203 );
xor ( n75206 , n74031 , n74052 );
nor ( n75207 , n9698 , n74843 );
and ( n75208 , n75206 , n75207 );
xor ( n75209 , n75206 , n75207 );
xor ( n75210 , n74035 , n74050 );
nor ( n75211 , n9707 , n74843 );
and ( n75212 , n75210 , n75211 );
xor ( n75213 , n75210 , n75211 );
xor ( n75214 , n74039 , n74048 );
nor ( n75215 , n9716 , n74843 );
and ( n75216 , n75214 , n75215 );
xor ( n75217 , n75214 , n75215 );
xor ( n75218 , n74043 , n74046 );
nor ( n75219 , n9725 , n74843 );
and ( n75220 , n75218 , n75219 );
xor ( n75221 , n75218 , n75219 );
xor ( n75222 , n74044 , n74045 );
nor ( n75223 , n9734 , n74843 );
and ( n75224 , n75222 , n75223 );
xor ( n75225 , n75222 , n75223 );
nor ( n75226 , n9752 , n73665 );
nor ( n75227 , n9743 , n74843 );
and ( n75228 , n75226 , n75227 );
and ( n75229 , n75225 , n75228 );
or ( n75230 , n75224 , n75229 );
and ( n75231 , n75221 , n75230 );
or ( n75232 , n75220 , n75231 );
and ( n75233 , n75217 , n75232 );
or ( n75234 , n75216 , n75233 );
and ( n75235 , n75213 , n75234 );
or ( n75236 , n75212 , n75235 );
and ( n75237 , n75209 , n75236 );
or ( n75238 , n75208 , n75237 );
and ( n75239 , n75205 , n75238 );
or ( n75240 , n75204 , n75239 );
and ( n75241 , n75201 , n75240 );
or ( n75242 , n75200 , n75241 );
and ( n75243 , n75197 , n75242 );
or ( n75244 , n75196 , n75243 );
and ( n75245 , n75193 , n75244 );
or ( n75246 , n75192 , n75245 );
and ( n75247 , n75189 , n75246 );
or ( n75248 , n75188 , n75247 );
and ( n75249 , n75185 , n75248 );
or ( n75250 , n75184 , n75249 );
and ( n75251 , n75181 , n75250 );
or ( n75252 , n75180 , n75251 );
and ( n75253 , n75177 , n75252 );
or ( n75254 , n75176 , n75253 );
and ( n75255 , n75173 , n75254 );
or ( n75256 , n75172 , n75255 );
and ( n75257 , n75169 , n75256 );
or ( n75258 , n75168 , n75257 );
and ( n75259 , n75165 , n75258 );
or ( n75260 , n75164 , n75259 );
and ( n75261 , n75161 , n75260 );
or ( n75262 , n75160 , n75261 );
and ( n75263 , n75157 , n75262 );
or ( n75264 , n75156 , n75263 );
and ( n75265 , n75153 , n75264 );
or ( n75266 , n75152 , n75265 );
and ( n75267 , n75149 , n75266 );
or ( n75268 , n75148 , n75267 );
and ( n75269 , n75145 , n75268 );
or ( n75270 , n75144 , n75269 );
and ( n75271 , n75141 , n75270 );
or ( n75272 , n75140 , n75271 );
and ( n75273 , n75137 , n75272 );
or ( n75274 , n75136 , n75273 );
and ( n75275 , n75133 , n75274 );
or ( n75276 , n75132 , n75275 );
and ( n75277 , n75129 , n75276 );
or ( n75278 , n75128 , n75277 );
and ( n75279 , n75125 , n75278 );
or ( n75280 , n75124 , n75279 );
and ( n75281 , n75121 , n75280 );
or ( n75282 , n75120 , n75281 );
and ( n75283 , n75117 , n75282 );
or ( n75284 , n75116 , n75283 );
and ( n75285 , n75113 , n75284 );
or ( n75286 , n75112 , n75285 );
and ( n75287 , n75109 , n75286 );
or ( n75288 , n75108 , n75287 );
and ( n75289 , n75105 , n75288 );
or ( n75290 , n75104 , n75289 );
and ( n75291 , n75101 , n75290 );
or ( n75292 , n75100 , n75291 );
and ( n75293 , n75097 , n75292 );
or ( n75294 , n75096 , n75293 );
and ( n75295 , n75093 , n75294 );
or ( n75296 , n75092 , n75295 );
and ( n75297 , n75089 , n75296 );
or ( n75298 , n75088 , n75297 );
and ( n75299 , n75085 , n75298 );
or ( n75300 , n75084 , n75299 );
and ( n75301 , n75081 , n75300 );
or ( n75302 , n75080 , n75301 );
and ( n75303 , n75077 , n75302 );
or ( n75304 , n75076 , n75303 );
and ( n75305 , n75073 , n75304 );
or ( n75306 , n75072 , n75305 );
and ( n75307 , n75069 , n75306 );
or ( n75308 , n75068 , n75307 );
and ( n75309 , n75065 , n75308 );
or ( n75310 , n75064 , n75309 );
and ( n75311 , n75061 , n75310 );
or ( n75312 , n75060 , n75311 );
and ( n75313 , n75057 , n75312 );
or ( n75314 , n75056 , n75313 );
and ( n75315 , n75053 , n75314 );
or ( n75316 , n75052 , n75315 );
and ( n75317 , n75049 , n75316 );
or ( n75318 , n75048 , n75317 );
and ( n75319 , n75045 , n75318 );
or ( n75320 , n75044 , n75319 );
and ( n75321 , n75041 , n75320 );
or ( n75322 , n75040 , n75321 );
and ( n75323 , n75037 , n75322 );
or ( n75324 , n75036 , n75323 );
and ( n75325 , n75033 , n75324 );
or ( n75326 , n75032 , n75325 );
and ( n75327 , n75029 , n75326 );
or ( n75328 , n75028 , n75327 );
and ( n75329 , n75025 , n75328 );
or ( n75330 , n75024 , n75329 );
and ( n75331 , n75021 , n75330 );
or ( n75332 , n75020 , n75331 );
and ( n75333 , n75017 , n75332 );
or ( n75334 , n75016 , n75333 );
and ( n75335 , n75013 , n75334 );
or ( n75336 , n75012 , n75335 );
and ( n75337 , n75009 , n75336 );
or ( n75338 , n75008 , n75337 );
and ( n75339 , n75005 , n75338 );
or ( n75340 , n75004 , n75339 );
and ( n75341 , n75001 , n75340 );
or ( n75342 , n75000 , n75341 );
and ( n75343 , n74997 , n75342 );
or ( n75344 , n74996 , n75343 );
and ( n75345 , n74993 , n75344 );
or ( n75346 , n74992 , n75345 );
and ( n75347 , n74989 , n75346 );
or ( n75348 , n74988 , n75347 );
and ( n75349 , n74985 , n75348 );
or ( n75350 , n74984 , n75349 );
and ( n75351 , n74981 , n75350 );
or ( n75352 , n74980 , n75351 );
and ( n75353 , n74977 , n75352 );
or ( n75354 , n74976 , n75353 );
and ( n75355 , n74973 , n75354 );
or ( n75356 , n74972 , n75355 );
and ( n75357 , n74969 , n75356 );
or ( n75358 , n74968 , n75357 );
and ( n75359 , n74965 , n75358 );
or ( n75360 , n74964 , n75359 );
and ( n75361 , n74961 , n75360 );
or ( n75362 , n74960 , n75361 );
and ( n75363 , n74957 , n75362 );
or ( n75364 , n74956 , n75363 );
and ( n75365 , n74953 , n75364 );
or ( n75366 , n74952 , n75365 );
and ( n75367 , n74949 , n75366 );
or ( n75368 , n74948 , n75367 );
and ( n75369 , n74945 , n75368 );
or ( n75370 , n74944 , n75369 );
and ( n75371 , n74941 , n75370 );
or ( n75372 , n74940 , n75371 );
and ( n75373 , n74937 , n75372 );
or ( n75374 , n74936 , n75373 );
and ( n75375 , n74933 , n75374 );
or ( n75376 , n74932 , n75375 );
and ( n75377 , n74929 , n75376 );
or ( n75378 , n74928 , n75377 );
and ( n75379 , n74925 , n75378 );
or ( n75380 , n74924 , n75379 );
and ( n75381 , n74921 , n75380 );
or ( n75382 , n74920 , n75381 );
and ( n75383 , n74917 , n75382 );
or ( n75384 , n74916 , n75383 );
and ( n75385 , n74913 , n75384 );
or ( n75386 , n74912 , n75385 );
and ( n75387 , n74909 , n75386 );
or ( n75388 , n74908 , n75387 );
and ( n75389 , n74905 , n75388 );
or ( n75390 , n74904 , n75389 );
and ( n75391 , n74901 , n75390 );
or ( n75392 , n74900 , n75391 );
and ( n75393 , n74897 , n75392 );
or ( n75394 , n74896 , n75393 );
and ( n75395 , n74893 , n75394 );
or ( n75396 , n74892 , n75395 );
and ( n75397 , n74889 , n75396 );
or ( n75398 , n74888 , n75397 );
and ( n75399 , n74885 , n75398 );
or ( n75400 , n74884 , n75399 );
and ( n75401 , n74881 , n75400 );
or ( n75402 , n74880 , n75401 );
and ( n75403 , n74877 , n75402 );
or ( n75404 , n74876 , n75403 );
and ( n75405 , n74873 , n75404 );
or ( n75406 , n74872 , n75405 );
and ( n75407 , n74869 , n75406 );
or ( n75408 , n74868 , n75407 );
and ( n75409 , n74865 , n75408 );
or ( n75410 , n74864 , n75409 );
and ( n75411 , n74861 , n75410 );
or ( n75412 , n74860 , n75411 );
and ( n75413 , n74857 , n75412 );
or ( n75414 , n74856 , n75413 );
and ( n75415 , n74853 , n75414 );
or ( n75416 , n74852 , n75415 );
and ( n75417 , n74849 , n75416 );
or ( n75418 , n74848 , n75417 );
xor ( n75419 , n74845 , n75418 );
and ( n75420 , n33403 , n8280 );
nor ( n75421 , n8281 , n75420 );
nor ( n75422 , n8737 , n32231 );
xor ( n75423 , n75421 , n75422 );
and ( n75424 , n74237 , n74238 );
and ( n75425 , n74239 , n74242 );
or ( n75426 , n75424 , n75425 );
xor ( n75427 , n75423 , n75426 );
nor ( n75428 , n9420 , n31083 );
xor ( n75429 , n75427 , n75428 );
and ( n75430 , n74243 , n74244 );
and ( n75431 , n74245 , n74248 );
or ( n75432 , n75430 , n75431 );
xor ( n75433 , n75429 , n75432 );
nor ( n75434 , n10312 , n29948 );
xor ( n75435 , n75433 , n75434 );
and ( n75436 , n74249 , n74250 );
and ( n75437 , n74251 , n74254 );
or ( n75438 , n75436 , n75437 );
xor ( n75439 , n75435 , n75438 );
nor ( n75440 , n11041 , n28833 );
xor ( n75441 , n75439 , n75440 );
and ( n75442 , n74255 , n74256 );
and ( n75443 , n74257 , n74260 );
or ( n75444 , n75442 , n75443 );
xor ( n75445 , n75441 , n75444 );
nor ( n75446 , n11790 , n27737 );
xor ( n75447 , n75445 , n75446 );
and ( n75448 , n74261 , n74262 );
and ( n75449 , n74263 , n74266 );
or ( n75450 , n75448 , n75449 );
xor ( n75451 , n75447 , n75450 );
nor ( n75452 , n12555 , n26660 );
xor ( n75453 , n75451 , n75452 );
and ( n75454 , n74267 , n74268 );
and ( n75455 , n74269 , n74272 );
or ( n75456 , n75454 , n75455 );
xor ( n75457 , n75453 , n75456 );
nor ( n75458 , n13340 , n25600 );
xor ( n75459 , n75457 , n75458 );
and ( n75460 , n74273 , n74274 );
and ( n75461 , n74275 , n74278 );
or ( n75462 , n75460 , n75461 );
xor ( n75463 , n75459 , n75462 );
nor ( n75464 , n14138 , n24564 );
xor ( n75465 , n75463 , n75464 );
and ( n75466 , n74279 , n74280 );
and ( n75467 , n74281 , n74284 );
or ( n75468 , n75466 , n75467 );
xor ( n75469 , n75465 , n75468 );
nor ( n75470 , n14959 , n23541 );
xor ( n75471 , n75469 , n75470 );
and ( n75472 , n74285 , n74286 );
and ( n75473 , n74287 , n74290 );
or ( n75474 , n75472 , n75473 );
xor ( n75475 , n75471 , n75474 );
nor ( n75476 , n15800 , n22541 );
xor ( n75477 , n75475 , n75476 );
and ( n75478 , n74291 , n74292 );
and ( n75479 , n74293 , n74296 );
or ( n75480 , n75478 , n75479 );
xor ( n75481 , n75477 , n75480 );
nor ( n75482 , n16660 , n21562 );
xor ( n75483 , n75481 , n75482 );
and ( n75484 , n74297 , n74298 );
and ( n75485 , n74299 , n74302 );
or ( n75486 , n75484 , n75485 );
xor ( n75487 , n75483 , n75486 );
nor ( n75488 , n17539 , n20601 );
xor ( n75489 , n75487 , n75488 );
and ( n75490 , n74303 , n74304 );
and ( n75491 , n74305 , n74308 );
or ( n75492 , n75490 , n75491 );
xor ( n75493 , n75489 , n75492 );
nor ( n75494 , n18439 , n19657 );
xor ( n75495 , n75493 , n75494 );
and ( n75496 , n74309 , n74310 );
and ( n75497 , n74311 , n74314 );
or ( n75498 , n75496 , n75497 );
xor ( n75499 , n75495 , n75498 );
nor ( n75500 , n19356 , n18734 );
xor ( n75501 , n75499 , n75500 );
and ( n75502 , n74315 , n74316 );
and ( n75503 , n74317 , n74320 );
or ( n75504 , n75502 , n75503 );
xor ( n75505 , n75501 , n75504 );
nor ( n75506 , n20294 , n17828 );
xor ( n75507 , n75505 , n75506 );
and ( n75508 , n74321 , n74322 );
and ( n75509 , n74323 , n74326 );
or ( n75510 , n75508 , n75509 );
xor ( n75511 , n75507 , n75510 );
nor ( n75512 , n21249 , n16943 );
xor ( n75513 , n75511 , n75512 );
and ( n75514 , n74327 , n74328 );
and ( n75515 , n74329 , n74332 );
or ( n75516 , n75514 , n75515 );
xor ( n75517 , n75513 , n75516 );
nor ( n75518 , n22222 , n16077 );
xor ( n75519 , n75517 , n75518 );
and ( n75520 , n74333 , n74334 );
and ( n75521 , n74335 , n74338 );
or ( n75522 , n75520 , n75521 );
xor ( n75523 , n75519 , n75522 );
nor ( n75524 , n23216 , n15230 );
xor ( n75525 , n75523 , n75524 );
and ( n75526 , n74339 , n74340 );
and ( n75527 , n74341 , n74344 );
or ( n75528 , n75526 , n75527 );
xor ( n75529 , n75525 , n75528 );
nor ( n75530 , n24233 , n14403 );
xor ( n75531 , n75529 , n75530 );
and ( n75532 , n74345 , n74346 );
and ( n75533 , n74347 , n74350 );
or ( n75534 , n75532 , n75533 );
xor ( n75535 , n75531 , n75534 );
nor ( n75536 , n25263 , n13599 );
xor ( n75537 , n75535 , n75536 );
and ( n75538 , n74351 , n74352 );
and ( n75539 , n74353 , n74356 );
or ( n75540 , n75538 , n75539 );
xor ( n75541 , n75537 , n75540 );
nor ( n75542 , n26317 , n12808 );
xor ( n75543 , n75541 , n75542 );
and ( n75544 , n74357 , n74358 );
and ( n75545 , n74359 , n74362 );
or ( n75546 , n75544 , n75545 );
xor ( n75547 , n75543 , n75546 );
nor ( n75548 , n27388 , n12037 );
xor ( n75549 , n75547 , n75548 );
and ( n75550 , n74363 , n74364 );
and ( n75551 , n74365 , n74368 );
or ( n75552 , n75550 , n75551 );
xor ( n75553 , n75549 , n75552 );
nor ( n75554 , n28478 , n11282 );
xor ( n75555 , n75553 , n75554 );
and ( n75556 , n74369 , n74370 );
and ( n75557 , n74371 , n74374 );
or ( n75558 , n75556 , n75557 );
xor ( n75559 , n75555 , n75558 );
nor ( n75560 , n29587 , n10547 );
xor ( n75561 , n75559 , n75560 );
and ( n75562 , n74375 , n74376 );
and ( n75563 , n74377 , n74380 );
or ( n75564 , n75562 , n75563 );
xor ( n75565 , n75561 , n75564 );
nor ( n75566 , n30716 , n9829 );
xor ( n75567 , n75565 , n75566 );
and ( n75568 , n74381 , n74382 );
and ( n75569 , n74383 , n74386 );
or ( n75570 , n75568 , n75569 );
xor ( n75571 , n75567 , n75570 );
nor ( n75572 , n31858 , n8955 );
xor ( n75573 , n75571 , n75572 );
and ( n75574 , n74387 , n74388 );
and ( n75575 , n74389 , n74392 );
or ( n75576 , n75574 , n75575 );
xor ( n75577 , n75573 , n75576 );
nor ( n75578 , n33024 , n603 );
xor ( n75579 , n75577 , n75578 );
and ( n75580 , n74393 , n74394 );
and ( n75581 , n74395 , n74398 );
or ( n75582 , n75580 , n75581 );
xor ( n75583 , n75579 , n75582 );
nor ( n75584 , n34215 , n652 );
xor ( n75585 , n75583 , n75584 );
and ( n75586 , n74399 , n74400 );
and ( n75587 , n74401 , n74404 );
or ( n75588 , n75586 , n75587 );
xor ( n75589 , n75585 , n75588 );
nor ( n75590 , n35410 , n624 );
xor ( n75591 , n75589 , n75590 );
and ( n75592 , n74405 , n74406 );
and ( n75593 , n74407 , n74410 );
or ( n75594 , n75592 , n75593 );
xor ( n75595 , n75591 , n75594 );
nor ( n75596 , n36611 , n648 );
xor ( n75597 , n75595 , n75596 );
and ( n75598 , n74411 , n74412 );
and ( n75599 , n74413 , n74416 );
or ( n75600 , n75598 , n75599 );
xor ( n75601 , n75597 , n75600 );
nor ( n75602 , n37816 , n686 );
xor ( n75603 , n75601 , n75602 );
and ( n75604 , n74417 , n74418 );
and ( n75605 , n74419 , n74422 );
or ( n75606 , n75604 , n75605 );
xor ( n75607 , n75603 , n75606 );
nor ( n75608 , n39018 , n735 );
xor ( n75609 , n75607 , n75608 );
and ( n75610 , n74423 , n74424 );
and ( n75611 , n74425 , n74428 );
or ( n75612 , n75610 , n75611 );
xor ( n75613 , n75609 , n75612 );
nor ( n75614 , n40223 , n798 );
xor ( n75615 , n75613 , n75614 );
and ( n75616 , n74429 , n74430 );
and ( n75617 , n74431 , n74434 );
or ( n75618 , n75616 , n75617 );
xor ( n75619 , n75615 , n75618 );
nor ( n75620 , n41428 , n870 );
xor ( n75621 , n75619 , n75620 );
and ( n75622 , n74435 , n74436 );
and ( n75623 , n74437 , n74440 );
or ( n75624 , n75622 , n75623 );
xor ( n75625 , n75621 , n75624 );
nor ( n75626 , n42632 , n960 );
xor ( n75627 , n75625 , n75626 );
and ( n75628 , n74441 , n74442 );
and ( n75629 , n74443 , n74446 );
or ( n75630 , n75628 , n75629 );
xor ( n75631 , n75627 , n75630 );
nor ( n75632 , n43834 , n1064 );
xor ( n75633 , n75631 , n75632 );
and ( n75634 , n74447 , n74448 );
and ( n75635 , n74449 , n74452 );
or ( n75636 , n75634 , n75635 );
xor ( n75637 , n75633 , n75636 );
nor ( n75638 , n45038 , n1178 );
xor ( n75639 , n75637 , n75638 );
and ( n75640 , n74453 , n74454 );
and ( n75641 , n74455 , n74458 );
or ( n75642 , n75640 , n75641 );
xor ( n75643 , n75639 , n75642 );
nor ( n75644 , n46239 , n1305 );
xor ( n75645 , n75643 , n75644 );
and ( n75646 , n74459 , n74460 );
and ( n75647 , n74461 , n74464 );
or ( n75648 , n75646 , n75647 );
xor ( n75649 , n75645 , n75648 );
nor ( n75650 , n47440 , n1447 );
xor ( n75651 , n75649 , n75650 );
and ( n75652 , n74465 , n74466 );
and ( n75653 , n74467 , n74470 );
or ( n75654 , n75652 , n75653 );
xor ( n75655 , n75651 , n75654 );
nor ( n75656 , n48641 , n1600 );
xor ( n75657 , n75655 , n75656 );
and ( n75658 , n74471 , n74472 );
and ( n75659 , n74473 , n74476 );
or ( n75660 , n75658 , n75659 );
xor ( n75661 , n75657 , n75660 );
nor ( n75662 , n49841 , n1768 );
xor ( n75663 , n75661 , n75662 );
and ( n75664 , n74477 , n74478 );
and ( n75665 , n74479 , n74482 );
or ( n75666 , n75664 , n75665 );
xor ( n75667 , n75663 , n75666 );
nor ( n75668 , n51040 , n1947 );
xor ( n75669 , n75667 , n75668 );
and ( n75670 , n74483 , n74484 );
and ( n75671 , n74485 , n74488 );
or ( n75672 , n75670 , n75671 );
xor ( n75673 , n75669 , n75672 );
nor ( n75674 , n52238 , n2139 );
xor ( n75675 , n75673 , n75674 );
and ( n75676 , n74489 , n74490 );
and ( n75677 , n74491 , n74494 );
or ( n75678 , n75676 , n75677 );
xor ( n75679 , n75675 , n75678 );
nor ( n75680 , n53432 , n2345 );
xor ( n75681 , n75679 , n75680 );
and ( n75682 , n74495 , n74496 );
and ( n75683 , n74497 , n74500 );
or ( n75684 , n75682 , n75683 );
xor ( n75685 , n75681 , n75684 );
nor ( n75686 , n54629 , n2568 );
xor ( n75687 , n75685 , n75686 );
and ( n75688 , n74501 , n74502 );
and ( n75689 , n74503 , n74506 );
or ( n75690 , n75688 , n75689 );
xor ( n75691 , n75687 , n75690 );
nor ( n75692 , n55826 , n2799 );
xor ( n75693 , n75691 , n75692 );
and ( n75694 , n74507 , n74508 );
and ( n75695 , n74509 , n74512 );
or ( n75696 , n75694 , n75695 );
xor ( n75697 , n75693 , n75696 );
nor ( n75698 , n57022 , n3045 );
xor ( n75699 , n75697 , n75698 );
and ( n75700 , n74513 , n74514 );
and ( n75701 , n74515 , n74518 );
or ( n75702 , n75700 , n75701 );
xor ( n75703 , n75699 , n75702 );
nor ( n75704 , n58217 , n3302 );
xor ( n75705 , n75703 , n75704 );
and ( n75706 , n74519 , n74520 );
and ( n75707 , n74521 , n74524 );
or ( n75708 , n75706 , n75707 );
xor ( n75709 , n75705 , n75708 );
nor ( n75710 , n59412 , n3572 );
xor ( n75711 , n75709 , n75710 );
and ( n75712 , n74525 , n74526 );
and ( n75713 , n74527 , n74530 );
or ( n75714 , n75712 , n75713 );
xor ( n75715 , n75711 , n75714 );
nor ( n75716 , n60600 , n3855 );
xor ( n75717 , n75715 , n75716 );
and ( n75718 , n74531 , n74532 );
and ( n75719 , n74533 , n74536 );
or ( n75720 , n75718 , n75719 );
xor ( n75721 , n75717 , n75720 );
nor ( n75722 , n61791 , n4153 );
xor ( n75723 , n75721 , n75722 );
and ( n75724 , n74537 , n74538 );
and ( n75725 , n74539 , n74542 );
or ( n75726 , n75724 , n75725 );
xor ( n75727 , n75723 , n75726 );
nor ( n75728 , n62982 , n4460 );
xor ( n75729 , n75727 , n75728 );
and ( n75730 , n74543 , n74544 );
and ( n75731 , n74545 , n74548 );
or ( n75732 , n75730 , n75731 );
xor ( n75733 , n75729 , n75732 );
nor ( n75734 , n64172 , n4788 );
xor ( n75735 , n75733 , n75734 );
and ( n75736 , n74549 , n74550 );
and ( n75737 , n74551 , n74554 );
or ( n75738 , n75736 , n75737 );
xor ( n75739 , n75735 , n75738 );
nor ( n75740 , n65360 , n5128 );
xor ( n75741 , n75739 , n75740 );
and ( n75742 , n74555 , n74556 );
and ( n75743 , n74557 , n74560 );
or ( n75744 , n75742 , n75743 );
xor ( n75745 , n75741 , n75744 );
nor ( n75746 , n66550 , n5479 );
xor ( n75747 , n75745 , n75746 );
and ( n75748 , n74561 , n74562 );
and ( n75749 , n74563 , n74566 );
or ( n75750 , n75748 , n75749 );
xor ( n75751 , n75747 , n75750 );
nor ( n75752 , n67736 , n5840 );
xor ( n75753 , n75751 , n75752 );
and ( n75754 , n74567 , n74568 );
and ( n75755 , n74569 , n74572 );
or ( n75756 , n75754 , n75755 );
xor ( n75757 , n75753 , n75756 );
nor ( n75758 , n68924 , n6214 );
xor ( n75759 , n75757 , n75758 );
and ( n75760 , n74573 , n74574 );
and ( n75761 , n74575 , n74578 );
or ( n75762 , n75760 , n75761 );
xor ( n75763 , n75759 , n75762 );
nor ( n75764 , n70110 , n6598 );
xor ( n75765 , n75763 , n75764 );
and ( n75766 , n74579 , n74580 );
and ( n75767 , n74581 , n74584 );
or ( n75768 , n75766 , n75767 );
xor ( n75769 , n75765 , n75768 );
nor ( n75770 , n71292 , n6999 );
xor ( n75771 , n75769 , n75770 );
and ( n75772 , n74585 , n74586 );
and ( n75773 , n74587 , n74590 );
or ( n75774 , n75772 , n75773 );
xor ( n75775 , n75771 , n75774 );
nor ( n75776 , n72472 , n7415 );
xor ( n75777 , n75775 , n75776 );
and ( n75778 , n74591 , n74592 );
and ( n75779 , n74593 , n74596 );
or ( n75780 , n75778 , n75779 );
xor ( n75781 , n75777 , n75780 );
nor ( n75782 , n73654 , n7843 );
xor ( n75783 , n75781 , n75782 );
and ( n75784 , n74597 , n74598 );
and ( n75785 , n74599 , n74602 );
or ( n75786 , n75784 , n75785 );
xor ( n75787 , n75783 , n75786 );
nor ( n75788 , n74832 , n8283 );
xor ( n75789 , n75787 , n75788 );
and ( n75790 , n74603 , n74604 );
and ( n75791 , n74605 , n74608 );
or ( n75792 , n75790 , n75791 );
xor ( n75793 , n75789 , n75792 );
and ( n75794 , n74621 , n74625 );
and ( n75795 , n74625 , n74818 );
and ( n75796 , n74621 , n74818 );
or ( n75797 , n75794 , n75795 , n75796 );
and ( n75798 , n33774 , n8243 );
not ( n75799 , n8243 );
nor ( n75800 , n75798 , n75799 );
xor ( n75801 , n75797 , n75800 );
and ( n75802 , n74631 , n74632 );
and ( n75803 , n74632 , n74700 );
and ( n75804 , n74631 , n74700 );
or ( n75805 , n75802 , n75803 , n75804 );
and ( n75806 , n74627 , n74701 );
and ( n75807 , n74701 , n74817 );
and ( n75808 , n74627 , n74817 );
or ( n75809 , n75806 , n75807 , n75808 );
xor ( n75810 , n75805 , n75809 );
and ( n75811 , n74712 , n74816 );
and ( n75812 , n74637 , n74641 );
and ( n75813 , n74641 , n74699 );
and ( n75814 , n74637 , n74699 );
or ( n75815 , n75812 , n75813 , n75814 );
and ( n75816 , n74716 , n74815 );
xor ( n75817 , n75815 , n75816 );
and ( n75818 , n74668 , n74672 );
and ( n75819 , n74672 , n74678 );
and ( n75820 , n74668 , n74678 );
or ( n75821 , n75818 , n75819 , n75820 );
and ( n75822 , n74646 , n74650 );
and ( n75823 , n74650 , n74698 );
and ( n75824 , n74646 , n74698 );
or ( n75825 , n75822 , n75823 , n75824 );
xor ( n75826 , n75821 , n75825 );
and ( n75827 , n74655 , n74659 );
and ( n75828 , n74659 , n74697 );
and ( n75829 , n74655 , n74697 );
or ( n75830 , n75827 , n75828 , n75829 );
and ( n75831 , n74724 , n74749 );
and ( n75832 , n74749 , n74784 );
and ( n75833 , n74724 , n74784 );
or ( n75834 , n75831 , n75832 , n75833 );
xor ( n75835 , n75830 , n75834 );
and ( n75836 , n74664 , n74679 );
and ( n75837 , n74679 , n74696 );
and ( n75838 , n74664 , n74696 );
or ( n75839 , n75836 , n75837 , n75838 );
and ( n75840 , n74728 , n74732 );
and ( n75841 , n74732 , n74748 );
and ( n75842 , n74728 , n74748 );
or ( n75843 , n75840 , n75841 , n75842 );
xor ( n75844 , n75839 , n75843 );
and ( n75845 , n74684 , n74689 );
and ( n75846 , n74689 , n74695 );
and ( n75847 , n74684 , n74695 );
or ( n75848 , n75845 , n75846 , n75847 );
and ( n75849 , n74674 , n74675 );
and ( n75850 , n74675 , n74677 );
and ( n75851 , n74674 , n74677 );
or ( n75852 , n75849 , n75850 , n75851 );
and ( n75853 , n74685 , n74686 );
and ( n75854 , n74686 , n74688 );
and ( n75855 , n74685 , n74688 );
or ( n75856 , n75853 , n75854 , n75855 );
xor ( n75857 , n75852 , n75856 );
and ( n75858 , n30695 , n10239 );
and ( n75859 , n31836 , n9348 );
xor ( n75860 , n75858 , n75859 );
and ( n75861 , n32649 , n8669 );
xor ( n75862 , n75860 , n75861 );
xor ( n75863 , n75857 , n75862 );
xor ( n75864 , n75848 , n75863 );
and ( n75865 , n74691 , n74692 );
and ( n75866 , n74692 , n74694 );
and ( n75867 , n74691 , n74694 );
or ( n75868 , n75865 , n75866 , n75867 );
and ( n75869 , n27361 , n12531 );
and ( n75870 , n28456 , n11718 );
xor ( n75871 , n75869 , n75870 );
and ( n75872 , n29559 , n10977 );
xor ( n75873 , n75871 , n75872 );
xor ( n75874 , n75868 , n75873 );
and ( n75875 , n24214 , n14838 );
and ( n75876 , n25243 , n14044 );
xor ( n75877 , n75875 , n75876 );
and ( n75878 , n26296 , n13256 );
xor ( n75879 , n75877 , n75878 );
xor ( n75880 , n75874 , n75879 );
xor ( n75881 , n75864 , n75880 );
xor ( n75882 , n75844 , n75881 );
xor ( n75883 , n75835 , n75882 );
xor ( n75884 , n75826 , n75883 );
xor ( n75885 , n75817 , n75884 );
xor ( n75886 , n75811 , n75885 );
and ( n75887 , n74709 , n74710 );
not ( n75888 , n8079 );
and ( n75889 , n34193 , n8079 );
nor ( n75890 , n75888 , n75889 );
xor ( n75891 , n75887 , n75890 );
and ( n75892 , n74720 , n74785 );
and ( n75893 , n74785 , n74814 );
and ( n75894 , n74720 , n74814 );
or ( n75895 , n75892 , n75893 , n75894 );
and ( n75896 , n74790 , n74813 );
and ( n75897 , n74754 , n74767 );
and ( n75898 , n74767 , n74783 );
and ( n75899 , n74754 , n74783 );
or ( n75900 , n75897 , n75898 , n75899 );
and ( n75901 , n74737 , n74741 );
and ( n75902 , n74741 , n74747 );
and ( n75903 , n74737 , n74747 );
or ( n75904 , n75901 , n75902 , n75903 );
and ( n75905 , n74758 , n74763 );
and ( n75906 , n74763 , n74766 );
and ( n75907 , n74758 , n74766 );
or ( n75908 , n75905 , n75906 , n75907 );
xor ( n75909 , n75904 , n75908 );
and ( n75910 , n74743 , n74744 );
and ( n75911 , n74744 , n74746 );
and ( n75912 , n74743 , n74746 );
or ( n75913 , n75910 , n75911 , n75912 );
and ( n75914 , n18144 , n19222 );
and ( n75915 , n19324 , n18407 );
and ( n75916 , n75914 , n75915 );
and ( n75917 , n75915 , n74765 );
and ( n75918 , n75914 , n74765 );
or ( n75919 , n75916 , n75917 , n75918 );
xor ( n75920 , n75913 , n75919 );
and ( n75921 , n21216 , n17422 );
and ( n75922 , n22186 , n16550 );
xor ( n75923 , n75921 , n75922 );
and ( n75924 , n22892 , n15691 );
xor ( n75925 , n75923 , n75924 );
xor ( n75926 , n75920 , n75925 );
xor ( n75927 , n75909 , n75926 );
xor ( n75928 , n75900 , n75927 );
and ( n75929 , n74772 , n74776 );
and ( n75930 , n74776 , n74782 );
and ( n75931 , n74772 , n74782 );
or ( n75932 , n75929 , n75930 , n75931 );
and ( n75933 , n74759 , n74760 );
and ( n75934 , n74760 , n74762 );
and ( n75935 , n74759 , n74762 );
or ( n75936 , n75933 , n75934 , n75935 );
and ( n75937 , n18144 , n20156 );
buf ( n75938 , n19324 );
xor ( n75939 , n75937 , n75938 );
and ( n75940 , n20233 , n18407 );
xor ( n75941 , n75939 , n75940 );
xor ( n75942 , n75936 , n75941 );
and ( n75943 , n15758 , n23075 );
and ( n75944 , n16637 , n22065 );
xor ( n75945 , n75943 , n75944 );
and ( n75946 , n17512 , n20976 );
xor ( n75947 , n75945 , n75946 );
xor ( n75948 , n75942 , n75947 );
xor ( n75949 , n75932 , n75948 );
and ( n75950 , n74807 , n74808 );
and ( n75951 , n74808 , n74810 );
and ( n75952 , n74807 , n74810 );
or ( n75953 , n75950 , n75951 , n75952 );
and ( n75954 , n74778 , n74779 );
and ( n75955 , n74779 , n74781 );
and ( n75956 , n74778 , n74781 );
or ( n75957 , n75954 , n75955 , n75956 );
xor ( n75958 , n75953 , n75957 );
and ( n75959 , n13322 , n26216 );
and ( n75960 , n14118 , n25163 );
xor ( n75961 , n75959 , n75960 );
and ( n75962 , n14938 , n24137 );
xor ( n75963 , n75961 , n75962 );
xor ( n75964 , n75958 , n75963 );
xor ( n75965 , n75949 , n75964 );
xor ( n75966 , n75928 , n75965 );
xor ( n75967 , n75896 , n75966 );
and ( n75968 , n74794 , n74795 );
and ( n75969 , n74795 , n74812 );
and ( n75970 , n74794 , n74812 );
or ( n75971 , n75968 , n75969 , n75970 );
and ( n75972 , n74800 , n74805 );
and ( n75973 , n74805 , n74811 );
and ( n75974 , n74800 , n74811 );
or ( n75975 , n75972 , n75973 , n75974 );
and ( n75976 , n74706 , n74711 );
xor ( n75977 , n75975 , n75976 );
and ( n75978 , n74801 , n74802 );
and ( n75979 , n74802 , n74804 );
and ( n75980 , n74801 , n74804 );
or ( n75981 , n75978 , n75979 , n75980 );
and ( n75982 , n11015 , n29508 );
and ( n75983 , n11769 , n28406 );
xor ( n75984 , n75982 , n75983 );
and ( n75985 , n12320 , n27296 );
xor ( n75986 , n75984 , n75985 );
xor ( n75987 , n75981 , n75986 );
and ( n75988 , n8718 , n32999 );
and ( n75989 , n9400 , n31761 );
xor ( n75990 , n75988 , n75989 );
and ( n75991 , n10291 , n30629 );
xor ( n75992 , n75990 , n75991 );
xor ( n75993 , n75987 , n75992 );
xor ( n75994 , n75977 , n75993 );
xor ( n75995 , n75971 , n75994 );
xor ( n75996 , n75967 , n75995 );
xor ( n75997 , n75895 , n75996 );
xor ( n75998 , n75891 , n75997 );
xor ( n75999 , n75886 , n75998 );
xor ( n76000 , n75810 , n75999 );
xor ( n76001 , n75801 , n76000 );
and ( n76002 , n74613 , n74616 );
and ( n76003 , n74616 , n74819 );
and ( n76004 , n74613 , n74819 );
or ( n76005 , n76002 , n76003 , n76004 );
xor ( n76006 , n76001 , n76005 );
and ( n76007 , n74820 , n74824 );
and ( n76008 , n74825 , n74828 );
or ( n76009 , n76007 , n76008 );
xor ( n76010 , n76006 , n76009 );
buf ( n76011 , n76010 );
buf ( n76012 , n76011 );
not ( n76013 , n76012 );
nor ( n76014 , n76013 , n8739 );
xor ( n76015 , n75793 , n76014 );
and ( n76016 , n74609 , n74833 );
and ( n76017 , n74834 , n74837 );
or ( n76018 , n76016 , n76017 );
xor ( n76019 , n76015 , n76018 );
buf ( n76020 , n76019 );
buf ( n76021 , n76020 );
not ( n76022 , n76021 );
buf ( n76023 , n597 );
not ( n76024 , n76023 );
nor ( n76025 , n76022 , n76024 );
xor ( n76026 , n75419 , n76025 );
xor ( n76027 , n74849 , n75416 );
nor ( n76028 , n74841 , n76024 );
and ( n76029 , n76027 , n76028 );
xor ( n76030 , n76027 , n76028 );
xor ( n76031 , n74853 , n75414 );
nor ( n76032 , n73663 , n76024 );
and ( n76033 , n76031 , n76032 );
xor ( n76034 , n76031 , n76032 );
xor ( n76035 , n74857 , n75412 );
nor ( n76036 , n72481 , n76024 );
and ( n76037 , n76035 , n76036 );
xor ( n76038 , n76035 , n76036 );
xor ( n76039 , n74861 , n75410 );
nor ( n76040 , n71301 , n76024 );
and ( n76041 , n76039 , n76040 );
xor ( n76042 , n76039 , n76040 );
xor ( n76043 , n74865 , n75408 );
nor ( n76044 , n70119 , n76024 );
and ( n76045 , n76043 , n76044 );
xor ( n76046 , n76043 , n76044 );
xor ( n76047 , n74869 , n75406 );
nor ( n76048 , n68933 , n76024 );
and ( n76049 , n76047 , n76048 );
xor ( n76050 , n76047 , n76048 );
xor ( n76051 , n74873 , n75404 );
nor ( n76052 , n67745 , n76024 );
and ( n76053 , n76051 , n76052 );
xor ( n76054 , n76051 , n76052 );
xor ( n76055 , n74877 , n75402 );
nor ( n76056 , n66559 , n76024 );
and ( n76057 , n76055 , n76056 );
xor ( n76058 , n76055 , n76056 );
xor ( n76059 , n74881 , n75400 );
nor ( n76060 , n65369 , n76024 );
and ( n76061 , n76059 , n76060 );
xor ( n76062 , n76059 , n76060 );
xor ( n76063 , n74885 , n75398 );
nor ( n76064 , n64181 , n76024 );
and ( n76065 , n76063 , n76064 );
xor ( n76066 , n76063 , n76064 );
xor ( n76067 , n74889 , n75396 );
nor ( n76068 , n62991 , n76024 );
and ( n76069 , n76067 , n76068 );
xor ( n76070 , n76067 , n76068 );
xor ( n76071 , n74893 , n75394 );
nor ( n76072 , n61800 , n76024 );
and ( n76073 , n76071 , n76072 );
xor ( n76074 , n76071 , n76072 );
xor ( n76075 , n74897 , n75392 );
nor ( n76076 , n60609 , n76024 );
and ( n76077 , n76075 , n76076 );
xor ( n76078 , n76075 , n76076 );
xor ( n76079 , n74901 , n75390 );
nor ( n76080 , n59421 , n76024 );
and ( n76081 , n76079 , n76080 );
xor ( n76082 , n76079 , n76080 );
xor ( n76083 , n74905 , n75388 );
nor ( n76084 , n58226 , n76024 );
and ( n76085 , n76083 , n76084 );
xor ( n76086 , n76083 , n76084 );
xor ( n76087 , n74909 , n75386 );
nor ( n76088 , n57031 , n76024 );
and ( n76089 , n76087 , n76088 );
xor ( n76090 , n76087 , n76088 );
xor ( n76091 , n74913 , n75384 );
nor ( n76092 , n55835 , n76024 );
and ( n76093 , n76091 , n76092 );
xor ( n76094 , n76091 , n76092 );
xor ( n76095 , n74917 , n75382 );
nor ( n76096 , n54638 , n76024 );
and ( n76097 , n76095 , n76096 );
xor ( n76098 , n76095 , n76096 );
xor ( n76099 , n74921 , n75380 );
nor ( n76100 , n53441 , n76024 );
and ( n76101 , n76099 , n76100 );
xor ( n76102 , n76099 , n76100 );
xor ( n76103 , n74925 , n75378 );
nor ( n76104 , n52247 , n76024 );
and ( n76105 , n76103 , n76104 );
xor ( n76106 , n76103 , n76104 );
xor ( n76107 , n74929 , n75376 );
nor ( n76108 , n51049 , n76024 );
and ( n76109 , n76107 , n76108 );
xor ( n76110 , n76107 , n76108 );
xor ( n76111 , n74933 , n75374 );
nor ( n76112 , n49850 , n76024 );
and ( n76113 , n76111 , n76112 );
xor ( n76114 , n76111 , n76112 );
xor ( n76115 , n74937 , n75372 );
nor ( n76116 , n48650 , n76024 );
and ( n76117 , n76115 , n76116 );
xor ( n76118 , n76115 , n76116 );
xor ( n76119 , n74941 , n75370 );
nor ( n76120 , n47449 , n76024 );
and ( n76121 , n76119 , n76120 );
xor ( n76122 , n76119 , n76120 );
xor ( n76123 , n74945 , n75368 );
nor ( n76124 , n46248 , n76024 );
and ( n76125 , n76123 , n76124 );
xor ( n76126 , n76123 , n76124 );
xor ( n76127 , n74949 , n75366 );
nor ( n76128 , n45047 , n76024 );
and ( n76129 , n76127 , n76128 );
xor ( n76130 , n76127 , n76128 );
xor ( n76131 , n74953 , n75364 );
nor ( n76132 , n43843 , n76024 );
and ( n76133 , n76131 , n76132 );
xor ( n76134 , n76131 , n76132 );
xor ( n76135 , n74957 , n75362 );
nor ( n76136 , n42641 , n76024 );
and ( n76137 , n76135 , n76136 );
xor ( n76138 , n76135 , n76136 );
xor ( n76139 , n74961 , n75360 );
nor ( n76140 , n41437 , n76024 );
and ( n76141 , n76139 , n76140 );
xor ( n76142 , n76139 , n76140 );
xor ( n76143 , n74965 , n75358 );
nor ( n76144 , n40232 , n76024 );
and ( n76145 , n76143 , n76144 );
xor ( n76146 , n76143 , n76144 );
xor ( n76147 , n74969 , n75356 );
nor ( n76148 , n39027 , n76024 );
and ( n76149 , n76147 , n76148 );
xor ( n76150 , n76147 , n76148 );
xor ( n76151 , n74973 , n75354 );
nor ( n76152 , n37825 , n76024 );
and ( n76153 , n76151 , n76152 );
xor ( n76154 , n76151 , n76152 );
xor ( n76155 , n74977 , n75352 );
nor ( n76156 , n36620 , n76024 );
and ( n76157 , n76155 , n76156 );
xor ( n76158 , n76155 , n76156 );
xor ( n76159 , n74981 , n75350 );
nor ( n76160 , n35419 , n76024 );
and ( n76161 , n76159 , n76160 );
xor ( n76162 , n76159 , n76160 );
xor ( n76163 , n74985 , n75348 );
nor ( n76164 , n34224 , n76024 );
and ( n76165 , n76163 , n76164 );
xor ( n76166 , n76163 , n76164 );
xor ( n76167 , n74989 , n75346 );
nor ( n76168 , n33033 , n76024 );
and ( n76169 , n76167 , n76168 );
xor ( n76170 , n76167 , n76168 );
xor ( n76171 , n74993 , n75344 );
nor ( n76172 , n31867 , n76024 );
and ( n76173 , n76171 , n76172 );
xor ( n76174 , n76171 , n76172 );
xor ( n76175 , n74997 , n75342 );
nor ( n76176 , n30725 , n76024 );
and ( n76177 , n76175 , n76176 );
xor ( n76178 , n76175 , n76176 );
xor ( n76179 , n75001 , n75340 );
nor ( n76180 , n29596 , n76024 );
and ( n76181 , n76179 , n76180 );
xor ( n76182 , n76179 , n76180 );
xor ( n76183 , n75005 , n75338 );
nor ( n76184 , n28487 , n76024 );
and ( n76185 , n76183 , n76184 );
xor ( n76186 , n76183 , n76184 );
xor ( n76187 , n75009 , n75336 );
nor ( n76188 , n27397 , n76024 );
and ( n76189 , n76187 , n76188 );
xor ( n76190 , n76187 , n76188 );
xor ( n76191 , n75013 , n75334 );
nor ( n76192 , n26326 , n76024 );
and ( n76193 , n76191 , n76192 );
xor ( n76194 , n76191 , n76192 );
xor ( n76195 , n75017 , n75332 );
nor ( n76196 , n25272 , n76024 );
and ( n76197 , n76195 , n76196 );
xor ( n76198 , n76195 , n76196 );
xor ( n76199 , n75021 , n75330 );
nor ( n76200 , n24242 , n76024 );
and ( n76201 , n76199 , n76200 );
xor ( n76202 , n76199 , n76200 );
xor ( n76203 , n75025 , n75328 );
nor ( n76204 , n23225 , n76024 );
and ( n76205 , n76203 , n76204 );
xor ( n76206 , n76203 , n76204 );
xor ( n76207 , n75029 , n75326 );
nor ( n76208 , n22231 , n76024 );
and ( n76209 , n76207 , n76208 );
xor ( n76210 , n76207 , n76208 );
xor ( n76211 , n75033 , n75324 );
nor ( n76212 , n21258 , n76024 );
and ( n76213 , n76211 , n76212 );
xor ( n76214 , n76211 , n76212 );
xor ( n76215 , n75037 , n75322 );
nor ( n76216 , n20303 , n76024 );
and ( n76217 , n76215 , n76216 );
xor ( n76218 , n76215 , n76216 );
xor ( n76219 , n75041 , n75320 );
nor ( n76220 , n19365 , n76024 );
and ( n76221 , n76219 , n76220 );
xor ( n76222 , n76219 , n76220 );
xor ( n76223 , n75045 , n75318 );
nor ( n76224 , n18448 , n76024 );
and ( n76225 , n76223 , n76224 );
xor ( n76226 , n76223 , n76224 );
xor ( n76227 , n75049 , n75316 );
nor ( n76228 , n17548 , n76024 );
and ( n76229 , n76227 , n76228 );
xor ( n76230 , n76227 , n76228 );
xor ( n76231 , n75053 , n75314 );
nor ( n76232 , n16669 , n76024 );
and ( n76233 , n76231 , n76232 );
xor ( n76234 , n76231 , n76232 );
xor ( n76235 , n75057 , n75312 );
nor ( n76236 , n15809 , n76024 );
and ( n76237 , n76235 , n76236 );
xor ( n76238 , n76235 , n76236 );
xor ( n76239 , n75061 , n75310 );
nor ( n76240 , n14968 , n76024 );
and ( n76241 , n76239 , n76240 );
xor ( n76242 , n76239 , n76240 );
xor ( n76243 , n75065 , n75308 );
nor ( n76244 , n14147 , n76024 );
and ( n76245 , n76243 , n76244 );
xor ( n76246 , n76243 , n76244 );
xor ( n76247 , n75069 , n75306 );
nor ( n76248 , n13349 , n76024 );
and ( n76249 , n76247 , n76248 );
xor ( n76250 , n76247 , n76248 );
xor ( n76251 , n75073 , n75304 );
nor ( n76252 , n12564 , n76024 );
and ( n76253 , n76251 , n76252 );
xor ( n76254 , n76251 , n76252 );
xor ( n76255 , n75077 , n75302 );
nor ( n76256 , n11799 , n76024 );
and ( n76257 , n76255 , n76256 );
xor ( n76258 , n76255 , n76256 );
xor ( n76259 , n75081 , n75300 );
nor ( n76260 , n11050 , n76024 );
and ( n76261 , n76259 , n76260 );
xor ( n76262 , n76259 , n76260 );
xor ( n76263 , n75085 , n75298 );
nor ( n76264 , n10321 , n76024 );
and ( n76265 , n76263 , n76264 );
xor ( n76266 , n76263 , n76264 );
xor ( n76267 , n75089 , n75296 );
nor ( n76268 , n9429 , n76024 );
and ( n76269 , n76267 , n76268 );
xor ( n76270 , n76267 , n76268 );
xor ( n76271 , n75093 , n75294 );
nor ( n76272 , n8949 , n76024 );
and ( n76273 , n76271 , n76272 );
xor ( n76274 , n76271 , n76272 );
xor ( n76275 , n75097 , n75292 );
nor ( n76276 , n9437 , n76024 );
and ( n76277 , n76275 , n76276 );
xor ( n76278 , n76275 , n76276 );
xor ( n76279 , n75101 , n75290 );
nor ( n76280 , n9446 , n76024 );
and ( n76281 , n76279 , n76280 );
xor ( n76282 , n76279 , n76280 );
xor ( n76283 , n75105 , n75288 );
nor ( n76284 , n9455 , n76024 );
and ( n76285 , n76283 , n76284 );
xor ( n76286 , n76283 , n76284 );
xor ( n76287 , n75109 , n75286 );
nor ( n76288 , n9464 , n76024 );
and ( n76289 , n76287 , n76288 );
xor ( n76290 , n76287 , n76288 );
xor ( n76291 , n75113 , n75284 );
nor ( n76292 , n9473 , n76024 );
and ( n76293 , n76291 , n76292 );
xor ( n76294 , n76291 , n76292 );
xor ( n76295 , n75117 , n75282 );
nor ( n76296 , n9482 , n76024 );
and ( n76297 , n76295 , n76296 );
xor ( n76298 , n76295 , n76296 );
xor ( n76299 , n75121 , n75280 );
nor ( n76300 , n9491 , n76024 );
and ( n76301 , n76299 , n76300 );
xor ( n76302 , n76299 , n76300 );
xor ( n76303 , n75125 , n75278 );
nor ( n76304 , n9500 , n76024 );
and ( n76305 , n76303 , n76304 );
xor ( n76306 , n76303 , n76304 );
xor ( n76307 , n75129 , n75276 );
nor ( n76308 , n9509 , n76024 );
and ( n76309 , n76307 , n76308 );
xor ( n76310 , n76307 , n76308 );
xor ( n76311 , n75133 , n75274 );
nor ( n76312 , n9518 , n76024 );
and ( n76313 , n76311 , n76312 );
xor ( n76314 , n76311 , n76312 );
xor ( n76315 , n75137 , n75272 );
nor ( n76316 , n9527 , n76024 );
and ( n76317 , n76315 , n76316 );
xor ( n76318 , n76315 , n76316 );
xor ( n76319 , n75141 , n75270 );
nor ( n76320 , n9536 , n76024 );
and ( n76321 , n76319 , n76320 );
xor ( n76322 , n76319 , n76320 );
xor ( n76323 , n75145 , n75268 );
nor ( n76324 , n9545 , n76024 );
and ( n76325 , n76323 , n76324 );
xor ( n76326 , n76323 , n76324 );
xor ( n76327 , n75149 , n75266 );
nor ( n76328 , n9554 , n76024 );
and ( n76329 , n76327 , n76328 );
xor ( n76330 , n76327 , n76328 );
xor ( n76331 , n75153 , n75264 );
nor ( n76332 , n9563 , n76024 );
and ( n76333 , n76331 , n76332 );
xor ( n76334 , n76331 , n76332 );
xor ( n76335 , n75157 , n75262 );
nor ( n76336 , n9572 , n76024 );
and ( n76337 , n76335 , n76336 );
xor ( n76338 , n76335 , n76336 );
xor ( n76339 , n75161 , n75260 );
nor ( n76340 , n9581 , n76024 );
and ( n76341 , n76339 , n76340 );
xor ( n76342 , n76339 , n76340 );
xor ( n76343 , n75165 , n75258 );
nor ( n76344 , n9590 , n76024 );
and ( n76345 , n76343 , n76344 );
xor ( n76346 , n76343 , n76344 );
xor ( n76347 , n75169 , n75256 );
nor ( n76348 , n9599 , n76024 );
and ( n76349 , n76347 , n76348 );
xor ( n76350 , n76347 , n76348 );
xor ( n76351 , n75173 , n75254 );
nor ( n76352 , n9608 , n76024 );
and ( n76353 , n76351 , n76352 );
xor ( n76354 , n76351 , n76352 );
xor ( n76355 , n75177 , n75252 );
nor ( n76356 , n9617 , n76024 );
and ( n76357 , n76355 , n76356 );
xor ( n76358 , n76355 , n76356 );
xor ( n76359 , n75181 , n75250 );
nor ( n76360 , n9626 , n76024 );
and ( n76361 , n76359 , n76360 );
xor ( n76362 , n76359 , n76360 );
xor ( n76363 , n75185 , n75248 );
nor ( n76364 , n9635 , n76024 );
and ( n76365 , n76363 , n76364 );
xor ( n76366 , n76363 , n76364 );
xor ( n76367 , n75189 , n75246 );
nor ( n76368 , n9644 , n76024 );
and ( n76369 , n76367 , n76368 );
xor ( n76370 , n76367 , n76368 );
xor ( n76371 , n75193 , n75244 );
nor ( n76372 , n9653 , n76024 );
and ( n76373 , n76371 , n76372 );
xor ( n76374 , n76371 , n76372 );
xor ( n76375 , n75197 , n75242 );
nor ( n76376 , n9662 , n76024 );
and ( n76377 , n76375 , n76376 );
xor ( n76378 , n76375 , n76376 );
xor ( n76379 , n75201 , n75240 );
nor ( n76380 , n9671 , n76024 );
and ( n76381 , n76379 , n76380 );
xor ( n76382 , n76379 , n76380 );
xor ( n76383 , n75205 , n75238 );
nor ( n76384 , n9680 , n76024 );
and ( n76385 , n76383 , n76384 );
xor ( n76386 , n76383 , n76384 );
xor ( n76387 , n75209 , n75236 );
nor ( n76388 , n9689 , n76024 );
and ( n76389 , n76387 , n76388 );
xor ( n76390 , n76387 , n76388 );
xor ( n76391 , n75213 , n75234 );
nor ( n76392 , n9698 , n76024 );
and ( n76393 , n76391 , n76392 );
xor ( n76394 , n76391 , n76392 );
xor ( n76395 , n75217 , n75232 );
nor ( n76396 , n9707 , n76024 );
and ( n76397 , n76395 , n76396 );
xor ( n76398 , n76395 , n76396 );
xor ( n76399 , n75221 , n75230 );
nor ( n76400 , n9716 , n76024 );
and ( n76401 , n76399 , n76400 );
xor ( n76402 , n76399 , n76400 );
xor ( n76403 , n75225 , n75228 );
nor ( n76404 , n9725 , n76024 );
and ( n76405 , n76403 , n76404 );
xor ( n76406 , n76403 , n76404 );
xor ( n76407 , n75226 , n75227 );
nor ( n76408 , n9734 , n76024 );
and ( n76409 , n76407 , n76408 );
xor ( n76410 , n76407 , n76408 );
nor ( n76411 , n9752 , n74843 );
nor ( n76412 , n9743 , n76024 );
and ( n76413 , n76411 , n76412 );
and ( n76414 , n76410 , n76413 );
or ( n76415 , n76409 , n76414 );
and ( n76416 , n76406 , n76415 );
or ( n76417 , n76405 , n76416 );
and ( n76418 , n76402 , n76417 );
or ( n76419 , n76401 , n76418 );
and ( n76420 , n76398 , n76419 );
or ( n76421 , n76397 , n76420 );
and ( n76422 , n76394 , n76421 );
or ( n76423 , n76393 , n76422 );
and ( n76424 , n76390 , n76423 );
or ( n76425 , n76389 , n76424 );
and ( n76426 , n76386 , n76425 );
or ( n76427 , n76385 , n76426 );
and ( n76428 , n76382 , n76427 );
or ( n76429 , n76381 , n76428 );
and ( n76430 , n76378 , n76429 );
or ( n76431 , n76377 , n76430 );
and ( n76432 , n76374 , n76431 );
or ( n76433 , n76373 , n76432 );
and ( n76434 , n76370 , n76433 );
or ( n76435 , n76369 , n76434 );
and ( n76436 , n76366 , n76435 );
or ( n76437 , n76365 , n76436 );
and ( n76438 , n76362 , n76437 );
or ( n76439 , n76361 , n76438 );
and ( n76440 , n76358 , n76439 );
or ( n76441 , n76357 , n76440 );
and ( n76442 , n76354 , n76441 );
or ( n76443 , n76353 , n76442 );
and ( n76444 , n76350 , n76443 );
or ( n76445 , n76349 , n76444 );
and ( n76446 , n76346 , n76445 );
or ( n76447 , n76345 , n76446 );
and ( n76448 , n76342 , n76447 );
or ( n76449 , n76341 , n76448 );
and ( n76450 , n76338 , n76449 );
or ( n76451 , n76337 , n76450 );
and ( n76452 , n76334 , n76451 );
or ( n76453 , n76333 , n76452 );
and ( n76454 , n76330 , n76453 );
or ( n76455 , n76329 , n76454 );
and ( n76456 , n76326 , n76455 );
or ( n76457 , n76325 , n76456 );
and ( n76458 , n76322 , n76457 );
or ( n76459 , n76321 , n76458 );
and ( n76460 , n76318 , n76459 );
or ( n76461 , n76317 , n76460 );
and ( n76462 , n76314 , n76461 );
or ( n76463 , n76313 , n76462 );
and ( n76464 , n76310 , n76463 );
or ( n76465 , n76309 , n76464 );
and ( n76466 , n76306 , n76465 );
or ( n76467 , n76305 , n76466 );
and ( n76468 , n76302 , n76467 );
or ( n76469 , n76301 , n76468 );
and ( n76470 , n76298 , n76469 );
or ( n76471 , n76297 , n76470 );
and ( n76472 , n76294 , n76471 );
or ( n76473 , n76293 , n76472 );
and ( n76474 , n76290 , n76473 );
or ( n76475 , n76289 , n76474 );
and ( n76476 , n76286 , n76475 );
or ( n76477 , n76285 , n76476 );
and ( n76478 , n76282 , n76477 );
or ( n76479 , n76281 , n76478 );
and ( n76480 , n76278 , n76479 );
or ( n76481 , n76277 , n76480 );
and ( n76482 , n76274 , n76481 );
or ( n76483 , n76273 , n76482 );
and ( n76484 , n76270 , n76483 );
or ( n76485 , n76269 , n76484 );
and ( n76486 , n76266 , n76485 );
or ( n76487 , n76265 , n76486 );
and ( n76488 , n76262 , n76487 );
or ( n76489 , n76261 , n76488 );
and ( n76490 , n76258 , n76489 );
or ( n76491 , n76257 , n76490 );
and ( n76492 , n76254 , n76491 );
or ( n76493 , n76253 , n76492 );
and ( n76494 , n76250 , n76493 );
or ( n76495 , n76249 , n76494 );
and ( n76496 , n76246 , n76495 );
or ( n76497 , n76245 , n76496 );
and ( n76498 , n76242 , n76497 );
or ( n76499 , n76241 , n76498 );
and ( n76500 , n76238 , n76499 );
or ( n76501 , n76237 , n76500 );
and ( n76502 , n76234 , n76501 );
or ( n76503 , n76233 , n76502 );
and ( n76504 , n76230 , n76503 );
or ( n76505 , n76229 , n76504 );
and ( n76506 , n76226 , n76505 );
or ( n76507 , n76225 , n76506 );
and ( n76508 , n76222 , n76507 );
or ( n76509 , n76221 , n76508 );
and ( n76510 , n76218 , n76509 );
or ( n76511 , n76217 , n76510 );
and ( n76512 , n76214 , n76511 );
or ( n76513 , n76213 , n76512 );
and ( n76514 , n76210 , n76513 );
or ( n76515 , n76209 , n76514 );
and ( n76516 , n76206 , n76515 );
or ( n76517 , n76205 , n76516 );
and ( n76518 , n76202 , n76517 );
or ( n76519 , n76201 , n76518 );
and ( n76520 , n76198 , n76519 );
or ( n76521 , n76197 , n76520 );
and ( n76522 , n76194 , n76521 );
or ( n76523 , n76193 , n76522 );
and ( n76524 , n76190 , n76523 );
or ( n76525 , n76189 , n76524 );
and ( n76526 , n76186 , n76525 );
or ( n76527 , n76185 , n76526 );
and ( n76528 , n76182 , n76527 );
or ( n76529 , n76181 , n76528 );
and ( n76530 , n76178 , n76529 );
or ( n76531 , n76177 , n76530 );
and ( n76532 , n76174 , n76531 );
or ( n76533 , n76173 , n76532 );
and ( n76534 , n76170 , n76533 );
or ( n76535 , n76169 , n76534 );
and ( n76536 , n76166 , n76535 );
or ( n76537 , n76165 , n76536 );
and ( n76538 , n76162 , n76537 );
or ( n76539 , n76161 , n76538 );
and ( n76540 , n76158 , n76539 );
or ( n76541 , n76157 , n76540 );
and ( n76542 , n76154 , n76541 );
or ( n76543 , n76153 , n76542 );
and ( n76544 , n76150 , n76543 );
or ( n76545 , n76149 , n76544 );
and ( n76546 , n76146 , n76545 );
or ( n76547 , n76145 , n76546 );
and ( n76548 , n76142 , n76547 );
or ( n76549 , n76141 , n76548 );
and ( n76550 , n76138 , n76549 );
or ( n76551 , n76137 , n76550 );
and ( n76552 , n76134 , n76551 );
or ( n76553 , n76133 , n76552 );
and ( n76554 , n76130 , n76553 );
or ( n76555 , n76129 , n76554 );
and ( n76556 , n76126 , n76555 );
or ( n76557 , n76125 , n76556 );
and ( n76558 , n76122 , n76557 );
or ( n76559 , n76121 , n76558 );
and ( n76560 , n76118 , n76559 );
or ( n76561 , n76117 , n76560 );
and ( n76562 , n76114 , n76561 );
or ( n76563 , n76113 , n76562 );
and ( n76564 , n76110 , n76563 );
or ( n76565 , n76109 , n76564 );
and ( n76566 , n76106 , n76565 );
or ( n76567 , n76105 , n76566 );
and ( n76568 , n76102 , n76567 );
or ( n76569 , n76101 , n76568 );
and ( n76570 , n76098 , n76569 );
or ( n76571 , n76097 , n76570 );
and ( n76572 , n76094 , n76571 );
or ( n76573 , n76093 , n76572 );
and ( n76574 , n76090 , n76573 );
or ( n76575 , n76089 , n76574 );
and ( n76576 , n76086 , n76575 );
or ( n76577 , n76085 , n76576 );
and ( n76578 , n76082 , n76577 );
or ( n76579 , n76081 , n76578 );
and ( n76580 , n76078 , n76579 );
or ( n76581 , n76077 , n76580 );
and ( n76582 , n76074 , n76581 );
or ( n76583 , n76073 , n76582 );
and ( n76584 , n76070 , n76583 );
or ( n76585 , n76069 , n76584 );
and ( n76586 , n76066 , n76585 );
or ( n76587 , n76065 , n76586 );
and ( n76588 , n76062 , n76587 );
or ( n76589 , n76061 , n76588 );
and ( n76590 , n76058 , n76589 );
or ( n76591 , n76057 , n76590 );
and ( n76592 , n76054 , n76591 );
or ( n76593 , n76053 , n76592 );
and ( n76594 , n76050 , n76593 );
or ( n76595 , n76049 , n76594 );
and ( n76596 , n76046 , n76595 );
or ( n76597 , n76045 , n76596 );
and ( n76598 , n76042 , n76597 );
or ( n76599 , n76041 , n76598 );
and ( n76600 , n76038 , n76599 );
or ( n76601 , n76037 , n76600 );
and ( n76602 , n76034 , n76601 );
or ( n76603 , n76033 , n76602 );
and ( n76604 , n76030 , n76603 );
or ( n76605 , n76029 , n76604 );
xor ( n76606 , n76026 , n76605 );
and ( n76607 , n33403 , n8736 );
nor ( n76608 , n8737 , n76607 );
nor ( n76609 , n9420 , n32231 );
xor ( n76610 , n76608 , n76609 );
and ( n76611 , n75421 , n75422 );
and ( n76612 , n75423 , n75426 );
or ( n76613 , n76611 , n76612 );
xor ( n76614 , n76610 , n76613 );
nor ( n76615 , n10312 , n31083 );
xor ( n76616 , n76614 , n76615 );
and ( n76617 , n75427 , n75428 );
and ( n76618 , n75429 , n75432 );
or ( n76619 , n76617 , n76618 );
xor ( n76620 , n76616 , n76619 );
nor ( n76621 , n11041 , n29948 );
xor ( n76622 , n76620 , n76621 );
and ( n76623 , n75433 , n75434 );
and ( n76624 , n75435 , n75438 );
or ( n76625 , n76623 , n76624 );
xor ( n76626 , n76622 , n76625 );
nor ( n76627 , n11790 , n28833 );
xor ( n76628 , n76626 , n76627 );
and ( n76629 , n75439 , n75440 );
and ( n76630 , n75441 , n75444 );
or ( n76631 , n76629 , n76630 );
xor ( n76632 , n76628 , n76631 );
nor ( n76633 , n12555 , n27737 );
xor ( n76634 , n76632 , n76633 );
and ( n76635 , n75445 , n75446 );
and ( n76636 , n75447 , n75450 );
or ( n76637 , n76635 , n76636 );
xor ( n76638 , n76634 , n76637 );
nor ( n76639 , n13340 , n26660 );
xor ( n76640 , n76638 , n76639 );
and ( n76641 , n75451 , n75452 );
and ( n76642 , n75453 , n75456 );
or ( n76643 , n76641 , n76642 );
xor ( n76644 , n76640 , n76643 );
nor ( n76645 , n14138 , n25600 );
xor ( n76646 , n76644 , n76645 );
and ( n76647 , n75457 , n75458 );
and ( n76648 , n75459 , n75462 );
or ( n76649 , n76647 , n76648 );
xor ( n76650 , n76646 , n76649 );
nor ( n76651 , n14959 , n24564 );
xor ( n76652 , n76650 , n76651 );
and ( n76653 , n75463 , n75464 );
and ( n76654 , n75465 , n75468 );
or ( n76655 , n76653 , n76654 );
xor ( n76656 , n76652 , n76655 );
nor ( n76657 , n15800 , n23541 );
xor ( n76658 , n76656 , n76657 );
and ( n76659 , n75469 , n75470 );
and ( n76660 , n75471 , n75474 );
or ( n76661 , n76659 , n76660 );
xor ( n76662 , n76658 , n76661 );
nor ( n76663 , n16660 , n22541 );
xor ( n76664 , n76662 , n76663 );
and ( n76665 , n75475 , n75476 );
and ( n76666 , n75477 , n75480 );
or ( n76667 , n76665 , n76666 );
xor ( n76668 , n76664 , n76667 );
nor ( n76669 , n17539 , n21562 );
xor ( n76670 , n76668 , n76669 );
and ( n76671 , n75481 , n75482 );
and ( n76672 , n75483 , n75486 );
or ( n76673 , n76671 , n76672 );
xor ( n76674 , n76670 , n76673 );
nor ( n76675 , n18439 , n20601 );
xor ( n76676 , n76674 , n76675 );
and ( n76677 , n75487 , n75488 );
and ( n76678 , n75489 , n75492 );
or ( n76679 , n76677 , n76678 );
xor ( n76680 , n76676 , n76679 );
nor ( n76681 , n19356 , n19657 );
xor ( n76682 , n76680 , n76681 );
and ( n76683 , n75493 , n75494 );
and ( n76684 , n75495 , n75498 );
or ( n76685 , n76683 , n76684 );
xor ( n76686 , n76682 , n76685 );
nor ( n76687 , n20294 , n18734 );
xor ( n76688 , n76686 , n76687 );
and ( n76689 , n75499 , n75500 );
and ( n76690 , n75501 , n75504 );
or ( n76691 , n76689 , n76690 );
xor ( n76692 , n76688 , n76691 );
nor ( n76693 , n21249 , n17828 );
xor ( n76694 , n76692 , n76693 );
and ( n76695 , n75505 , n75506 );
and ( n76696 , n75507 , n75510 );
or ( n76697 , n76695 , n76696 );
xor ( n76698 , n76694 , n76697 );
nor ( n76699 , n22222 , n16943 );
xor ( n76700 , n76698 , n76699 );
and ( n76701 , n75511 , n75512 );
and ( n76702 , n75513 , n75516 );
or ( n76703 , n76701 , n76702 );
xor ( n76704 , n76700 , n76703 );
nor ( n76705 , n23216 , n16077 );
xor ( n76706 , n76704 , n76705 );
and ( n76707 , n75517 , n75518 );
and ( n76708 , n75519 , n75522 );
or ( n76709 , n76707 , n76708 );
xor ( n76710 , n76706 , n76709 );
nor ( n76711 , n24233 , n15230 );
xor ( n76712 , n76710 , n76711 );
and ( n76713 , n75523 , n75524 );
and ( n76714 , n75525 , n75528 );
or ( n76715 , n76713 , n76714 );
xor ( n76716 , n76712 , n76715 );
nor ( n76717 , n25263 , n14403 );
xor ( n76718 , n76716 , n76717 );
and ( n76719 , n75529 , n75530 );
and ( n76720 , n75531 , n75534 );
or ( n76721 , n76719 , n76720 );
xor ( n76722 , n76718 , n76721 );
nor ( n76723 , n26317 , n13599 );
xor ( n76724 , n76722 , n76723 );
and ( n76725 , n75535 , n75536 );
and ( n76726 , n75537 , n75540 );
or ( n76727 , n76725 , n76726 );
xor ( n76728 , n76724 , n76727 );
nor ( n76729 , n27388 , n12808 );
xor ( n76730 , n76728 , n76729 );
and ( n76731 , n75541 , n75542 );
and ( n76732 , n75543 , n75546 );
or ( n76733 , n76731 , n76732 );
xor ( n76734 , n76730 , n76733 );
nor ( n76735 , n28478 , n12037 );
xor ( n76736 , n76734 , n76735 );
and ( n76737 , n75547 , n75548 );
and ( n76738 , n75549 , n75552 );
or ( n76739 , n76737 , n76738 );
xor ( n76740 , n76736 , n76739 );
nor ( n76741 , n29587 , n11282 );
xor ( n76742 , n76740 , n76741 );
and ( n76743 , n75553 , n75554 );
and ( n76744 , n75555 , n75558 );
or ( n76745 , n76743 , n76744 );
xor ( n76746 , n76742 , n76745 );
nor ( n76747 , n30716 , n10547 );
xor ( n76748 , n76746 , n76747 );
and ( n76749 , n75559 , n75560 );
and ( n76750 , n75561 , n75564 );
or ( n76751 , n76749 , n76750 );
xor ( n76752 , n76748 , n76751 );
nor ( n76753 , n31858 , n9829 );
xor ( n76754 , n76752 , n76753 );
and ( n76755 , n75565 , n75566 );
and ( n76756 , n75567 , n75570 );
or ( n76757 , n76755 , n76756 );
xor ( n76758 , n76754 , n76757 );
nor ( n76759 , n33024 , n8955 );
xor ( n76760 , n76758 , n76759 );
and ( n76761 , n75571 , n75572 );
and ( n76762 , n75573 , n75576 );
or ( n76763 , n76761 , n76762 );
xor ( n76764 , n76760 , n76763 );
nor ( n76765 , n34215 , n603 );
xor ( n76766 , n76764 , n76765 );
and ( n76767 , n75577 , n75578 );
and ( n76768 , n75579 , n75582 );
or ( n76769 , n76767 , n76768 );
xor ( n76770 , n76766 , n76769 );
nor ( n76771 , n35410 , n652 );
xor ( n76772 , n76770 , n76771 );
and ( n76773 , n75583 , n75584 );
and ( n76774 , n75585 , n75588 );
or ( n76775 , n76773 , n76774 );
xor ( n76776 , n76772 , n76775 );
nor ( n76777 , n36611 , n624 );
xor ( n76778 , n76776 , n76777 );
and ( n76779 , n75589 , n75590 );
and ( n76780 , n75591 , n75594 );
or ( n76781 , n76779 , n76780 );
xor ( n76782 , n76778 , n76781 );
nor ( n76783 , n37816 , n648 );
xor ( n76784 , n76782 , n76783 );
and ( n76785 , n75595 , n75596 );
and ( n76786 , n75597 , n75600 );
or ( n76787 , n76785 , n76786 );
xor ( n76788 , n76784 , n76787 );
nor ( n76789 , n39018 , n686 );
xor ( n76790 , n76788 , n76789 );
and ( n76791 , n75601 , n75602 );
and ( n76792 , n75603 , n75606 );
or ( n76793 , n76791 , n76792 );
xor ( n76794 , n76790 , n76793 );
nor ( n76795 , n40223 , n735 );
xor ( n76796 , n76794 , n76795 );
and ( n76797 , n75607 , n75608 );
and ( n76798 , n75609 , n75612 );
or ( n76799 , n76797 , n76798 );
xor ( n76800 , n76796 , n76799 );
nor ( n76801 , n41428 , n798 );
xor ( n76802 , n76800 , n76801 );
and ( n76803 , n75613 , n75614 );
and ( n76804 , n75615 , n75618 );
or ( n76805 , n76803 , n76804 );
xor ( n76806 , n76802 , n76805 );
nor ( n76807 , n42632 , n870 );
xor ( n76808 , n76806 , n76807 );
and ( n76809 , n75619 , n75620 );
and ( n76810 , n75621 , n75624 );
or ( n76811 , n76809 , n76810 );
xor ( n76812 , n76808 , n76811 );
nor ( n76813 , n43834 , n960 );
xor ( n76814 , n76812 , n76813 );
and ( n76815 , n75625 , n75626 );
and ( n76816 , n75627 , n75630 );
or ( n76817 , n76815 , n76816 );
xor ( n76818 , n76814 , n76817 );
nor ( n76819 , n45038 , n1064 );
xor ( n76820 , n76818 , n76819 );
and ( n76821 , n75631 , n75632 );
and ( n76822 , n75633 , n75636 );
or ( n76823 , n76821 , n76822 );
xor ( n76824 , n76820 , n76823 );
nor ( n76825 , n46239 , n1178 );
xor ( n76826 , n76824 , n76825 );
and ( n76827 , n75637 , n75638 );
and ( n76828 , n75639 , n75642 );
or ( n76829 , n76827 , n76828 );
xor ( n76830 , n76826 , n76829 );
nor ( n76831 , n47440 , n1305 );
xor ( n76832 , n76830 , n76831 );
and ( n76833 , n75643 , n75644 );
and ( n76834 , n75645 , n75648 );
or ( n76835 , n76833 , n76834 );
xor ( n76836 , n76832 , n76835 );
nor ( n76837 , n48641 , n1447 );
xor ( n76838 , n76836 , n76837 );
and ( n76839 , n75649 , n75650 );
and ( n76840 , n75651 , n75654 );
or ( n76841 , n76839 , n76840 );
xor ( n76842 , n76838 , n76841 );
nor ( n76843 , n49841 , n1600 );
xor ( n76844 , n76842 , n76843 );
and ( n76845 , n75655 , n75656 );
and ( n76846 , n75657 , n75660 );
or ( n76847 , n76845 , n76846 );
xor ( n76848 , n76844 , n76847 );
nor ( n76849 , n51040 , n1768 );
xor ( n76850 , n76848 , n76849 );
and ( n76851 , n75661 , n75662 );
and ( n76852 , n75663 , n75666 );
or ( n76853 , n76851 , n76852 );
xor ( n76854 , n76850 , n76853 );
nor ( n76855 , n52238 , n1947 );
xor ( n76856 , n76854 , n76855 );
and ( n76857 , n75667 , n75668 );
and ( n76858 , n75669 , n75672 );
or ( n76859 , n76857 , n76858 );
xor ( n76860 , n76856 , n76859 );
nor ( n76861 , n53432 , n2139 );
xor ( n76862 , n76860 , n76861 );
and ( n76863 , n75673 , n75674 );
and ( n76864 , n75675 , n75678 );
or ( n76865 , n76863 , n76864 );
xor ( n76866 , n76862 , n76865 );
nor ( n76867 , n54629 , n2345 );
xor ( n76868 , n76866 , n76867 );
and ( n76869 , n75679 , n75680 );
and ( n76870 , n75681 , n75684 );
or ( n76871 , n76869 , n76870 );
xor ( n76872 , n76868 , n76871 );
nor ( n76873 , n55826 , n2568 );
xor ( n76874 , n76872 , n76873 );
and ( n76875 , n75685 , n75686 );
and ( n76876 , n75687 , n75690 );
or ( n76877 , n76875 , n76876 );
xor ( n76878 , n76874 , n76877 );
nor ( n76879 , n57022 , n2799 );
xor ( n76880 , n76878 , n76879 );
and ( n76881 , n75691 , n75692 );
and ( n76882 , n75693 , n75696 );
or ( n76883 , n76881 , n76882 );
xor ( n76884 , n76880 , n76883 );
nor ( n76885 , n58217 , n3045 );
xor ( n76886 , n76884 , n76885 );
and ( n76887 , n75697 , n75698 );
and ( n76888 , n75699 , n75702 );
or ( n76889 , n76887 , n76888 );
xor ( n76890 , n76886 , n76889 );
nor ( n76891 , n59412 , n3302 );
xor ( n76892 , n76890 , n76891 );
and ( n76893 , n75703 , n75704 );
and ( n76894 , n75705 , n75708 );
or ( n76895 , n76893 , n76894 );
xor ( n76896 , n76892 , n76895 );
nor ( n76897 , n60600 , n3572 );
xor ( n76898 , n76896 , n76897 );
and ( n76899 , n75709 , n75710 );
and ( n76900 , n75711 , n75714 );
or ( n76901 , n76899 , n76900 );
xor ( n76902 , n76898 , n76901 );
nor ( n76903 , n61791 , n3855 );
xor ( n76904 , n76902 , n76903 );
and ( n76905 , n75715 , n75716 );
and ( n76906 , n75717 , n75720 );
or ( n76907 , n76905 , n76906 );
xor ( n76908 , n76904 , n76907 );
nor ( n76909 , n62982 , n4153 );
xor ( n76910 , n76908 , n76909 );
and ( n76911 , n75721 , n75722 );
and ( n76912 , n75723 , n75726 );
or ( n76913 , n76911 , n76912 );
xor ( n76914 , n76910 , n76913 );
nor ( n76915 , n64172 , n4460 );
xor ( n76916 , n76914 , n76915 );
and ( n76917 , n75727 , n75728 );
and ( n76918 , n75729 , n75732 );
or ( n76919 , n76917 , n76918 );
xor ( n76920 , n76916 , n76919 );
nor ( n76921 , n65360 , n4788 );
xor ( n76922 , n76920 , n76921 );
and ( n76923 , n75733 , n75734 );
and ( n76924 , n75735 , n75738 );
or ( n76925 , n76923 , n76924 );
xor ( n76926 , n76922 , n76925 );
nor ( n76927 , n66550 , n5128 );
xor ( n76928 , n76926 , n76927 );
and ( n76929 , n75739 , n75740 );
and ( n76930 , n75741 , n75744 );
or ( n76931 , n76929 , n76930 );
xor ( n76932 , n76928 , n76931 );
nor ( n76933 , n67736 , n5479 );
xor ( n76934 , n76932 , n76933 );
and ( n76935 , n75745 , n75746 );
and ( n76936 , n75747 , n75750 );
or ( n76937 , n76935 , n76936 );
xor ( n76938 , n76934 , n76937 );
nor ( n76939 , n68924 , n5840 );
xor ( n76940 , n76938 , n76939 );
and ( n76941 , n75751 , n75752 );
and ( n76942 , n75753 , n75756 );
or ( n76943 , n76941 , n76942 );
xor ( n76944 , n76940 , n76943 );
nor ( n76945 , n70110 , n6214 );
xor ( n76946 , n76944 , n76945 );
and ( n76947 , n75757 , n75758 );
and ( n76948 , n75759 , n75762 );
or ( n76949 , n76947 , n76948 );
xor ( n76950 , n76946 , n76949 );
nor ( n76951 , n71292 , n6598 );
xor ( n76952 , n76950 , n76951 );
and ( n76953 , n75763 , n75764 );
and ( n76954 , n75765 , n75768 );
or ( n76955 , n76953 , n76954 );
xor ( n76956 , n76952 , n76955 );
nor ( n76957 , n72472 , n6999 );
xor ( n76958 , n76956 , n76957 );
and ( n76959 , n75769 , n75770 );
and ( n76960 , n75771 , n75774 );
or ( n76961 , n76959 , n76960 );
xor ( n76962 , n76958 , n76961 );
nor ( n76963 , n73654 , n7415 );
xor ( n76964 , n76962 , n76963 );
and ( n76965 , n75775 , n75776 );
and ( n76966 , n75777 , n75780 );
or ( n76967 , n76965 , n76966 );
xor ( n76968 , n76964 , n76967 );
nor ( n76969 , n74832 , n7843 );
xor ( n76970 , n76968 , n76969 );
and ( n76971 , n75781 , n75782 );
and ( n76972 , n75783 , n75786 );
or ( n76973 , n76971 , n76972 );
xor ( n76974 , n76970 , n76973 );
nor ( n76975 , n76013 , n8283 );
xor ( n76976 , n76974 , n76975 );
and ( n76977 , n75787 , n75788 );
and ( n76978 , n75789 , n75792 );
or ( n76979 , n76977 , n76978 );
xor ( n76980 , n76976 , n76979 );
and ( n76981 , n75805 , n75809 );
and ( n76982 , n75809 , n75999 );
and ( n76983 , n75805 , n75999 );
or ( n76984 , n76981 , n76982 , n76983 );
and ( n76985 , n33774 , n8669 );
not ( n76986 , n8669 );
nor ( n76987 , n76985 , n76986 );
xor ( n76988 , n76984 , n76987 );
and ( n76989 , n75815 , n75816 );
and ( n76990 , n75816 , n75884 );
and ( n76991 , n75815 , n75884 );
or ( n76992 , n76989 , n76990 , n76991 );
and ( n76993 , n75811 , n75885 );
and ( n76994 , n75885 , n75998 );
and ( n76995 , n75811 , n75998 );
or ( n76996 , n76993 , n76994 , n76995 );
xor ( n76997 , n76992 , n76996 );
and ( n76998 , n75891 , n75997 );
and ( n76999 , n75821 , n75825 );
and ( n77000 , n75825 , n75883 );
and ( n77001 , n75821 , n75883 );
or ( n77002 , n76999 , n77000 , n77001 );
and ( n77003 , n75895 , n75996 );
xor ( n77004 , n77002 , n77003 );
and ( n77005 , n75852 , n75856 );
and ( n77006 , n75856 , n75862 );
and ( n77007 , n75852 , n75862 );
or ( n77008 , n77005 , n77006 , n77007 );
and ( n77009 , n75830 , n75834 );
and ( n77010 , n75834 , n75882 );
and ( n77011 , n75830 , n75882 );
or ( n77012 , n77009 , n77010 , n77011 );
xor ( n77013 , n77008 , n77012 );
and ( n77014 , n75839 , n75843 );
and ( n77015 , n75843 , n75881 );
and ( n77016 , n75839 , n75881 );
or ( n77017 , n77014 , n77015 , n77016 );
and ( n77018 , n75900 , n75927 );
and ( n77019 , n75927 , n75965 );
and ( n77020 , n75900 , n75965 );
or ( n77021 , n77018 , n77019 , n77020 );
xor ( n77022 , n77017 , n77021 );
and ( n77023 , n75848 , n75863 );
and ( n77024 , n75863 , n75880 );
and ( n77025 , n75848 , n75880 );
or ( n77026 , n77023 , n77024 , n77025 );
and ( n77027 , n75904 , n75908 );
and ( n77028 , n75908 , n75926 );
and ( n77029 , n75904 , n75926 );
or ( n77030 , n77027 , n77028 , n77029 );
xor ( n77031 , n77026 , n77030 );
and ( n77032 , n75868 , n75873 );
and ( n77033 , n75873 , n75879 );
and ( n77034 , n75868 , n75879 );
or ( n77035 , n77032 , n77033 , n77034 );
and ( n77036 , n75858 , n75859 );
and ( n77037 , n75859 , n75861 );
and ( n77038 , n75858 , n75861 );
or ( n77039 , n77036 , n77037 , n77038 );
and ( n77040 , n75869 , n75870 );
and ( n77041 , n75870 , n75872 );
and ( n77042 , n75869 , n75872 );
or ( n77043 , n77040 , n77041 , n77042 );
xor ( n77044 , n77039 , n77043 );
and ( n77045 , n30695 , n10977 );
and ( n77046 , n31836 , n10239 );
xor ( n77047 , n77045 , n77046 );
and ( n77048 , n32649 , n9348 );
xor ( n77049 , n77047 , n77048 );
xor ( n77050 , n77044 , n77049 );
xor ( n77051 , n77035 , n77050 );
and ( n77052 , n75875 , n75876 );
and ( n77053 , n75876 , n75878 );
and ( n77054 , n75875 , n75878 );
or ( n77055 , n77052 , n77053 , n77054 );
and ( n77056 , n27361 , n13256 );
and ( n77057 , n28456 , n12531 );
xor ( n77058 , n77056 , n77057 );
and ( n77059 , n29559 , n11718 );
xor ( n77060 , n77058 , n77059 );
xor ( n77061 , n77055 , n77060 );
and ( n77062 , n24214 , n15691 );
and ( n77063 , n25243 , n14838 );
xor ( n77064 , n77062 , n77063 );
and ( n77065 , n26296 , n14044 );
xor ( n77066 , n77064 , n77065 );
xor ( n77067 , n77061 , n77066 );
xor ( n77068 , n77051 , n77067 );
xor ( n77069 , n77031 , n77068 );
xor ( n77070 , n77022 , n77069 );
xor ( n77071 , n77013 , n77070 );
xor ( n77072 , n77004 , n77071 );
xor ( n77073 , n76998 , n77072 );
and ( n77074 , n75896 , n75966 );
and ( n77075 , n75966 , n75995 );
and ( n77076 , n75896 , n75995 );
or ( n77077 , n77074 , n77075 , n77076 );
and ( n77078 , n75971 , n75994 );
and ( n77079 , n75932 , n75948 );
and ( n77080 , n75948 , n75964 );
and ( n77081 , n75932 , n75964 );
or ( n77082 , n77079 , n77080 , n77081 );
and ( n77083 , n75913 , n75919 );
and ( n77084 , n75919 , n75925 );
and ( n77085 , n75913 , n75925 );
or ( n77086 , n77083 , n77084 , n77085 );
and ( n77087 , n75936 , n75941 );
and ( n77088 , n75941 , n75947 );
and ( n77089 , n75936 , n75947 );
or ( n77090 , n77087 , n77088 , n77089 );
xor ( n77091 , n77086 , n77090 );
and ( n77092 , n75921 , n75922 );
and ( n77093 , n75922 , n75924 );
and ( n77094 , n75921 , n75924 );
or ( n77095 , n77092 , n77093 , n77094 );
and ( n77096 , n75937 , n75938 );
and ( n77097 , n75938 , n75940 );
and ( n77098 , n75937 , n75940 );
or ( n77099 , n77096 , n77097 , n77098 );
xor ( n77100 , n77095 , n77099 );
and ( n77101 , n21216 , n18407 );
and ( n77102 , n22186 , n17422 );
xor ( n77103 , n77101 , n77102 );
and ( n77104 , n22892 , n16550 );
xor ( n77105 , n77103 , n77104 );
xor ( n77106 , n77100 , n77105 );
xor ( n77107 , n77091 , n77106 );
xor ( n77108 , n77082 , n77107 );
and ( n77109 , n75953 , n75957 );
and ( n77110 , n75957 , n75963 );
and ( n77111 , n75953 , n75963 );
or ( n77112 , n77109 , n77110 , n77111 );
and ( n77113 , n75943 , n75944 );
and ( n77114 , n75944 , n75946 );
and ( n77115 , n75943 , n75946 );
or ( n77116 , n77113 , n77114 , n77115 );
and ( n77117 , n18144 , n20976 );
and ( n77118 , n19324 , n20156 );
xor ( n77119 , n77117 , n77118 );
and ( n77120 , n20233 , n19222 );
xor ( n77121 , n77119 , n77120 );
xor ( n77122 , n77116 , n77121 );
and ( n77123 , n15758 , n24137 );
and ( n77124 , n16637 , n23075 );
xor ( n77125 , n77123 , n77124 );
and ( n77126 , n17512 , n22065 );
xor ( n77127 , n77125 , n77126 );
xor ( n77128 , n77122 , n77127 );
xor ( n77129 , n77112 , n77128 );
and ( n77130 , n75959 , n75960 );
and ( n77131 , n75960 , n75962 );
and ( n77132 , n75959 , n75962 );
or ( n77133 , n77130 , n77131 , n77132 );
and ( n77134 , n75982 , n75983 );
and ( n77135 , n75983 , n75985 );
and ( n77136 , n75982 , n75985 );
or ( n77137 , n77134 , n77135 , n77136 );
xor ( n77138 , n77133 , n77137 );
and ( n77139 , n13322 , n27296 );
and ( n77140 , n14118 , n26216 );
xor ( n77141 , n77139 , n77140 );
and ( n77142 , n14938 , n25163 );
xor ( n77143 , n77141 , n77142 );
xor ( n77144 , n77138 , n77143 );
xor ( n77145 , n77129 , n77144 );
xor ( n77146 , n77108 , n77145 );
xor ( n77147 , n77078 , n77146 );
and ( n77148 , n75975 , n75976 );
and ( n77149 , n75976 , n75993 );
and ( n77150 , n75975 , n75993 );
or ( n77151 , n77148 , n77149 , n77150 );
and ( n77152 , n75981 , n75986 );
and ( n77153 , n75986 , n75992 );
and ( n77154 , n75981 , n75992 );
or ( n77155 , n77152 , n77153 , n77154 );
and ( n77156 , n75887 , n75890 );
xor ( n77157 , n77155 , n77156 );
and ( n77158 , n75988 , n75989 );
and ( n77159 , n75989 , n75991 );
and ( n77160 , n75988 , n75991 );
or ( n77161 , n77158 , n77159 , n77160 );
and ( n77162 , n11015 , n30629 );
and ( n77163 , n11769 , n29508 );
xor ( n77164 , n77162 , n77163 );
and ( n77165 , n12320 , n28406 );
xor ( n77166 , n77164 , n77165 );
xor ( n77167 , n77161 , n77166 );
not ( n77168 , n8718 );
and ( n77169 , n34193 , n8718 );
nor ( n77170 , n77168 , n77169 );
and ( n77171 , n9400 , n32999 );
xor ( n77172 , n77170 , n77171 );
and ( n77173 , n10291 , n31761 );
xor ( n77174 , n77172 , n77173 );
xor ( n77175 , n77167 , n77174 );
xor ( n77176 , n77157 , n77175 );
xor ( n77177 , n77151 , n77176 );
xor ( n77178 , n77147 , n77177 );
xor ( n77179 , n77077 , n77178 );
xor ( n77180 , n77073 , n77179 );
xor ( n77181 , n76997 , n77180 );
xor ( n77182 , n76988 , n77181 );
and ( n77183 , n75797 , n75800 );
and ( n77184 , n75800 , n76000 );
and ( n77185 , n75797 , n76000 );
or ( n77186 , n77183 , n77184 , n77185 );
xor ( n77187 , n77182 , n77186 );
and ( n77188 , n76001 , n76005 );
and ( n77189 , n76006 , n76009 );
or ( n77190 , n77188 , n77189 );
xor ( n77191 , n77187 , n77190 );
buf ( n77192 , n77191 );
buf ( n77193 , n77192 );
not ( n77194 , n77193 );
and ( n77195 , n77194 , n8738 );
nor ( n77196 , n77195 , n8739 );
xor ( n77197 , n76980 , n77196 );
and ( n77198 , n75793 , n76014 );
and ( n77199 , n76015 , n76018 );
or ( n77200 , n77198 , n77199 );
xor ( n77201 , n77197 , n77200 );
buf ( n77202 , n77201 );
buf ( n77203 , n77202 );
not ( n77204 , n77203 );
buf ( n77205 , n598 );
and ( n77206 , n77204 , n77205 );
not ( n77207 , n77205 );
nor ( n77208 , n77206 , n77207 );
xor ( n77209 , n76606 , n77208 );
xor ( n77210 , n76030 , n76603 );
nor ( n77211 , n76022 , n77207 );
and ( n77212 , n77210 , n77211 );
xor ( n77213 , n77210 , n77211 );
xor ( n77214 , n76034 , n76601 );
nor ( n77215 , n74841 , n77207 );
and ( n77216 , n77214 , n77215 );
xor ( n77217 , n77214 , n77215 );
xor ( n77218 , n76038 , n76599 );
nor ( n77219 , n73663 , n77207 );
and ( n77220 , n77218 , n77219 );
xor ( n77221 , n77218 , n77219 );
xor ( n77222 , n76042 , n76597 );
nor ( n77223 , n72481 , n77207 );
and ( n77224 , n77222 , n77223 );
xor ( n77225 , n77222 , n77223 );
xor ( n77226 , n76046 , n76595 );
nor ( n77227 , n71301 , n77207 );
and ( n77228 , n77226 , n77227 );
xor ( n77229 , n77226 , n77227 );
xor ( n77230 , n76050 , n76593 );
nor ( n77231 , n70119 , n77207 );
and ( n77232 , n77230 , n77231 );
xor ( n77233 , n77230 , n77231 );
xor ( n77234 , n76054 , n76591 );
nor ( n77235 , n68933 , n77207 );
and ( n77236 , n77234 , n77235 );
xor ( n77237 , n77234 , n77235 );
xor ( n77238 , n76058 , n76589 );
nor ( n77239 , n67745 , n77207 );
and ( n77240 , n77238 , n77239 );
xor ( n77241 , n77238 , n77239 );
xor ( n77242 , n76062 , n76587 );
nor ( n77243 , n66559 , n77207 );
and ( n77244 , n77242 , n77243 );
xor ( n77245 , n77242 , n77243 );
xor ( n77246 , n76066 , n76585 );
nor ( n77247 , n65369 , n77207 );
and ( n77248 , n77246 , n77247 );
xor ( n77249 , n77246 , n77247 );
xor ( n77250 , n76070 , n76583 );
nor ( n77251 , n64181 , n77207 );
and ( n77252 , n77250 , n77251 );
xor ( n77253 , n77250 , n77251 );
xor ( n77254 , n76074 , n76581 );
nor ( n77255 , n62991 , n77207 );
and ( n77256 , n77254 , n77255 );
xor ( n77257 , n77254 , n77255 );
xor ( n77258 , n76078 , n76579 );
nor ( n77259 , n61800 , n77207 );
and ( n77260 , n77258 , n77259 );
xor ( n77261 , n77258 , n77259 );
xor ( n77262 , n76082 , n76577 );
nor ( n77263 , n60609 , n77207 );
and ( n77264 , n77262 , n77263 );
xor ( n77265 , n77262 , n77263 );
xor ( n77266 , n76086 , n76575 );
nor ( n77267 , n59421 , n77207 );
and ( n77268 , n77266 , n77267 );
xor ( n77269 , n77266 , n77267 );
xor ( n77270 , n76090 , n76573 );
nor ( n77271 , n58226 , n77207 );
and ( n77272 , n77270 , n77271 );
xor ( n77273 , n77270 , n77271 );
xor ( n77274 , n76094 , n76571 );
nor ( n77275 , n57031 , n77207 );
and ( n77276 , n77274 , n77275 );
xor ( n77277 , n77274 , n77275 );
xor ( n77278 , n76098 , n76569 );
nor ( n77279 , n55835 , n77207 );
and ( n77280 , n77278 , n77279 );
xor ( n77281 , n77278 , n77279 );
xor ( n77282 , n76102 , n76567 );
nor ( n77283 , n54638 , n77207 );
and ( n77284 , n77282 , n77283 );
xor ( n77285 , n77282 , n77283 );
xor ( n77286 , n76106 , n76565 );
nor ( n77287 , n53441 , n77207 );
and ( n77288 , n77286 , n77287 );
xor ( n77289 , n77286 , n77287 );
xor ( n77290 , n76110 , n76563 );
nor ( n77291 , n52247 , n77207 );
and ( n77292 , n77290 , n77291 );
xor ( n77293 , n77290 , n77291 );
xor ( n77294 , n76114 , n76561 );
nor ( n77295 , n51049 , n77207 );
and ( n77296 , n77294 , n77295 );
xor ( n77297 , n77294 , n77295 );
xor ( n77298 , n76118 , n76559 );
nor ( n77299 , n49850 , n77207 );
and ( n77300 , n77298 , n77299 );
xor ( n77301 , n77298 , n77299 );
xor ( n77302 , n76122 , n76557 );
nor ( n77303 , n48650 , n77207 );
and ( n77304 , n77302 , n77303 );
xor ( n77305 , n77302 , n77303 );
xor ( n77306 , n76126 , n76555 );
nor ( n77307 , n47449 , n77207 );
and ( n77308 , n77306 , n77307 );
xor ( n77309 , n77306 , n77307 );
xor ( n77310 , n76130 , n76553 );
nor ( n77311 , n46248 , n77207 );
and ( n77312 , n77310 , n77311 );
xor ( n77313 , n77310 , n77311 );
xor ( n77314 , n76134 , n76551 );
nor ( n77315 , n45047 , n77207 );
and ( n77316 , n77314 , n77315 );
xor ( n77317 , n77314 , n77315 );
xor ( n77318 , n76138 , n76549 );
nor ( n77319 , n43843 , n77207 );
and ( n77320 , n77318 , n77319 );
xor ( n77321 , n77318 , n77319 );
xor ( n77322 , n76142 , n76547 );
nor ( n77323 , n42641 , n77207 );
and ( n77324 , n77322 , n77323 );
xor ( n77325 , n77322 , n77323 );
xor ( n77326 , n76146 , n76545 );
nor ( n77327 , n41437 , n77207 );
and ( n77328 , n77326 , n77327 );
xor ( n77329 , n77326 , n77327 );
xor ( n77330 , n76150 , n76543 );
nor ( n77331 , n40232 , n77207 );
and ( n77332 , n77330 , n77331 );
xor ( n77333 , n77330 , n77331 );
xor ( n77334 , n76154 , n76541 );
nor ( n77335 , n39027 , n77207 );
and ( n77336 , n77334 , n77335 );
xor ( n77337 , n77334 , n77335 );
xor ( n77338 , n76158 , n76539 );
nor ( n77339 , n37825 , n77207 );
and ( n77340 , n77338 , n77339 );
xor ( n77341 , n77338 , n77339 );
xor ( n77342 , n76162 , n76537 );
nor ( n77343 , n36620 , n77207 );
and ( n77344 , n77342 , n77343 );
xor ( n77345 , n77342 , n77343 );
xor ( n77346 , n76166 , n76535 );
nor ( n77347 , n35419 , n77207 );
and ( n77348 , n77346 , n77347 );
xor ( n77349 , n77346 , n77347 );
xor ( n77350 , n76170 , n76533 );
nor ( n77351 , n34224 , n77207 );
and ( n77352 , n77350 , n77351 );
xor ( n77353 , n77350 , n77351 );
xor ( n77354 , n76174 , n76531 );
nor ( n77355 , n33033 , n77207 );
and ( n77356 , n77354 , n77355 );
xor ( n77357 , n77354 , n77355 );
xor ( n77358 , n76178 , n76529 );
nor ( n77359 , n31867 , n77207 );
and ( n77360 , n77358 , n77359 );
xor ( n77361 , n77358 , n77359 );
xor ( n77362 , n76182 , n76527 );
nor ( n77363 , n30725 , n77207 );
and ( n77364 , n77362 , n77363 );
xor ( n77365 , n77362 , n77363 );
xor ( n77366 , n76186 , n76525 );
nor ( n77367 , n29596 , n77207 );
and ( n77368 , n77366 , n77367 );
xor ( n77369 , n77366 , n77367 );
xor ( n77370 , n76190 , n76523 );
nor ( n77371 , n28487 , n77207 );
and ( n77372 , n77370 , n77371 );
xor ( n77373 , n77370 , n77371 );
xor ( n77374 , n76194 , n76521 );
nor ( n77375 , n27397 , n77207 );
and ( n77376 , n77374 , n77375 );
xor ( n77377 , n77374 , n77375 );
xor ( n77378 , n76198 , n76519 );
nor ( n77379 , n26326 , n77207 );
and ( n77380 , n77378 , n77379 );
xor ( n77381 , n77378 , n77379 );
xor ( n77382 , n76202 , n76517 );
nor ( n77383 , n25272 , n77207 );
and ( n77384 , n77382 , n77383 );
xor ( n77385 , n77382 , n77383 );
xor ( n77386 , n76206 , n76515 );
nor ( n77387 , n24242 , n77207 );
and ( n77388 , n77386 , n77387 );
xor ( n77389 , n77386 , n77387 );
xor ( n77390 , n76210 , n76513 );
nor ( n77391 , n23225 , n77207 );
and ( n77392 , n77390 , n77391 );
xor ( n77393 , n77390 , n77391 );
xor ( n77394 , n76214 , n76511 );
nor ( n77395 , n22231 , n77207 );
and ( n77396 , n77394 , n77395 );
xor ( n77397 , n77394 , n77395 );
xor ( n77398 , n76218 , n76509 );
nor ( n77399 , n21258 , n77207 );
and ( n77400 , n77398 , n77399 );
xor ( n77401 , n77398 , n77399 );
xor ( n77402 , n76222 , n76507 );
nor ( n77403 , n20303 , n77207 );
and ( n77404 , n77402 , n77403 );
xor ( n77405 , n77402 , n77403 );
xor ( n77406 , n76226 , n76505 );
nor ( n77407 , n19365 , n77207 );
and ( n77408 , n77406 , n77407 );
xor ( n77409 , n77406 , n77407 );
xor ( n77410 , n76230 , n76503 );
nor ( n77411 , n18448 , n77207 );
and ( n77412 , n77410 , n77411 );
xor ( n77413 , n77410 , n77411 );
xor ( n77414 , n76234 , n76501 );
nor ( n77415 , n17548 , n77207 );
and ( n77416 , n77414 , n77415 );
xor ( n77417 , n77414 , n77415 );
xor ( n77418 , n76238 , n76499 );
nor ( n77419 , n16669 , n77207 );
and ( n77420 , n77418 , n77419 );
xor ( n77421 , n77418 , n77419 );
xor ( n77422 , n76242 , n76497 );
nor ( n77423 , n15809 , n77207 );
and ( n77424 , n77422 , n77423 );
xor ( n77425 , n77422 , n77423 );
xor ( n77426 , n76246 , n76495 );
nor ( n77427 , n14968 , n77207 );
and ( n77428 , n77426 , n77427 );
xor ( n77429 , n77426 , n77427 );
xor ( n77430 , n76250 , n76493 );
nor ( n77431 , n14147 , n77207 );
and ( n77432 , n77430 , n77431 );
xor ( n77433 , n77430 , n77431 );
xor ( n77434 , n76254 , n76491 );
nor ( n77435 , n13349 , n77207 );
and ( n77436 , n77434 , n77435 );
xor ( n77437 , n77434 , n77435 );
xor ( n77438 , n76258 , n76489 );
nor ( n77439 , n12564 , n77207 );
and ( n77440 , n77438 , n77439 );
xor ( n77441 , n77438 , n77439 );
xor ( n77442 , n76262 , n76487 );
nor ( n77443 , n11799 , n77207 );
and ( n77444 , n77442 , n77443 );
xor ( n77445 , n77442 , n77443 );
xor ( n77446 , n76266 , n76485 );
nor ( n77447 , n11050 , n77207 );
and ( n77448 , n77446 , n77447 );
xor ( n77449 , n77446 , n77447 );
xor ( n77450 , n76270 , n76483 );
nor ( n77451 , n10321 , n77207 );
and ( n77452 , n77450 , n77451 );
xor ( n77453 , n77450 , n77451 );
xor ( n77454 , n76274 , n76481 );
nor ( n77455 , n9429 , n77207 );
and ( n77456 , n77454 , n77455 );
xor ( n77457 , n77454 , n77455 );
xor ( n77458 , n76278 , n76479 );
nor ( n77459 , n8949 , n77207 );
and ( n77460 , n77458 , n77459 );
xor ( n77461 , n77458 , n77459 );
xor ( n77462 , n76282 , n76477 );
nor ( n77463 , n9437 , n77207 );
and ( n77464 , n77462 , n77463 );
xor ( n77465 , n77462 , n77463 );
xor ( n77466 , n76286 , n76475 );
nor ( n77467 , n9446 , n77207 );
and ( n77468 , n77466 , n77467 );
xor ( n77469 , n77466 , n77467 );
xor ( n77470 , n76290 , n76473 );
nor ( n77471 , n9455 , n77207 );
and ( n77472 , n77470 , n77471 );
xor ( n77473 , n77470 , n77471 );
xor ( n77474 , n76294 , n76471 );
nor ( n77475 , n9464 , n77207 );
and ( n77476 , n77474 , n77475 );
xor ( n77477 , n77474 , n77475 );
xor ( n77478 , n76298 , n76469 );
nor ( n77479 , n9473 , n77207 );
and ( n77480 , n77478 , n77479 );
xor ( n77481 , n77478 , n77479 );
xor ( n77482 , n76302 , n76467 );
nor ( n77483 , n9482 , n77207 );
and ( n77484 , n77482 , n77483 );
xor ( n77485 , n77482 , n77483 );
xor ( n77486 , n76306 , n76465 );
nor ( n77487 , n9491 , n77207 );
and ( n77488 , n77486 , n77487 );
xor ( n77489 , n77486 , n77487 );
xor ( n77490 , n76310 , n76463 );
nor ( n77491 , n9500 , n77207 );
and ( n77492 , n77490 , n77491 );
xor ( n77493 , n77490 , n77491 );
xor ( n77494 , n76314 , n76461 );
nor ( n77495 , n9509 , n77207 );
and ( n77496 , n77494 , n77495 );
xor ( n77497 , n77494 , n77495 );
xor ( n77498 , n76318 , n76459 );
nor ( n77499 , n9518 , n77207 );
and ( n77500 , n77498 , n77499 );
xor ( n77501 , n77498 , n77499 );
xor ( n77502 , n76322 , n76457 );
nor ( n77503 , n9527 , n77207 );
and ( n77504 , n77502 , n77503 );
xor ( n77505 , n77502 , n77503 );
xor ( n77506 , n76326 , n76455 );
nor ( n77507 , n9536 , n77207 );
and ( n77508 , n77506 , n77507 );
xor ( n77509 , n77506 , n77507 );
xor ( n77510 , n76330 , n76453 );
nor ( n77511 , n9545 , n77207 );
and ( n77512 , n77510 , n77511 );
xor ( n77513 , n77510 , n77511 );
xor ( n77514 , n76334 , n76451 );
nor ( n77515 , n9554 , n77207 );
and ( n77516 , n77514 , n77515 );
xor ( n77517 , n77514 , n77515 );
xor ( n77518 , n76338 , n76449 );
nor ( n77519 , n9563 , n77207 );
and ( n77520 , n77518 , n77519 );
xor ( n77521 , n77518 , n77519 );
xor ( n77522 , n76342 , n76447 );
nor ( n77523 , n9572 , n77207 );
and ( n77524 , n77522 , n77523 );
xor ( n77525 , n77522 , n77523 );
xor ( n77526 , n76346 , n76445 );
nor ( n77527 , n9581 , n77207 );
and ( n77528 , n77526 , n77527 );
xor ( n77529 , n77526 , n77527 );
xor ( n77530 , n76350 , n76443 );
nor ( n77531 , n9590 , n77207 );
and ( n77532 , n77530 , n77531 );
xor ( n77533 , n77530 , n77531 );
xor ( n77534 , n76354 , n76441 );
nor ( n77535 , n9599 , n77207 );
and ( n77536 , n77534 , n77535 );
xor ( n77537 , n77534 , n77535 );
xor ( n77538 , n76358 , n76439 );
nor ( n77539 , n9608 , n77207 );
and ( n77540 , n77538 , n77539 );
xor ( n77541 , n77538 , n77539 );
xor ( n77542 , n76362 , n76437 );
nor ( n77543 , n9617 , n77207 );
and ( n77544 , n77542 , n77543 );
xor ( n77545 , n77542 , n77543 );
xor ( n77546 , n76366 , n76435 );
nor ( n77547 , n9626 , n77207 );
and ( n77548 , n77546 , n77547 );
xor ( n77549 , n77546 , n77547 );
xor ( n77550 , n76370 , n76433 );
nor ( n77551 , n9635 , n77207 );
and ( n77552 , n77550 , n77551 );
xor ( n77553 , n77550 , n77551 );
xor ( n77554 , n76374 , n76431 );
nor ( n77555 , n9644 , n77207 );
and ( n77556 , n77554 , n77555 );
xor ( n77557 , n77554 , n77555 );
xor ( n77558 , n76378 , n76429 );
nor ( n77559 , n9653 , n77207 );
and ( n77560 , n77558 , n77559 );
xor ( n77561 , n77558 , n77559 );
xor ( n77562 , n76382 , n76427 );
nor ( n77563 , n9662 , n77207 );
and ( n77564 , n77562 , n77563 );
xor ( n77565 , n77562 , n77563 );
xor ( n77566 , n76386 , n76425 );
nor ( n77567 , n9671 , n77207 );
and ( n77568 , n77566 , n77567 );
xor ( n77569 , n77566 , n77567 );
xor ( n77570 , n76390 , n76423 );
nor ( n77571 , n9680 , n77207 );
and ( n77572 , n77570 , n77571 );
xor ( n77573 , n77570 , n77571 );
xor ( n77574 , n76394 , n76421 );
nor ( n77575 , n9689 , n77207 );
and ( n77576 , n77574 , n77575 );
xor ( n77577 , n77574 , n77575 );
xor ( n77578 , n76398 , n76419 );
nor ( n77579 , n9698 , n77207 );
and ( n77580 , n77578 , n77579 );
xor ( n77581 , n77578 , n77579 );
xor ( n77582 , n76402 , n76417 );
nor ( n77583 , n9707 , n77207 );
and ( n77584 , n77582 , n77583 );
xor ( n77585 , n77582 , n77583 );
xor ( n77586 , n76406 , n76415 );
nor ( n77587 , n9716 , n77207 );
and ( n77588 , n77586 , n77587 );
xor ( n77589 , n77586 , n77587 );
xor ( n77590 , n76410 , n76413 );
nor ( n77591 , n9725 , n77207 );
and ( n77592 , n77590 , n77591 );
xor ( n77593 , n77590 , n77591 );
xor ( n77594 , n76411 , n76412 );
nor ( n77595 , n9734 , n77207 );
and ( n77596 , n77594 , n77595 );
xor ( n77597 , n77594 , n77595 );
nor ( n77598 , n9752 , n76024 );
nor ( n77599 , n9743 , n77207 );
and ( n77600 , n77598 , n77599 );
and ( n77601 , n77597 , n77600 );
or ( n77602 , n77596 , n77601 );
and ( n77603 , n77593 , n77602 );
or ( n77604 , n77592 , n77603 );
and ( n77605 , n77589 , n77604 );
or ( n77606 , n77588 , n77605 );
and ( n77607 , n77585 , n77606 );
or ( n77608 , n77584 , n77607 );
and ( n77609 , n77581 , n77608 );
or ( n77610 , n77580 , n77609 );
and ( n77611 , n77577 , n77610 );
or ( n77612 , n77576 , n77611 );
and ( n77613 , n77573 , n77612 );
or ( n77614 , n77572 , n77613 );
and ( n77615 , n77569 , n77614 );
or ( n77616 , n77568 , n77615 );
and ( n77617 , n77565 , n77616 );
or ( n77618 , n77564 , n77617 );
and ( n77619 , n77561 , n77618 );
or ( n77620 , n77560 , n77619 );
and ( n77621 , n77557 , n77620 );
or ( n77622 , n77556 , n77621 );
and ( n77623 , n77553 , n77622 );
or ( n77624 , n77552 , n77623 );
and ( n77625 , n77549 , n77624 );
or ( n77626 , n77548 , n77625 );
and ( n77627 , n77545 , n77626 );
or ( n77628 , n77544 , n77627 );
and ( n77629 , n77541 , n77628 );
or ( n77630 , n77540 , n77629 );
and ( n77631 , n77537 , n77630 );
or ( n77632 , n77536 , n77631 );
and ( n77633 , n77533 , n77632 );
or ( n77634 , n77532 , n77633 );
and ( n77635 , n77529 , n77634 );
or ( n77636 , n77528 , n77635 );
and ( n77637 , n77525 , n77636 );
or ( n77638 , n77524 , n77637 );
and ( n77639 , n77521 , n77638 );
or ( n77640 , n77520 , n77639 );
and ( n77641 , n77517 , n77640 );
or ( n77642 , n77516 , n77641 );
and ( n77643 , n77513 , n77642 );
or ( n77644 , n77512 , n77643 );
and ( n77645 , n77509 , n77644 );
or ( n77646 , n77508 , n77645 );
and ( n77647 , n77505 , n77646 );
or ( n77648 , n77504 , n77647 );
and ( n77649 , n77501 , n77648 );
or ( n77650 , n77500 , n77649 );
and ( n77651 , n77497 , n77650 );
or ( n77652 , n77496 , n77651 );
and ( n77653 , n77493 , n77652 );
or ( n77654 , n77492 , n77653 );
and ( n77655 , n77489 , n77654 );
or ( n77656 , n77488 , n77655 );
and ( n77657 , n77485 , n77656 );
or ( n77658 , n77484 , n77657 );
and ( n77659 , n77481 , n77658 );
or ( n77660 , n77480 , n77659 );
and ( n77661 , n77477 , n77660 );
or ( n77662 , n77476 , n77661 );
and ( n77663 , n77473 , n77662 );
or ( n77664 , n77472 , n77663 );
and ( n77665 , n77469 , n77664 );
or ( n77666 , n77468 , n77665 );
and ( n77667 , n77465 , n77666 );
or ( n77668 , n77464 , n77667 );
and ( n77669 , n77461 , n77668 );
or ( n77670 , n77460 , n77669 );
and ( n77671 , n77457 , n77670 );
or ( n77672 , n77456 , n77671 );
and ( n77673 , n77453 , n77672 );
or ( n77674 , n77452 , n77673 );
and ( n77675 , n77449 , n77674 );
or ( n77676 , n77448 , n77675 );
and ( n77677 , n77445 , n77676 );
or ( n77678 , n77444 , n77677 );
and ( n77679 , n77441 , n77678 );
or ( n77680 , n77440 , n77679 );
and ( n77681 , n77437 , n77680 );
or ( n77682 , n77436 , n77681 );
and ( n77683 , n77433 , n77682 );
or ( n77684 , n77432 , n77683 );
and ( n77685 , n77429 , n77684 );
or ( n77686 , n77428 , n77685 );
and ( n77687 , n77425 , n77686 );
or ( n77688 , n77424 , n77687 );
and ( n77689 , n77421 , n77688 );
or ( n77690 , n77420 , n77689 );
and ( n77691 , n77417 , n77690 );
or ( n77692 , n77416 , n77691 );
and ( n77693 , n77413 , n77692 );
or ( n77694 , n77412 , n77693 );
and ( n77695 , n77409 , n77694 );
or ( n77696 , n77408 , n77695 );
and ( n77697 , n77405 , n77696 );
or ( n77698 , n77404 , n77697 );
and ( n77699 , n77401 , n77698 );
or ( n77700 , n77400 , n77699 );
and ( n77701 , n77397 , n77700 );
or ( n77702 , n77396 , n77701 );
and ( n77703 , n77393 , n77702 );
or ( n77704 , n77392 , n77703 );
and ( n77705 , n77389 , n77704 );
or ( n77706 , n77388 , n77705 );
and ( n77707 , n77385 , n77706 );
or ( n77708 , n77384 , n77707 );
and ( n77709 , n77381 , n77708 );
or ( n77710 , n77380 , n77709 );
and ( n77711 , n77377 , n77710 );
or ( n77712 , n77376 , n77711 );
and ( n77713 , n77373 , n77712 );
or ( n77714 , n77372 , n77713 );
and ( n77715 , n77369 , n77714 );
or ( n77716 , n77368 , n77715 );
and ( n77717 , n77365 , n77716 );
or ( n77718 , n77364 , n77717 );
and ( n77719 , n77361 , n77718 );
or ( n77720 , n77360 , n77719 );
and ( n77721 , n77357 , n77720 );
or ( n77722 , n77356 , n77721 );
and ( n77723 , n77353 , n77722 );
or ( n77724 , n77352 , n77723 );
and ( n77725 , n77349 , n77724 );
or ( n77726 , n77348 , n77725 );
and ( n77727 , n77345 , n77726 );
or ( n77728 , n77344 , n77727 );
and ( n77729 , n77341 , n77728 );
or ( n77730 , n77340 , n77729 );
and ( n77731 , n77337 , n77730 );
or ( n77732 , n77336 , n77731 );
and ( n77733 , n77333 , n77732 );
or ( n77734 , n77332 , n77733 );
and ( n77735 , n77329 , n77734 );
or ( n77736 , n77328 , n77735 );
and ( n77737 , n77325 , n77736 );
or ( n77738 , n77324 , n77737 );
and ( n77739 , n77321 , n77738 );
or ( n77740 , n77320 , n77739 );
and ( n77741 , n77317 , n77740 );
or ( n77742 , n77316 , n77741 );
and ( n77743 , n77313 , n77742 );
or ( n77744 , n77312 , n77743 );
and ( n77745 , n77309 , n77744 );
or ( n77746 , n77308 , n77745 );
and ( n77747 , n77305 , n77746 );
or ( n77748 , n77304 , n77747 );
and ( n77749 , n77301 , n77748 );
or ( n77750 , n77300 , n77749 );
and ( n77751 , n77297 , n77750 );
or ( n77752 , n77296 , n77751 );
and ( n77753 , n77293 , n77752 );
or ( n77754 , n77292 , n77753 );
and ( n77755 , n77289 , n77754 );
or ( n77756 , n77288 , n77755 );
and ( n77757 , n77285 , n77756 );
or ( n77758 , n77284 , n77757 );
and ( n77759 , n77281 , n77758 );
or ( n77760 , n77280 , n77759 );
and ( n77761 , n77277 , n77760 );
or ( n77762 , n77276 , n77761 );
and ( n77763 , n77273 , n77762 );
or ( n77764 , n77272 , n77763 );
and ( n77765 , n77269 , n77764 );
or ( n77766 , n77268 , n77765 );
and ( n77767 , n77265 , n77766 );
or ( n77768 , n77264 , n77767 );
and ( n77769 , n77261 , n77768 );
or ( n77770 , n77260 , n77769 );
and ( n77771 , n77257 , n77770 );
or ( n77772 , n77256 , n77771 );
and ( n77773 , n77253 , n77772 );
or ( n77774 , n77252 , n77773 );
and ( n77775 , n77249 , n77774 );
or ( n77776 , n77248 , n77775 );
and ( n77777 , n77245 , n77776 );
or ( n77778 , n77244 , n77777 );
and ( n77779 , n77241 , n77778 );
or ( n77780 , n77240 , n77779 );
and ( n77781 , n77237 , n77780 );
or ( n77782 , n77236 , n77781 );
and ( n77783 , n77233 , n77782 );
or ( n77784 , n77232 , n77783 );
and ( n77785 , n77229 , n77784 );
or ( n77786 , n77228 , n77785 );
and ( n77787 , n77225 , n77786 );
or ( n77788 , n77224 , n77787 );
and ( n77789 , n77221 , n77788 );
or ( n77790 , n77220 , n77789 );
and ( n77791 , n77217 , n77790 );
or ( n77792 , n77216 , n77791 );
and ( n77793 , n77213 , n77792 );
or ( n77794 , n77212 , n77793 );
xor ( n77795 , n77209 , n77794 );
buf ( n77796 , n77795 );
buf ( n77797 , n77796 );
xor ( n77798 , n77213 , n77792 );
buf ( n77799 , n77798 );
buf ( n77800 , n77799 );
xor ( n77801 , n77217 , n77790 );
buf ( n77802 , n77801 );
buf ( n77803 , n77802 );
xor ( n77804 , n77221 , n77788 );
buf ( n77805 , n77804 );
buf ( n77806 , n77805 );
xor ( n77807 , n77225 , n77786 );
buf ( n77808 , n77807 );
buf ( n77809 , n77808 );
xor ( n77810 , n77229 , n77784 );
buf ( n77811 , n77810 );
buf ( n77812 , n77811 );
xor ( n77813 , n77233 , n77782 );
buf ( n77814 , n77813 );
buf ( n77815 , n77814 );
xor ( n77816 , n77237 , n77780 );
buf ( n77817 , n77816 );
buf ( n77818 , n77817 );
xor ( n77819 , n77241 , n77778 );
buf ( n77820 , n77819 );
buf ( n77821 , n77820 );
xor ( n77822 , n77245 , n77776 );
buf ( n77823 , n77822 );
buf ( n77824 , n77823 );
endmodule
