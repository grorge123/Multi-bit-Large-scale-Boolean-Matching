module top( n5 , n16 , n23 , n24 , n31 , n38 , n41 , n44 , n46 ,
n53 , n55 , n57 , n62 , n63 , n68 , n71 , n72 , n78 , n79 ,
n84 , n92 , n96 , n98 , n101 , n106 , n107 , n120 , n123 , n126 ,
n136 , n142 , n144 , n145 , n153 , n165 , n177 , n182 , n216 , n220 );
    input n16 , n23 , n24 , n31 , n38 , n41 , n44 , n46 , n53 ,
n55 , n57 , n62 , n68 , n71 , n72 , n79 , n84 , n92 , n96 ,
n98 , n101 , n106 , n107 , n120 , n123 , n136 , n145 , n165 , n177 ,
n182 , n216 , n220 ;
    output n5 , n63 , n78 , n126 , n142 , n144 , n153 ;
    wire n0 , n1 , n2 , n3 , n4 , n6 , n7 , n8 , n9 ,
n10 , n11 , n12 , n13 , n14 , n15 , n17 , n18 , n19 , n20 ,
n21 , n22 , n25 , n26 , n27 , n28 , n29 , n30 , n32 , n33 ,
n34 , n35 , n36 , n37 , n39 , n40 , n42 , n43 , n45 , n47 ,
n48 , n49 , n50 , n51 , n52 , n54 , n56 , n58 , n59 , n60 ,
n61 , n64 , n65 , n66 , n67 , n69 , n70 , n73 , n74 , n75 ,
n76 , n77 , n80 , n81 , n82 , n83 , n85 , n86 , n87 , n88 ,
n89 , n90 , n91 , n93 , n94 , n95 , n97 , n99 , n100 , n102 ,
n103 , n104 , n105 , n108 , n109 , n110 , n111 , n112 , n113 , n114 ,
n115 , n116 , n117 , n118 , n119 , n121 , n122 , n124 , n125 , n127 ,
n128 , n129 , n130 , n131 , n132 , n133 , n134 , n135 , n137 , n138 ,
n139 , n140 , n141 , n143 , n146 , n147 , n148 , n149 , n150 , n151 ,
n152 , n154 , n155 , n156 , n157 , n158 , n159 , n160 , n161 , n162 ,
n163 , n164 , n166 , n167 , n168 , n169 , n170 , n171 , n172 , n173 ,
n174 , n175 , n176 , n178 , n179 , n180 , n181 , n183 , n184 , n185 ,
n186 , n187 , n188 , n189 , n190 , n191 , n192 , n193 , n194 , n195 ,
n196 , n197 , n198 , n199 , n200 , n201 , n202 , n203 , n204 , n205 ,
n206 , n207 , n208 , n209 , n210 , n211 , n212 , n213 , n214 , n215 ,
n217 , n218 , n219 , n221 , n222 , n223 , n224 , n225 , n226 , n227 ,
n228 , n229 , n230 ;
    not g0 ( n17 , n38 );
    and g1 ( n211 , n18 , n116 );
    not g2 ( n193 , n195 );
    and g3 ( n81 , n118 , n84 );
    or g4 ( n75 , n173 , n113 );
    and g5 ( n180 , n132 , n55 );
    and g6 ( n89 , n125 , n136 );
    or g7 ( n103 , n164 , n131 );
    and g8 ( n127 , n226 , n176 );
    nor g9 ( n155 , n198 , n179 );
    not g10 ( n18 , n195 );
    and g11 ( n21 , n180 , n59 );
    and g12 ( n42 , n121 , n170 );
    and g13 ( n209 , n159 , n98 );
    nor g14 ( n28 , n107 , n70 );
    and g15 ( n135 , n139 , n96 );
    or g16 ( n100 , n209 , n1 );
    or g17 ( n172 , n8 , n230 );
    or g18 ( n78 , n97 , n115 );
    or g19 ( n186 , n229 , n86 );
    and g20 ( n111 , n28 , n68 );
    not g21 ( n88 , n37 );
    not g22 ( n95 , n129 );
    and g23 ( n199 , n193 , n71 );
    nor g24 ( n2 , n190 , n118 );
    not g25 ( n47 , n61 );
    or g26 ( n179 , n199 , n81 );
    nor g27 ( n200 , n58 , n194 );
    and g28 ( n205 , n155 , n38 );
    nor g29 ( n26 , n75 , n115 );
    not g30 ( n105 , n170 );
    and g31 ( n152 , n153 , n120 );
    and g32 ( n131 , n88 , n31 );
    not g33 ( n201 , n212 );
    and g34 ( n80 , n227 , n53 );
    not g35 ( n217 , n67 );
    or g36 ( n51 , n41 , n7 );
    and g37 ( n109 , n218 , n10 );
    nor g38 ( n11 , n33 , n64 );
    and g39 ( n215 , n80 , n50 );
    not g40 ( n52 , n106 );
    not g41 ( n159 , n47 );
    nor g42 ( n114 , n157 , n125 );
    nor g43 ( n110 , n79 , n82 );
    and g44 ( n83 , n95 , n79 );
    or g45 ( n133 , n171 , n2 );
    and g46 ( n162 , n66 , n9 );
    not g47 ( n112 , n182 );
    nor g48 ( n138 , n89 , n102 );
    not g49 ( n174 , n217 );
    or g50 ( n39 , n50 , n204 );
    and g51 ( n99 , n0 , n35 );
    or g52 ( n116 , n71 , n17 );
    and g53 ( n50 , n25 , n53 );
    and g54 ( n70 , n5 , n206 );
    and g55 ( n194 , n138 , n53 );
    and g56 ( n160 , n6 , n11 );
    and g57 ( n82 , n159 , n163 );
    and g58 ( n212 , n223 , n51 );
    and g59 ( n161 , n193 , n165 );
    and g60 ( n183 , n171 , n162 );
    nor g61 ( n6 , n181 , n196 );
    or g62 ( n158 , n80 , n137 );
    and g63 ( n91 , n29 , n48 );
    and g64 ( n29 , n210 , n38 );
    or g65 ( n204 , n29 , n221 );
    or g66 ( n102 , n166 , n60 );
    or g67 ( n35 , n169 , n180 );
    and g68 ( n169 , n168 , n182 );
    or g69 ( n32 , n147 , n191 );
    nor g70 ( n25 , n136 , n54 );
    or g71 ( n33 , n119 , n85 );
    and g72 ( n154 , n141 , n51 );
    or g73 ( n73 , n46 , n112 );
    nor g74 ( n139 , n62 , n186 );
    nor g75 ( n227 , n177 , n54 );
    or g76 ( n143 , n172 , n78 );
    nor g77 ( n184 , n31 , n128 );
    or g78 ( n141 , n44 , n77 );
    and g79 ( n59 , n110 , n55 );
    and g80 ( n27 , n213 , n230 );
    and g81 ( n178 , n137 , n111 );
    not g82 ( n124 , n145 );
    or g83 ( n22 , n111 , n108 );
    or g84 ( n148 , n52 , n76 );
    and g85 ( n86 , n153 , n32 );
    not g86 ( n45 , n195 );
    not g87 ( n153 , n49 );
    not g88 ( n214 , n75 );
    not g89 ( n173 , n68 );
    not g90 ( n66 , n190 );
    and g91 ( n74 , n169 , n189 );
    not g92 ( n9 , n92 );
    or g93 ( n134 , n83 , n222 );
    and g94 ( n208 , n34 , n36 );
    not g95 ( n7 , n84 );
    or g96 ( n163 , n165 , n56 );
    or g97 ( n170 , n147 , n104 );
    nor g98 ( n30 , n182 , n143 );
    and g99 ( n54 , n45 , n141 );
    and g100 ( n128 , n90 , n10 );
    not g101 ( n130 , n103 );
    nor g102 ( n157 , n48 , n34 );
    not g103 ( n225 , n13 );
    not g104 ( n5 , n192 );
    nor g105 ( n15 , n185 , n140 );
    and g106 ( n34 , n184 , n84 );
    not g107 ( n12 , n101 );
    and g108 ( n48 , n228 , n7 );
    not g109 ( n10 , n185 );
    and g110 ( n140 , n195 , n84 );
    and g111 ( n171 , n66 , n24 );
    or g112 ( n206 , n57 , n173 );
    and g113 ( n226 , n20 , n116 );
    and g114 ( n4 , n87 , n73 );
    not g115 ( n122 , n211 );
    and g116 ( n63 , n149 , n103 );
    not g117 ( n13 , n40 );
    and g118 ( n20 , n154 , n73 );
    or g119 ( n207 , n91 , n208 );
    or g120 ( n164 , n15 , n152 );
    and g121 ( n166 , n45 , n44 );
    and g122 ( n228 , n122 , n38 );
    not g123 ( n67 , n203 );
    nor g124 ( n121 , n200 , n26 );
    buf g125 ( n0 , n203 );
    nor g126 ( n65 , n189 , n39 );
    not g127 ( n40 , n76 );
    and g128 ( n189 , n175 , n182 );
    nor g129 ( n132 , n16 , n82 );
    nor g130 ( n168 , n220 , n4 );
    nor g131 ( n175 , n123 , n4 );
    nor g132 ( n156 , n216 , n70 );
    or g133 ( n119 , n215 , n178 );
    and g134 ( n94 , n127 , n163 );
    not g135 ( n56 , n55 );
    and g136 ( n60 , n225 , n177 );
    and g137 ( n187 , n201 , n52 );
    or g138 ( n149 , n3 , n42 );
    and g139 ( n76 , n160 , n219 );
    not g140 ( n142 , n13 );
    and g141 ( n198 , n146 , n23 );
    and g142 ( n19 , n146 , n72 );
    and g143 ( n3 , n148 , n201 );
    and g144 ( n185 , n12 , n84 );
    nor g145 ( n144 , n205 , n30 );
    or g146 ( n167 , n74 , n21 );
    and g147 ( n117 , n18 , n57 );
    or g148 ( n181 , n167 , n99 );
    or g149 ( n190 , n124 , n87 );
    or g150 ( n230 , n194 , n214 );
    nor g151 ( n210 , n23 , n211 );
    or g152 ( n191 , n72 , n229 );
    and g153 ( n150 , n88 , n216 );
    not g154 ( n8 , n58 );
    or g155 ( n113 , n224 , n93 );
    nor g156 ( n126 , n97 , n27 );
    and g157 ( n36 , n43 , n84 );
    or g158 ( n64 , n207 , n114 );
    or g159 ( n176 , n98 , n147 );
    or g160 ( n196 , n183 , n135 );
    not g161 ( n129 , n67 );
    nor g162 ( n43 , n120 , n128 );
    and g163 ( n218 , n94 , n206 );
    not g164 ( n213 , n115 );
    and g165 ( n137 , n156 , n68 );
    or g166 ( n104 , n19 , n100 );
    not g167 ( n146 , n129 );
    not g168 ( n61 , n109 );
    not g169 ( n49 , n174 );
    or g170 ( n97 , n130 , n3 );
    not g171 ( n188 , n32 );
    and g172 ( n203 , n65 , n212 );
    or g173 ( n197 , n59 , n22 );
    not g174 ( n223 , n140 );
    and g175 ( n202 , n133 , n151 );
    or g176 ( n221 , n36 , n197 );
    not g177 ( n90 , n47 );
    buf g178 ( n195 , n109 );
    and g179 ( n229 , n90 , n176 );
    and g180 ( n85 , n0 , n158 );
    not g181 ( n147 , n96 );
    and g182 ( n69 , n225 , n16 );
    not g183 ( n87 , n192 );
    and g184 ( n224 , n95 , n107 );
    or g185 ( n151 , n9 , n0 );
    not g186 ( n125 , n217 );
    or g187 ( n108 , n188 , n162 );
    or g188 ( n93 , n117 , n150 );
    or g189 ( n115 , n202 , n105 );
    not g190 ( n77 , n53 );
    and g191 ( n1 , n142 , n62 );
    or g192 ( n58 , n56 , n134 );
    not g193 ( n192 , n61 );
    not g194 ( n37 , n40 );
    or g195 ( n222 , n161 , n69 );
    nor g196 ( n219 , n187 , n14 );
    not g197 ( n118 , n37 );
    and g198 ( n14 , n0 , n171 );
endmodule
